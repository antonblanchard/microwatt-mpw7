* NGSPICE file created from RAM32_1RW1R.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlclkp_1 abstract view
.subckt sky130_fd_sc_hd__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

.subckt RAM32_1RW1R A0[0] A0[1] A0[2] A0[3] A0[4] A1[0] A1[1] A1[2] A1[3] A1[4] CLK
+ Di0[0] Di0[10] Di0[11] Di0[12] Di0[13] Di0[14] Di0[15] Di0[16] Di0[17] Di0[18] Di0[19]
+ Di0[1] Di0[20] Di0[21] Di0[22] Di0[23] Di0[24] Di0[25] Di0[26] Di0[27] Di0[28] Di0[29]
+ Di0[2] Di0[30] Di0[31] Di0[32] Di0[33] Di0[34] Di0[35] Di0[36] Di0[37] Di0[38] Di0[39]
+ Di0[3] Di0[40] Di0[41] Di0[42] Di0[43] Di0[44] Di0[45] Di0[46] Di0[47] Di0[48] Di0[49]
+ Di0[4] Di0[50] Di0[51] Di0[52] Di0[53] Di0[54] Di0[55] Di0[56] Di0[57] Di0[58] Di0[59]
+ Di0[5] Di0[60] Di0[61] Di0[62] Di0[63] Di0[6] Di0[7] Di0[8] Di0[9] Do0[0] Do0[10]
+ Do0[11] Do0[12] Do0[13] Do0[14] Do0[15] Do0[16] Do0[17] Do0[18] Do0[19] Do0[1] Do0[20]
+ Do0[21] Do0[22] Do0[23] Do0[24] Do0[25] Do0[26] Do0[27] Do0[28] Do0[29] Do0[2] Do0[30]
+ Do0[31] Do0[32] Do0[33] Do0[34] Do0[35] Do0[36] Do0[37] Do0[38] Do0[39] Do0[3] Do0[40]
+ Do0[41] Do0[42] Do0[43] Do0[44] Do0[45] Do0[46] Do0[47] Do0[48] Do0[49] Do0[4] Do0[50]
+ Do0[51] Do0[52] Do0[53] Do0[54] Do0[55] Do0[56] Do0[57] Do0[58] Do0[59] Do0[5] Do0[60]
+ Do0[61] Do0[62] Do0[63] Do0[6] Do0[7] Do0[8] Do0[9] Do1[0] Do1[10] Do1[11] Do1[12]
+ Do1[13] Do1[14] Do1[15] Do1[16] Do1[17] Do1[18] Do1[19] Do1[1] Do1[20] Do1[21] Do1[22]
+ Do1[23] Do1[24] Do1[25] Do1[26] Do1[27] Do1[28] Do1[29] Do1[2] Do1[30] Do1[31] Do1[32]
+ Do1[33] Do1[34] Do1[35] Do1[36] Do1[37] Do1[38] Do1[39] Do1[3] Do1[40] Do1[41] Do1[42]
+ Do1[43] Do1[44] Do1[45] Do1[46] Do1[47] Do1[48] Do1[49] Do1[4] Do1[50] Do1[51] Do1[52]
+ Do1[53] Do1[54] Do1[55] Do1[56] Do1[57] Do1[58] Do1[59] Do1[5] Do1[60] Do1[61] Do1[62]
+ Do1[63] Do1[6] Do1[7] Do1[8] Do1[9] EN0 EN1 VGND VPWR WE0[0] WE0[1] WE0[2] WE0[3]
+ WE0[4] WE0[5] WE0[6] WE0[7]
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_3_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_24_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XA0BUF\[0\] A0[0] VGND VGND VPWR VPWR A0BUF\[0\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_12_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_12_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_22_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_9_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.CLKBUF CLKBUF/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.CLKBUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_34_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.DEC1.AND0 SLICE\[2\].RAM8.DEC1.AND7/A SLICE\[2\].RAM8.DEC1.AND7/B
+ SLICE\[2\].RAM8.DEC1.AND7/C SLICE\[2\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC1.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
Xtap_34_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.DEC1.ENBUF DEC1.AND0/Y VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC1.AND7/D
+ sky130_fd_sc_hd__clkbuf_2
Xfill_29_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WEBUF\[7\] WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WEBUF\[7\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_10_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_10_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_19_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_19_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_19_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_1_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[2\] Do0_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF0\[58\]/Z
+ VGND VGND VPWR VPWR Do0[58] sky130_fd_sc_hd__dfxtp_1
Xfill_23_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_23_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_23_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_6_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[1\].FLOATBUF0\[14\] TIE0\[1\]/LO FBUFENBUF0\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_6_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_22_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_15_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[5\].FLOATBUF0\[45\] TIE0\[5\]/LO FBUFENBUF0\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV SLICE\[1\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[2\] BYTE\[2\].FLOATBUF1\[18\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV SLICE\[0\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_21_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[4\].DIODE\[5\] BYTE\[4\].FLOATBUF0\[37\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_18_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_18_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF SLICE\[0\].RAM8.DEC0.AND2/X VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_6_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[1\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
Xfill_6_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_20_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[3\] Do1_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF1\[11\]/Z
+ VGND VGND VPWR VPWR Do1[11] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_13_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_16_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_32_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_20_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_20_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[6\] Do0_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF0\[30\]/Z
+ VGND VGND VPWR VPWR Do0[30] sky130_fd_sc_hd__dfxtp_1
Xtap_3_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_29_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_29_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.DEC1.ABUF\[2\] A1BUF\[2\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC1.AND7/C
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XDIBUF\[50\] Di0[50] VGND VGND VPWR VPWR DIBUF\[50\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_9_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_8_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WEBUF\[4\] WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WEBUF\[4\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_33_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_27_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV SLICE\[0\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_15_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_15_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.SEL1BUF SLICE\[2\].RAM8.DEC1.AND0/Y VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[0\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_31_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_31_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.DEC0.AND4 SLICE\[1\].RAM8.DEC0.AND7/A SLICE\[1\].RAM8.DEC0.AND7/B
+ SLICE\[1\].RAM8.DEC0.AND7/C SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[3\].FLOATBUF0\[26\] TIE0\[3\]/LO FBUFENBUF0\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_3_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XFBUFENBUF0\[5\] EN0 VGND VGND VPWR VPWR FBUFENBUF0\[5\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[7\].FLOATBUF0\[57\] TIE0\[7\]/LO FBUFENBUF0\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_7_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_31_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_24_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_17_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_26_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_9_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo1_REG.OUTREG_BYTE\[7\].DIODE\[2\] BYTE\[7\].FLOATBUF1\[58\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[13\] Di0[13] VGND VGND VPWR VPWR DIBUF\[13\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_5_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_5_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[0\].FLOATBUF1\[5\] TIE1\[0\]/LO FBUFENBUF1\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_3_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_24_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_12_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_12_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[6\].Do_FF\[3\] Do1_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF1\[51\]/Z
+ VGND VGND VPWR VPWR Do1[51] sky130_fd_sc_hd__dfxtp_1
Xfill_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV SLICE\[1\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_9_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_9_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.DEC1.AND1 SLICE\[2\].RAM8.DEC1.AND7/C SLICE\[2\].RAM8.DEC1.AND7/B
+ SLICE\[2\].RAM8.DEC1.AND7/A SLICE\[2\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC1.AND1/X
+ sky130_fd_sc_hd__and4bb_2
Xtap_34_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV SLICE\[0\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_10_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[2\] BYTE\[1\].FLOATBUF0\[10\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_19_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_19_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_19_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_1_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_23_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo1_REG.Do_CLKBUF\[7\] Do1_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do1_REG.Do_CLKBUF\[7\]/X
+ sky130_fd_sc_hd__clkbuf_4
Xfill_23_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_23_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_6_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF SLICE\[0\].RAM8.DEC0.AND1/X VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_6_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[6\] BYTE\[3\].FLOATBUF1\[30\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_22_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XTIE0\[7\] VGND VGND VPWR VPWR TIE0\[7\]/HI TIE0\[7\]/LO sky130_fd_sc_hd__conb_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_15_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[3\] Do0_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF0\[3\]/Z
+ VGND VGND VPWR VPWR Do0[3] sky130_fd_sc_hd__dfxtp_1
Xtap_21_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_18_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_18_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_11_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.DEC0.ENBUF DEC0.AND0/Y VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.AND7/D
+ sky130_fd_sc_hd__clkbuf_2
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[7\] Do1_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF1\[23\]/Z
+ VGND VGND VPWR VPWR Do1[23] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_6_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_20_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_16_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_32_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIODE_A0\[0\] A0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_20_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_20_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV SLICE\[1\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_3_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_29_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XWEBUF\[0\] WE0[0] VGND VGND VPWR VPWR WEBUF\[0\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[43\] Di0[43] VGND VGND VPWR VPWR DIBUF\[43\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_9_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_8_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[3\].FLOATBUF1\[31\] TIE1\[3\]/LO FBUFENBUF1\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_33_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_26_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_27_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_27_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[7\].FLOATBUF1\[62\] TIE1\[7\]/LO FBUFENBUF1\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_15_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_31_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_31_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_31_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.DEC0.AND5 SLICE\[1\].RAM8.DEC0.AND7/B SLICE\[1\].RAM8.DEC0.AND7/A
+ SLICE\[1\].RAM8.DEC0.AND7/C SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_3_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[6\].DIODE\[2\] BYTE\[6\].FLOATBUF0\[50\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WEBUF\[0\] WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[0\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_7_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xtap_13_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.SEL1BUF SLICE\[1\].RAM8.DEC1.AND7/X VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[7\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_31_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_24_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_17_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[0\] Do1_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF1\[24\]/Z
+ VGND VGND VPWR VPWR Do1[24] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_26_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_26_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_9_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV SLICE\[1\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_9_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV SLICE\[0\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[3\] Do0_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF0\[43\]/Z
+ VGND VGND VPWR VPWR Do0[43] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_5_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_24_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF SLICE\[0\].RAM8.DEC0.AND0/Y VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_12_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_12_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[3\] BYTE\[0\].FLOATBUF1\[3\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XDo1_REG.OUTREG_BYTE\[7\].Do_FF\[7\] Do1_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF1\[63\]/Z
+ VGND VGND VPWR VPWR Do1[63] sky130_fd_sc_hd__dfxtp_1
Xtap_22_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XBYTE\[0\].FLOATBUF0\[0\] TIE0\[0\]/LO FBUFENBUF0\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
Xfill_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_14_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_9_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_9_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_34_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.DEC1.AND2 SLICE\[2\].RAM8.DEC1.AND7/C SLICE\[2\].RAM8.DEC1.AND7/A
+ SLICE\[2\].RAM8.DEC1.AND7/B SLICE\[2\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC1.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_34_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[1\].FLOATBUF1\[12\] TIE1\[1\]/LO FBUFENBUF1\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[6\] BYTE\[2\].FLOATBUF0\[22\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfill_29_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XBYTE\[5\].FLOATBUF1\[43\] TIE1\[5\]/LO FBUFENBUF1\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_19_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_19_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_1_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_23_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_23_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_6_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_6_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV SLICE\[2\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[7\] Do0_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF0\[15\]/Z
+ VGND VGND VPWR VPWR Do0[15] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_27_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV SLICE\[1\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_18_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_18_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_18_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_11_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_6_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_13_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_32_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_20_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_3_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_29_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_29_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_22_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XDIBUF\[36\] Di0[36] VGND VGND VPWR VPWR DIBUF\[36\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_9_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_8_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.SEL1BUF SLICE\[1\].RAM8.DEC1.AND6/X VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[6\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XBYTE\[3\].FLOATBUF1\[24\] TIE1\[3\]/LO FBUFENBUF1\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[4\].FLOATBUF1\[39\] TIE1\[4\]/LO FBUFENBUF1\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[3\] Di0[3] VGND VGND VPWR VPWR DIBUF\[3\]/X sky130_fd_sc_hd__clkbuf_16
XDo1_REG.OUTREG_BYTE\[5\].DIODE\[3\] BYTE\[5\].FLOATBUF1\[43\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_26_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_27_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_27_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV SLICE\[1\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_15_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_15_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_31_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_31_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.DEC0.AND6 SLICE\[1\].RAM8.DEC0.AND7/A SLICE\[1\].RAM8.DEC0.AND7/B
+ SLICE\[1\].RAM8.DEC0.AND7/C SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_3_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XDo0_REG.OUTREG_BYTE\[7\].DIODE\[6\] BYTE\[7\].FLOATBUF0\[62\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[0\] Do0_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF0\[16\]/Z
+ VGND VGND VPWR VPWR Do0[16] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_7_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[4\].Do_FF\[4\] Do1_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF1\[36\]/Z
+ VGND VGND VPWR VPWR Do1[36] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_31_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_24_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_26_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_9_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[3\].FLOATBUF0\[31\] TIE0\[3\]/LO FBUFENBUF0\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[7\] Do0_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF0\[55\]/Z
+ VGND VGND VPWR VPWR Do0[55] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[7\].FLOATBUF0\[62\] TIE0\[7\]/LO FBUFENBUF0\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[7\] BYTE\[1\].FLOATBUF1\[15\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_12_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XEN1BUF EN1 VGND VGND VPWR VPWR EN1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_22_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_15_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_8_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_0_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_14_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_9_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_9_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV SLICE\[2\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.DEC1.AND3 SLICE\[2\].RAM8.DEC1.AND7/C SLICE\[2\].RAM8.DEC1.AND7/B
+ SLICE\[2\].RAM8.DEC1.AND7/A SLICE\[2\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC1.AND3/X
+ sky130_fd_sc_hd__and4b_2
Xtap_34_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_29_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_10_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV SLICE\[1\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_19_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_19_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_1_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_23_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_23_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_6_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_6_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_25_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_27_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WEBUF\[5\] WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WEBUF\[5\]/X
+ sky130_fd_sc_hd__clkbuf_2
Xtap_21_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_18_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[0\] Do0_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF0\[56\]/Z
+ VGND VGND VPWR VPWR Do0[56] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_11_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[1\].FLOATBUF0\[12\] TIE0\[1\]/LO FBUFENBUF0\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_11_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_6_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_6_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_20_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.SEL1BUF SLICE\[1\].RAM8.DEC1.AND5/X VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[5\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_13_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[5\].FLOATBUF0\[43\] TIE0\[5\]/LO FBUFENBUF0\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[0\] BYTE\[2\].FLOATBUF1\[16\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_32_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_32_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_20_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_3_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_3_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_29_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_29_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo0_REG.OUTREG_BYTE\[4\].DIODE\[3\] BYTE\[4\].FLOATBUF0\[35\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV SLICE\[2\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[6\].DIODE\[7\] BYTE\[6\].FLOATBUF1\[55\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfill_9_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[1\] Do1_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF1\[9\]/Z
+ VGND VGND VPWR VPWR Do1[9] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_11_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDIBUF\[29\] Di0[29] VGND VGND VPWR VPWR DIBUF\[29\]/X sky130_fd_sc_hd__clkbuf_16
XDIODE_A1\[3\] A0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_27_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_27_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
Xfill_15_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_31_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[4\] Do0_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF0\[28\]/Z
+ VGND VGND VPWR VPWR Do0[28] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.DEC0.AND7 SLICE\[1\].RAM8.DEC0.AND7/A SLICE\[1\].RAM8.DEC0.AND7/B
+ SLICE\[1\].RAM8.DEC0.AND7/C SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_17_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.DEC1.ABUF\[0\] A1BUF\[0\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC1.AND7/A
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_7_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[1\].FLOATBUF0\[8\] TIE0\[1\]/LO FBUFENBUF0\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_13_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WEBUF\[2\] WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WEBUF\[2\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_31_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_0_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_17_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[7\] BYTE\[0\].FLOATBUF0\[7\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_9_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV SLICE\[2\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_28_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBYTE\[3\].FLOATBUF0\[24\] TIE0\[3\]/LO FBUFENBUF0\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[4\].FLOATBUF0\[39\] TIE0\[4\]/LO FBUFENBUF0\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XFBUFENBUF0\[3\] EN0 VGND VGND VPWR VPWR FBUFENBUF0\[3\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV SLICE\[1\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_5_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_12_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_12_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XA1BUF\[3\] A1[3] VGND VGND VPWR VPWR DEC1.AND3/B sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_8_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_14_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_30_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_9_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo1_REG.OUTREG_BYTE\[7\].DIODE\[0\] BYTE\[7\].FLOATBUF1\[56\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_30_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.DEC1.AND4 SLICE\[2\].RAM8.DEC1.AND7/A SLICE\[2\].RAM8.DEC1.AND7/B
+ SLICE\[2\].RAM8.DEC1.AND7/C SLICE\[2\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC1.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_34_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDIBUF\[11\] Di0[11] VGND VGND VPWR VPWR DIBUF\[11\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_10_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_19_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[0\].FLOATBUF1\[3\] TIE1\[0\]/LO FBUFENBUF1\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_1_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_23_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_6_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_6_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_20_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_25_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.SEL1BUF SLICE\[1\].RAM8.DEC1.AND4/X VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[4\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[6\].Do_FF\[1\] Do1_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF1\[49\]/Z
+ VGND VGND VPWR VPWR Do1[49] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV SLICE\[3\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XDIBUF\[59\] Di0[59] VGND VGND VPWR VPWR DIBUF\[59\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_27_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_21_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[0\] BYTE\[1\].FLOATBUF0\[8\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV SLICE\[2\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_18_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_33_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.Do_CLKBUF\[5\] Do1_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do1_REG.Do_CLKBUF\[5\]/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_11_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_6_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[4\] BYTE\[3\].FLOATBUF1\[28\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_20_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XTIE0\[5\] VGND VGND VPWR VPWR TIE0\[5\]/HI TIE0\[5\]/LO sky130_fd_sc_hd__conb_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_13_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[5\].DIODE\[7\] BYTE\[5\].FLOATBUF0\[47\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[1\] Do0_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF0\[1\]/Z
+ VGND VGND VPWR VPWR Do0[1] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_20_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_20_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_3_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_3_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_29_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[5\] Do1_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF1\[21\]/Z
+ VGND VGND VPWR VPWR Do1[21] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_9_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_11_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_27_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_27_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_15_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_31_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV SLICE\[2\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_17_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[41\] Di0[41] VGND VGND VPWR VPWR DIBUF\[41\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_7_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_31_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_17_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[7\].FLOATBUF1\[60\] TIE1\[7\]/LO FBUFENBUF1\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_9_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_28_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.DEC1.ABUF\[1\] A1BUF\[1\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC1.AND7/B
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[6\].DIODE\[0\] BYTE\[6\].FLOATBUF0\[48\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_24_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_5_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_12_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_12_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_22_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.SEL1BUF SLICE\[1\].RAM8.DEC1.AND3/X VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[3\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_14_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_30_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_30_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_9_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_9_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV SLICE\[3\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.DEC1.AND5 SLICE\[2\].RAM8.DEC1.AND7/B SLICE\[2\].RAM8.DEC1.AND7/A
+ SLICE\[2\].RAM8.DEC1.AND7/C SLICE\[2\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC1.AND5/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_29_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[1\] Do0_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF0\[41\]/Z
+ VGND VGND VPWR VPWR Do0[41] sky130_fd_sc_hd__dfxtp_1
XCLKBUF CLK VGND VGND VPWR VPWR CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_19_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV SLICE\[2\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_23_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_6_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[1\] BYTE\[0\].FLOATBUF1\[1\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[7\].Do_FF\[5\] Do1_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF1\[61\]/Z
+ VGND VGND VPWR VPWR Do1[61] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_20_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_6_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[1\].FLOATBUF1\[10\] TIE1\[1\]/LO FBUFENBUF1\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[4\] BYTE\[2\].FLOATBUF0\[20\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfill_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBYTE\[5\].FLOATBUF1\[41\] TIE1\[5\]/LO FBUFENBUF1\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.DEC1.ENBUF DEC1.AND3/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC1.AND7/D
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[4\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_18_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_18_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_33_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_11_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_6_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[5\] Do0_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF0\[13\]/Z
+ VGND VGND VPWR VPWR Do0[13] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_32_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_16_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_20_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_20_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_3_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_3_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV SLICE\[3\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_9_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_11_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_27_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_27_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_15_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_15_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_31_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_17_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDIBUF\[34\] Di0[34] VGND VGND VPWR VPWR DIBUF\[34\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_7_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[4\].FLOATBUF1\[37\] TIE1\[4\]/LO FBUFENBUF1\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[1\] Di0[1] VGND VGND VPWR VPWR DIBUF\[1\]/X sky130_fd_sc_hd__clkbuf_16
XDo1_REG.OUTREG_BYTE\[5\].DIODE\[1\] BYTE\[5\].FLOATBUF1\[41\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_24_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.SEL1BUF SLICE\[1\].RAM8.DEC1.AND2/X VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[2\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_26_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_9_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_9_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV SLICE\[3\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_28_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[7\].DIODE\[4\] BYTE\[7\].FLOATBUF0\[60\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV SLICE\[2\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WEBUF\[6\] WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WEBUF\[6\]/X
+ sky130_fd_sc_hd__clkbuf_2
Xtap_24_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_5_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[4\].Do_FF\[2\] Do1_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF1\[34\]/Z
+ VGND VGND VPWR VPWR Do1[34] sky130_fd_sc_hd__dfxtp_1
Xfill_12_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_22_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_14_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFBUFENBUF1\[6\] EN1 VGND VGND VPWR VPWR FBUFENBUF1\[6\]/X sky130_fd_sc_hd__clkbuf_2
Xtap_14_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_30_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_30_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[5\] Do0_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF0\[53\]/Z
+ VGND VGND VPWR VPWR Do0[53] sky130_fd_sc_hd__dfxtp_1
Xtap_34_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.DEC1.AND6 SLICE\[2\].RAM8.DEC1.AND7/A SLICE\[2\].RAM8.DEC1.AND7/B
+ SLICE\[2\].RAM8.DEC1.AND7/C SLICE\[2\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC1.AND6/X
+ sky130_fd_sc_hd__and4b_2
Xfill_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[7\].FLOATBUF0\[60\] TIE0\[7\]/LO FBUFENBUF0\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[7\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
Xtap_19_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[5\] BYTE\[1\].FLOATBUF1\[13\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_23_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_23_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_6_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_20_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_25_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_25_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_27_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_1_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.Do_CLKBUF\[7\] Do0_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do0_REG.Do_CLKBUF\[7\]/X
+ sky130_fd_sc_hd__clkbuf_4
XBYTE\[2\].FLOATBUF1\[18\] TIE1\[2\]/LO FBUFENBUF1\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[6\] Do1_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF1\[6\]/Z
+ VGND VGND VPWR VPWR Do1[6] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[6\].FLOATBUF1\[49\] TIE1\[6\]/LO FBUFENBUF1\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_18_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_18_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV SLICE\[3\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_33_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_11_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_11_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_32_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_18_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WEBUF\[3\] WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WEBUF\[3\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_20_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_3_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_29_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_22_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[1\].FLOATBUF0\[10\] TIE0\[1\]/LO FBUFENBUF0\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_9_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBYTE\[5\].FLOATBUF0\[41\] TIE0\[5\]/LO FBUFENBUF0\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.DEC0.ENBUF DEC0.AND3/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.AND7/D
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_27_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.SEL1BUF SLICE\[1\].RAM8.DEC1.AND1/X VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[1\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_15_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_15_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_31_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_31_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV SLICE\[3\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XDo0_REG.OUTREG_BYTE\[4\].DIODE\[1\] BYTE\[4\].FLOATBUF0\[33\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_17_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_17_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_33_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.DEC0.ABUF\[1\] A0BUF\[1\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.AND7/B
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[6\].DIODE\[5\] BYTE\[6\].FLOATBUF1\[53\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfill_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDIBUF\[27\] Di0[27] VGND VGND VPWR VPWR DIBUF\[27\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIODE_A1\[1\] A0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_26_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_9_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_9_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[2\] Do0_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF0\[26\]/Z
+ VGND VGND VPWR VPWR Do0[26] sky130_fd_sc_hd__dfxtp_1
Xtap_29_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[5\].Do_FF\[6\] Do1_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF1\[46\]/Z
+ VGND VGND VPWR VPWR Do1[46] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_4_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_5_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WEBUF\[0\] WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WEBUF\[0\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_22_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_8_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_14_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[5\] BYTE\[0\].FLOATBUF0\[5\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_30_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_30_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_34_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.DEC1.AND7 SLICE\[2\].RAM8.DEC1.AND7/A SLICE\[2\].RAM8.DEC1.AND7/B
+ SLICE\[2\].RAM8.DEC1.AND7/C SLICE\[2\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC1.AND7/X
+ sky130_fd_sc_hd__and4_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[4\].FLOATBUF0\[37\] TIE0\[4\]/LO FBUFENBUF0\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_29_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.DEC1.AND0 SLICE\[0\].RAM8.DEC1.AND7/A SLICE\[0\].RAM8.DEC1.AND7/B
+ SLICE\[0\].RAM8.DEC1.AND7/C SLICE\[0\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC1.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XFBUFENBUF0\[1\] EN0 VGND VGND VPWR VPWR FBUFENBUF0\[1\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV SLICE\[3\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_3_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_23_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_6_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_6_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XA1BUF\[1\] A1[1] VGND VGND VPWR VPWR A1BUF\[1\]/X sky130_fd_sc_hd__clkbuf_2
Xtap_6_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_20_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_25_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_27_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[0\].FLOATBUF1\[1\] TIE1\[0\]/LO FBUFENBUF1\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_18_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_33_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_11_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.SEL1BUF SLICE\[1\].RAM8.DEC1.AND0/Y VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[0\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[57\] Di0[57] VGND VGND VPWR VPWR DIBUF\[57\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_25_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_18_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.DEC1.ABUF\[2\] A1BUF\[2\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC1.AND7/C
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_3_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_3_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_29_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_22_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.Do_CLKBUF\[3\] Do1_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do1_REG.Do_CLKBUF\[3\]/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV SLICE\[0\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_10_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[2\].FLOATBUF0\[18\] TIE0\[2\]/LO FBUFENBUF0\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[2\] BYTE\[3\].FLOATBUF1\[26\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XTIE0\[3\] VGND VGND VPWR VPWR TIE0\[3\]/HI TIE0\[3\]/LO sky130_fd_sc_hd__conb_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_11_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[6\].FLOATBUF0\[49\] TIE0\[6\]/LO FBUFENBUF0\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_7_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_30_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_15_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[5\].DIODE\[5\] BYTE\[5\].FLOATBUF0\[45\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_31_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_31_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_17_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_33_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[3\] Do1_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF1\[19\]/Z
+ VGND VGND VPWR VPWR Do1[19] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_7_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[6\] Do0_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF0\[38\]/Z
+ VGND VGND VPWR VPWR Do0[38] sky130_fd_sc_hd__dfxtp_1
Xfill_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_26_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_9_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_9_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_28_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_4_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV SLICE\[3\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_5_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_22_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_8_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_14_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_14_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_14_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_14_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_30_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.DEC1.AND1 SLICE\[0\].RAM8.DEC1.AND7/C SLICE\[0\].RAM8.DEC1.AND7/B
+ SLICE\[0\].RAM8.DEC1.AND7/A SLICE\[0\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC1.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_3_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_23_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_6_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_6_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_20_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_25_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_13_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_27_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_1_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_1_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV SLICE\[0\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_11_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_11_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[7\].Do_FF\[3\] Do1_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF1\[59\]/Z
+ VGND VGND VPWR VPWR Do1[59] sky130_fd_sc_hd__dfxtp_1
Xtap_11_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_32_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XWEBUF\[7\] WE0[7] VGND VGND VPWR VPWR WEBUF\[7\]/X sky130_fd_sc_hd__clkbuf_2
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[2\] BYTE\[2\].FLOATBUF0\[18\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfill_25_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[2\].FLOATBUF1\[23\] TIE1\[2\]/LO FBUFENBUF1\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_18_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_3_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_3_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_29_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[6\].FLOATBUF1\[54\] TIE1\[6\]/LO FBUFENBUF1\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_29_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[4\].DIODE\[6\] BYTE\[4\].FLOATBUF1\[38\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_22_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_10_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.SEL1BUF SLICE\[0\].RAM8.DEC1.AND7/X VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[7\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_11_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_7_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_7_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WEBUF\[7\] WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[7\]/X
+ sky130_fd_sc_hd__clkbuf_2
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[3\] Do0_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF0\[11\]/Z
+ VGND VGND VPWR VPWR Do0[11] sky130_fd_sc_hd__dfxtp_1
Xfill_30_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_23_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_31_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_17_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_17_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[7\] Do1_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF1\[31\]/Z
+ VGND VGND VPWR VPWR Do1[31] sky130_fd_sc_hd__dfxtp_1
Xtap_33_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_33_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_7_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV SLICE\[0\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_0_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_26_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[0\].FLOATBUF0\[7\] TIE0\[0\]/LO FBUFENBUF0\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_4_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_4_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[32\] Di0[32] VGND VGND VPWR VPWR DIBUF\[32\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_5_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[4\].FLOATBUF1\[35\] TIE1\[4\]/LO FBUFENBUF1\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_22_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_8_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_14_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_14_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_30_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_34_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XDo0_REG.OUTREG_BYTE\[7\].DIODE\[2\] BYTE\[7\].FLOATBUF0\[58\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XBYTE\[1\].FLOATBUF1\[9\] TIE1\[1\]/LO FBUFENBUF1\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.DEC1.AND2 SLICE\[0\].RAM8.DEC1.AND7/C SLICE\[0\].RAM8.DEC1.AND7/A
+ SLICE\[0\].RAM8.DEC1.AND7/B SLICE\[0\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC1.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WEBUF\[4\] WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WEBUF\[4\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_3_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV SLICE\[0\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_6_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDo1_REG.OUTREG_BYTE\[4\].Do_FF\[0\] Do1_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF1\[32\]/Z
+ VGND VGND VPWR VPWR Do1[32] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_6_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_6_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_20_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_13_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_25_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_6_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_25_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XFBUFENBUF1\[4\] EN1 VGND VGND VPWR VPWR FBUFENBUF1\[4\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_13_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_13_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[3\] Do0_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF0\[51\]/Z
+ VGND VGND VPWR VPWR Do0[51] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_27_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_1_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.DEC0.ABUF\[2\] A0BUF\[2\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.AND7/C
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[3\] BYTE\[1\].FLOATBUF1\[11\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_33_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_33_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.SEL1BUF SLICE\[0\].RAM8.DEC1.AND6/X VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[6\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_11_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[6\] BYTE\[3\].FLOATBUF0\[30\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_32_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_25_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_18_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.Do_CLKBUF\[5\] Do0_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do0_REG.Do_CLKBUF\[5\]/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[2\].FLOATBUF1\[16\] TIE1\[2\]/LO FBUFENBUF1\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_3_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[4\] Do1_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF1\[4\]/Z
+ VGND VGND VPWR VPWR Do1[4] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_29_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_22_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_10_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_10_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV SLICE\[1\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[7\] Do0_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF0\[23\]/Z
+ VGND VGND VPWR VPWR Do0[23] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV SLICE\[0\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_7_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_7_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[62\] Di0[62] VGND VGND VPWR VPWR DIBUF\[62\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_30_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_23_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_16_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WEBUF\[1\] WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WEBUF\[1\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XTIE1\[6\] VGND VGND VPWR VPWR TIE1\[6\]/HI TIE1\[6\]/LO sky130_fd_sc_hd__conb_1
Xtap_33_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_21_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_21_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[2\].FLOATBUF0\[23\] TIE0\[2\]/LO FBUFENBUF0\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[6\].FLOATBUF0\[54\] TIE0\[6\]/LO FBUFENBUF0\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_9_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_29_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_28_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_16_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_16_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_32_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_4_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_4_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[6\].DIODE\[3\] BYTE\[6\].FLOATBUF1\[51\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfill_5_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[25\] Di0[25] VGND VGND VPWR VPWR DIBUF\[25\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV SLICE\[0\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_15_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_8_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_14_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_14_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[0\] Do0_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF0\[24\]/Z
+ VGND VGND VPWR VPWR Do0[24] sky130_fd_sc_hd__dfxtp_1
Xtap_34_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_27_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_1_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.DEC1.AND3 SLICE\[0\].RAM8.DEC1.AND7/C SLICE\[0\].RAM8.DEC1.AND7/B
+ SLICE\[0\].RAM8.DEC1.AND7/A SLICE\[0\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC1.AND3/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[5\].Do_FF\[4\] Do1_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF1\[44\]/Z
+ VGND VGND VPWR VPWR Do1[44] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_3_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_6_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_6_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.SEL1BUF SLICE\[0\].RAM8.DEC1.AND5/X VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[5\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_20_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[3\] BYTE\[0\].FLOATBUF0\[3\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[7\] Do0_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF0\[63\]/Z
+ VGND VGND VPWR VPWR Do0[63] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_13_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[4\].FLOATBUF0\[35\] TIE0\[4\]/LO FBUFENBUF0\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_27_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_1_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[7\] BYTE\[2\].FLOATBUF1\[23\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_1_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_33_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_11_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_11_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV SLICE\[1\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_11_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_4_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_24_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_24_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV SLICE\[0\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_32_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_25_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_18_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_3_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_3_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_10_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_19_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_7_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[55\] Di0[55] VGND VGND VPWR VPWR DIBUF\[55\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_30_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_16_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.DEC1.ABUF\[0\] A1BUF\[0\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC1.AND7/A
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_17_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_33_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.Do_CLKBUF\[1\] Do1_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do1_REG.Do_CLKBUF\[1\]/X
+ sky130_fd_sc_hd__clkbuf_4
Xfill_21_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_21_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_4_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[2\].FLOATBUF0\[16\] TIE0\[2\]/LO FBUFENBUF0\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[0\] BYTE\[3\].FLOATBUF1\[24\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XTIE0\[1\] VGND VGND VPWR VPWR TIE0\[1\]/HI TIE0\[1\]/LO sky130_fd_sc_hd__conb_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_0_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV SLICE\[1\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_9_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_9_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[5\].DIODE\[3\] BYTE\[5\].FLOATBUF0\[43\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_16_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_32_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[7\].DIODE\[7\] BYTE\[7\].FLOATBUF1\[63\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[1\] Do1_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF1\[17\]/Z
+ VGND VGND VPWR VPWR Do1[17] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_4_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_4_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[18\] Di0[18] VGND VGND VPWR VPWR DIBUF\[18\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.SEL1BUF SLICE\[0\].RAM8.DEC1.AND4/X VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[4\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_8_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[4\] Do0_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF0\[36\]/Z
+ VGND VGND VPWR VPWR Do0[36] sky130_fd_sc_hd__dfxtp_1
Xtap_14_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_30_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_27_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_1_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_27_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.DEC1.AND4 SLICE\[0\].RAM8.DEC1.AND7/A SLICE\[0\].RAM8.DEC1.AND7/B
+ SLICE\[0\].RAM8.DEC1.AND7/C SLICE\[0\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC1.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_3_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_6_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_6_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV SLICE\[1\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[7\] BYTE\[1\].FLOATBUF0\[15\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_20_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_13_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.DEC0.AND0 SLICE\[2\].RAM8.DEC0.AND7/A SLICE\[2\].RAM8.DEC0.AND7/B
+ SLICE\[2\].RAM8.DEC0.AND7/C SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
Xtap_6_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_13_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV SLICE\[0\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_1_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_1_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfill_33_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_11_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_11_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_24_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_24_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_7_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_32_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_25_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_18_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_3_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_3_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_22_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_10_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[7\].Do_FF\[1\] Do1_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF1\[57\]/Z
+ VGND VGND VPWR VPWR Do1[57] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_10_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_19_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_19_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV SLICE\[2\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_2_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_7_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_7_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV SLICE\[1\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XWEBUF\[5\] WE0[5] VGND VGND VPWR VPWR WEBUF\[5\]/X sky130_fd_sc_hd__clkbuf_2
Xfill_30_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[0\] BYTE\[2\].FLOATBUF0\[16\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfill_23_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[48\] Di0[48] VGND VGND VPWR VPWR DIBUF\[48\]/X sky130_fd_sc_hd__clkbuf_16
XBYTE\[2\].FLOATBUF1\[21\] TIE1\[2\]/LO FBUFENBUF1\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_16_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XBYTE\[6\].FLOATBUF1\[52\] TIE1\[6\]/LO FBUFENBUF1\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_17_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[4\].DIODE\[4\] BYTE\[4\].FLOATBUF1\[36\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_21_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_21_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_4_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.SEL1BUF SLICE\[0\].RAM8.DEC1.AND3/X VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[3\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XDo0_REG.OUTREG_BYTE\[6\].DIODE\[7\] BYTE\[6\].FLOATBUF0\[55\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WEBUF\[5\] WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[5\]/X
+ sky130_fd_sc_hd__clkbuf_2
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[1\] Do0_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF0\[9\]/Z
+ VGND VGND VPWR VPWR Do0[9] sky130_fd_sc_hd__dfxtp_1
Xtap_0_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_21_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_9_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_29_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[5\] Do1_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF1\[29\]/Z
+ VGND VGND VPWR VPWR Do1[29] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_16_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_32_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_32_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_4_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_4_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_5_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV SLICE\[1\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_14_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF SLICE\[3\].RAM8.DEC0.AND7/X VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_30_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_30_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_30_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_27_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[0\].FLOATBUF0\[5\] TIE0\[0\]/LO FBUFENBUF0\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_1_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_27_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_27_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.DEC1.AND5 SLICE\[0\].RAM8.DEC1.AND7/B SLICE\[0\].RAM8.DEC1.AND7/A
+ SLICE\[0\].RAM8.DEC1.AND7/C SLICE\[0\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC1.AND5/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_3_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[30\] Di0[30] VGND VGND VPWR VPWR DIBUF\[30\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_6_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[4\].FLOATBUF1\[33\] TIE1\[4\]/LO FBUFENBUF1\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_20_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_25_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.DEC0.AND1 SLICE\[2\].RAM8.DEC0.AND7/C SLICE\[2\].RAM8.DEC0.AND7/B
+ SLICE\[2\].RAM8.DEC0.AND7/A SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
Xtap_6_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_13_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_13_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[7\].DIODE\[0\] BYTE\[7\].FLOATBUF0\[56\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_1_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_1_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WEBUF\[2\] WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WEBUF\[2\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_1_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_11_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_33_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_11_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_11_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV SLICE\[2\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_4_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XFBUFENBUF1\[2\] EN1 VGND VGND VPWR VPWR FBUFENBUF1\[2\]/X sky130_fd_sc_hd__clkbuf_2
Xfill_24_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_24_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_24_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV SLICE\[1\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[1\] Do0_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF0\[49\]/Z
+ VGND VGND VPWR VPWR Do0[49] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_32_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_18_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.DEC0.ABUF\[0\] A0BUF\[0\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.AND7/A
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_3_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_3_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[1\] BYTE\[1\].FLOATBUF1\[9\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_10_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_10_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_19_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_19_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[4\] BYTE\[3\].FLOATBUF0\[28\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[2\].W.SEL1BUF SLICE\[0\].RAM8.DEC1.AND2/X VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[2\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_7_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_30_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_23_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XDo0_REG.Do_CLKBUF\[3\] Do0_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do0_REG.Do_CLKBUF\[3\]/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[3\].FLOATBUF1\[29\] TIE1\[3\]/LO FBUFENBUF1\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[8\] Di0[8] VGND VGND VPWR VPWR DIBUF\[8\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[2\] Do1_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF1\[2\]/Z
+ VGND VGND VPWR VPWR Do1[2] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_17_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_33_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_21_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_21_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[5\] Do0_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF0\[21\]/Z
+ VGND VGND VPWR VPWR Do0[21] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_0_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[60\] Di0[60] VGND VGND VPWR VPWR DIBUF\[60\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_21_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xtap_9_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF SLICE\[3\].RAM8.DEC0.AND6/X VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV SLICE\[2\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_16_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTIE1\[4\] VGND VGND VPWR VPWR TIE1\[4\]/HI TIE1\[4\]/LO sky130_fd_sc_hd__conb_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_16_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_32_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_32_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[2\].FLOATBUF0\[21\] TIE0\[2\]/LO FBUFENBUF0\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_4_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_4_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBYTE\[6\].FLOATBUF0\[52\] TIE0\[6\]/LO FBUFENBUF0\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_14_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_30_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_30_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_30_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_34_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_27_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_1_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_27_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_27_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDEC1.AND0 DEC1.AND3/B DEC1.AND3/A EN1BUF/X VGND VGND VPWR VPWR DEC1.AND0/Y sky130_fd_sc_hd__nor3b_2
XSLICE\[0\].RAM8.DEC1.AND6 SLICE\[0\].RAM8.DEC1.AND7/A SLICE\[0\].RAM8.DEC1.AND7/B
+ SLICE\[0\].RAM8.DEC1.AND7/C SLICE\[0\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC1.AND6/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[6\].DIODE\[1\] BYTE\[6\].FLOATBUF1\[49\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_3_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XDIBUF\[23\] Di0[23] VGND VGND VPWR VPWR DIBUF\[23\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_6_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_13_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV SLICE\[2\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_25_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.DEC0.AND2 SLICE\[2\].RAM8.DEC0.AND7/C SLICE\[2\].RAM8.DEC0.AND7/A
+ SLICE\[2\].RAM8.DEC0.AND7/B SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
Xtap_6_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_25_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XA0BUF\[3\] A0[3] VGND VGND VPWR VPWR DEC0.AND3/B sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_13_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV SLICE\[1\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_1_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[5\].Do_FF\[2\] Do1_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF1\[42\]/Z
+ VGND VGND VPWR VPWR Do1[42] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_1_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_11_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.CLKBUF CLKBUF/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.CLKBUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_11_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_4_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[1\] BYTE\[0\].FLOATBUF0\[1\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_24_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_24_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[5\] Do0_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF0\[61\]/Z
+ VGND VGND VPWR VPWR Do0[61] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.SEL1BUF SLICE\[0\].RAM8.DEC1.AND1/X VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[1\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_7_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_32_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBYTE\[4\].FLOATBUF0\[33\] TIE0\[4\]/LO FBUFENBUF0\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_25_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[5\] BYTE\[2\].FLOATBUF1\[21\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_3_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_10_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_19_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_19_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV SLICE\[3\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_12_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_7_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_7_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_30_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_23_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[6\] Do1_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF1\[14\]/Z
+ VGND VGND VPWR VPWR Do1[14] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF SLICE\[3\].RAM8.DEC0.AND5/X VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV SLICE\[2\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_16_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.DEC0.ABUF\[1\] A0BUF\[1\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.AND7/B
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_21_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_21_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_4_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_4_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[53\] Di0[53] VGND VGND VPWR VPWR DIBUF\[53\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_21_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.DEC1.ENBUF DEC1.AND1/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC1.AND7/D
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WEBUF\[7\] WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WEBUF\[7\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_29_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_28_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_16_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_16_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_32_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_32_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[3\].FLOATBUF0\[29\] TIE0\[3\]/LO FBUFENBUF0\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_4_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_34_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV SLICE\[2\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_14_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[5\].DIODE\[1\] BYTE\[5\].FLOATBUF0\[41\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_30_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_30_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_34_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_27_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_1_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_1_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_27_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.DEC1.AND7 SLICE\[0\].RAM8.DEC1.AND7/A SLICE\[0\].RAM8.DEC1.AND7/B
+ SLICE\[0\].RAM8.DEC1.AND7/C SLICE\[0\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC1.AND7/X
+ sky130_fd_sc_hd__and4_2
XDEC1.AND1 DEC1.AND3/A DEC1.AND3/B EN1BUF/X VGND VGND VPWR VPWR DEC1.AND1/X sky130_fd_sc_hd__and3b_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[7\].DIODE\[5\] BYTE\[7\].FLOATBUF1\[61\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_20_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_3_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[16\] Di0[16] VGND VGND VPWR VPWR DIBUF\[16\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_6_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_25_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.DEC0.AND3 SLICE\[2\].RAM8.DEC0.AND7/C SLICE\[2\].RAM8.DEC0.AND7/B
+ SLICE\[2\].RAM8.DEC0.AND7/A SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
Xtap_6_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[2\] Do0_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF0\[34\]/Z
+ VGND VGND VPWR VPWR Do0[34] sky130_fd_sc_hd__dfxtp_1
Xtap_25_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[0\].W.SEL1BUF SLICE\[0\].RAM8.DEC1.AND0/Y VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[0\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_13_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_13_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_25_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_1_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_15_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[6\].Do_FF\[6\] Do1_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF1\[54\]/Z
+ VGND VGND VPWR VPWR Do1[54] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_1_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_11_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[5\] BYTE\[1\].FLOATBUF0\[13\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_11_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_4_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV SLICE\[3\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_24_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_24_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.DEC1.ABUF\[2\] A1BUF\[2\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC1.AND7/C
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_7_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_25_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF SLICE\[3\].RAM8.DEC0.AND4/X VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_18_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV SLICE\[2\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_22_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_22_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[6\] Do0_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF0\[6\]/Z
+ VGND VGND VPWR VPWR Do0[6] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_10_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_19_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_19_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_2_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.DEC1.AND0 SLICE\[3\].RAM8.DEC1.AND7/A SLICE\[3\].RAM8.DEC1.AND7/B
+ SLICE\[3\].RAM8.DEC1.AND7/C SLICE\[3\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC1.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_12_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_7_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_23_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_16_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_17_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_33_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDIODE_A0\[3\] A0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_21_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_4_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_23_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XWEBUF\[3\] WE0[3] VGND VGND VPWR VPWR WEBUF\[3\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_21_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[46\] Di0[46] VGND VGND VPWR VPWR DIBUF\[46\]/X sky130_fd_sc_hd__clkbuf_16
Xtap_9_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV SLICE\[3\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_28_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBYTE\[6\].FLOATBUF1\[50\] TIE1\[6\]/LO FBUFENBUF1\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_16_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[4\].DIODE\[2\] BYTE\[4\].FLOATBUF1\[34\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_32_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_4_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[6\].DIODE\[5\] BYTE\[6\].FLOATBUF0\[53\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WEBUF\[3\] WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[3\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_14_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_30_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_27_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[3\] Do1_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF1\[27\]/Z
+ VGND VGND VPWR VPWR Do1[27] sky130_fd_sc_hd__dfxtp_1
Xfill_27_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_27_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDEC1.AND2 DEC1.AND3/B DEC1.AND3/A EN1BUF/X VGND VGND VPWR VPWR DEC1.AND2/X sky130_fd_sc_hd__and3b_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_20_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.DEC0.ENBUF DEC0.AND1/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.AND7/D
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_3_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[6\] Do0_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF0\[46\]/Z
+ VGND VGND VPWR VPWR Do0[46] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_25_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.DEC0.AND4 SLICE\[2\].RAM8.DEC0.AND7/A SLICE\[2\].RAM8.DEC0.AND7/B
+ SLICE\[2\].RAM8.DEC0.AND7/C SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_25_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV SLICE\[3\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_13_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[6\] BYTE\[0\].FLOATBUF1\[6\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_25_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[0\].FLOATBUF0\[3\] TIE0\[0\]/LO FBUFENBUF0\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_18_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF SLICE\[3\].RAM8.DEC0.AND3/X VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV SLICE\[2\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_1_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_15_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_15_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_31_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[1\].FLOATBUF1\[15\] TIE1\[1\]/LO FBUFENBUF1\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_1_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_33_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[5\].FLOATBUF1\[46\] TIE1\[5\]/LO FBUFENBUF1\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_11_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_4_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_24_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_30_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_26_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_18_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIODE_CLK CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WEBUF\[0\] WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WEBUF\[0\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_22_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_10_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_10_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_19_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_19_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_2_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XFBUFENBUF1\[0\] EN1 VGND VGND VPWR VPWR FBUFENBUF1\[0\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.DEC1.AND1 SLICE\[3\].RAM8.DEC1.AND7/C SLICE\[3\].RAM8.DEC1.AND7/B
+ SLICE\[3\].RAM8.DEC1.AND7/A SLICE\[3\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC1.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_12_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_7_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_30_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_16_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV SLICE\[3\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_17_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_33_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_33_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_21_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_21_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_4_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_23_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[2\] BYTE\[3\].FLOATBUF0\[26\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_21_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[39\] Di0[39] VGND VGND VPWR VPWR DIBUF\[39\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XDo0_REG.Do_CLKBUF\[1\] Do0_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do0_REG.Do_CLKBUF\[1\]/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[3\].FLOATBUF1\[27\] TIE1\[3\]/LO FBUFENBUF1\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[6\] Di0[6] VGND VGND VPWR VPWR DIBUF\[6\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[5\].DIODE\[6\] BYTE\[5\].FLOATBUF1\[46\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[0\] Do1_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF1\[0\]/Z
+ VGND VGND VPWR VPWR Do1[0] sky130_fd_sc_hd__dfxtp_1
Xtap_29_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XBYTE\[7\].FLOATBUF1\[58\] TIE1\[7\]/LO FBUFENBUF1\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_16_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_32_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_32_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_18_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_4_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
Xtap_34_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[3\] Do0_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF0\[19\]/Z
+ VGND VGND VPWR VPWR Do0[19] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV SLICE\[3\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_14_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_12_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_30_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[4\].Do_FF\[7\] Do1_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF1\[39\]/Z
+ VGND VGND VPWR VPWR Do1[39] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_27_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_1_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_1_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF SLICE\[3\].RAM8.DEC0.AND2/X VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XTIE1\[2\] VGND VGND VPWR VPWR TIE1\[2\]/HI TIE1\[2\]/LO sky130_fd_sc_hd__conb_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDEC1.AND3 DEC1.AND3/A DEC1.AND3/B EN1BUF/X VGND VGND VPWR VPWR DEC1.AND3/X sky130_fd_sc_hd__and3_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_20_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_33_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[6\].FLOATBUF0\[50\] TIE0\[6\]/LO FBUFENBUF0\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_25_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.DEC0.AND5 SLICE\[2\].RAM8.DEC0.AND7/B SLICE\[2\].RAM8.DEC0.AND7/A
+ SLICE\[2\].RAM8.DEC0.AND7/C SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
Xtap_25_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_13_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.DEC0.ABUF\[2\] A0BUF\[2\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.AND7/C
+ sky130_fd_sc_hd__clkbuf_2
Xtap_32_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_25_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_1_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_1_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_15_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_31_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_1_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[21\] Di0[21] VGND VGND VPWR VPWR DIBUF\[21\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_33_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_11_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_11_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XA0BUF\[1\] A0[1] VGND VGND VPWR VPWR A0BUF\[1\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_24_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_7_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_30_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_23_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_26_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV SLICE\[3\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XDo0_REG.Root_CLKBUF CLKBUF/X VGND VGND VPWR VPWR Do0_REG.Root_CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo1_REG.OUTREG_BYTE\[5\].Do_FF\[0\] Do1_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF1\[40\]/Z
+ VGND VGND VPWR VPWR Do1[40] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_10_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_10_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_19_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_2_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[3\] Do0_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF0\[59\]/Z
+ VGND VGND VPWR VPWR Do0[59] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.DEC1.AND2 SLICE\[3\].RAM8.DEC1.AND7/C SLICE\[3\].RAM8.DEC1.AND7/A
+ SLICE\[3\].RAM8.DEC1.AND7/B SLICE\[3\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC1.AND2/X
+ sky130_fd_sc_hd__and4bb_2
Xtap_12_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[1\].FLOATBUF0\[15\] TIE0\[1\]/LO FBUFENBUF0\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_7_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_7_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_23_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_16_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[5\].FLOATBUF0\[46\] TIE0\[5\]/LO FBUFENBUF0\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[3\] BYTE\[2\].FLOATBUF1\[19\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_17_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_33_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_21_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_21_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_4_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[7\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XDo0_REG.OUTREG_BYTE\[4\].DIODE\[6\] BYTE\[4\].FLOATBUF0\[38\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_0_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_23_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_21_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[4\] Do1_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF1\[12\]/Z
+ VGND VGND VPWR VPWR Do1[12] sky130_fd_sc_hd__dfxtp_1
Xfill_14_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV SLICE\[0\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF SLICE\[3\].RAM8.DEC0.AND1/X VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_16_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[7\] Do0_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF0\[31\]/Z
+ VGND VGND VPWR VPWR Do0[31] sky130_fd_sc_hd__dfxtp_1
Xtap_18_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[51\] Di0[51] VGND VGND VPWR VPWR DIBUF\[51\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_14_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_12_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_30_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WEBUF\[5\] WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WEBUF\[5\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_1_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_1_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_20_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_29_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[3\].FLOATBUF0\[27\] TIE0\[3\]/LO FBUFENBUF0\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XFBUFENBUF0\[6\] EN0 VGND VGND VPWR VPWR FBUFENBUF0\[6\]/X sky130_fd_sc_hd__clkbuf_2
Xfill_33_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[7\].FLOATBUF0\[58\] TIE0\[7\]/LO FBUFENBUF0\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_25_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.DEC0.AND6 SLICE\[2\].RAM8.DEC0.AND7/A SLICE\[2\].RAM8.DEC0.AND7/B
+ SLICE\[2\].RAM8.DEC0.AND7/C SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
Xtap_25_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_13_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_13_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_32_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_25_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_15_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_31_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV SLICE\[3\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[7\].DIODE\[3\] BYTE\[7\].FLOATBUF1\[59\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[14\] Di0[14] VGND VGND VPWR VPWR DIBUF\[14\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_33_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[0\].FLOATBUF1\[6\] TIE1\[0\]/LO FBUFENBUF1\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[0\] Do0_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF0\[32\]/Z
+ VGND VGND VPWR VPWR Do0[32] sky130_fd_sc_hd__dfxtp_1
Xfill_24_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_30_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XDo1_REG.OUTREG_BYTE\[6\].Do_FF\[4\] Do1_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF1\[52\]/Z
+ VGND VGND VPWR VPWR Do1[52] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_22_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_10_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[3\] BYTE\[1\].FLOATBUF0\[11\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_19_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.DEC1.AND3 SLICE\[3\].RAM8.DEC1.AND7/C SLICE\[3\].RAM8.DEC1.AND7/B
+ SLICE\[3\].RAM8.DEC1.AND7/A SLICE\[3\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC1.AND3/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.DEC1.ABUF\[0\] A1BUF\[0\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC1.AND7/A
+ sky130_fd_sc_hd__clkbuf_2
Xtap_12_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_12_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_7_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_7_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[7\] BYTE\[3\].FLOATBUF1\[31\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_16_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV SLICE\[0\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF SLICE\[3\].RAM8.DEC0.AND0/Y VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_33_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[4\] Do0_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF0\[4\]/Z
+ VGND VGND VPWR VPWR Do0[4] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_21_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_21_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_4_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_0_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_23_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_21_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_14_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_16_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_16_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_32_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIODE_A0\[1\] A0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_18_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_34_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XWEBUF\[1\] WE0[1] VGND VGND VPWR VPWR WEBUF\[1\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[44\] Di0[44] VGND VGND VPWR VPWR DIBUF\[44\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_12_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_30_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_34_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_1_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_1_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_27_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[7\].FLOATBUF1\[63\] TIE1\[7\]/LO FBUFENBUF1\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[4\].DIODE\[0\] BYTE\[4\].FLOATBUF1\[32\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_20_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV SLICE\[0\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[6\].DIODE\[3\] BYTE\[6\].FLOATBUF0\[51\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WEBUF\[1\] WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[1\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_25_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.DEC0.AND7 SLICE\[2\].RAM8.DEC0.AND7/A SLICE\[2\].RAM8.DEC0.AND7/B
+ SLICE\[2\].RAM8.DEC0.AND7/C SLICE\[2\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_8_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.DEC0.AND0 SLICE\[0\].RAM8.DEC0.AND7/A SLICE\[0\].RAM8.DEC0.AND7/B
+ SLICE\[0\].RAM8.DEC0.AND7/C SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_13_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_13_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[1\] Do1_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF1\[25\]/Z
+ VGND VGND VPWR VPWR Do1[25] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_31_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_1_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[4\] Do0_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF0\[44\]/Z
+ VGND VGND VPWR VPWR Do0[44] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_24_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_24_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_7_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[4\] BYTE\[0\].FLOATBUF1\[4\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_30_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
Xtap_23_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[0\].FLOATBUF0\[1\] TIE0\[0\]/LO FBUFENBUF0\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_26_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_26_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV SLICE\[0\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[1\].FLOATBUF1\[13\] TIE1\[1\]/LO FBUFENBUF1\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[7\] BYTE\[2\].FLOATBUF0\[23\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfill_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBYTE\[5\].FLOATBUF1\[44\] TIE1\[5\]/LO FBUFENBUF1\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_19_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.DEC1.AND4 SLICE\[3\].RAM8.DEC1.AND7/A SLICE\[3\].RAM8.DEC1.AND7/B
+ SLICE\[3\].RAM8.DEC1.AND7/C SLICE\[3\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC1.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_12_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_7_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_16_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_28_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_21_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_4_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_0_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_23_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF SLICE\[2\].RAM8.DEC0.AND7/X VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_14_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV SLICE\[1\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_32_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV SLICE\[0\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_34_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_34_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[0\] BYTE\[3\].FLOATBUF0\[24\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[37\] Di0[37] VGND VGND VPWR VPWR DIBUF\[37\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[3\].FLOATBUF1\[25\] TIE1\[3\]/LO FBUFENBUF1\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[4\] Di0[4] VGND VGND VPWR VPWR DIBUF\[4\]/X sky130_fd_sc_hd__clkbuf_16
XDo1_REG.OUTREG_BYTE\[5\].DIODE\[4\] BYTE\[5\].FLOATBUF1\[44\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_27_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[7\].FLOATBUF1\[56\] TIE1\[7\]/LO FBUFENBUF1\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_20_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_20_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[7\].DIODE\[7\] BYTE\[7\].FLOATBUF0\[63\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[1\] Do0_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF0\[17\]/Z
+ VGND VGND VPWR VPWR Do0[17] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_8_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.DEC0.AND1 SLICE\[0\].RAM8.DEC0.AND7/C SLICE\[0\].RAM8.DEC0.AND7/B
+ SLICE\[0\].RAM8.DEC0.AND7/A SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_13_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[4\].Do_FF\[5\] Do1_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF1\[37\]/Z
+ VGND VGND VPWR VPWR Do1[37] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_25_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[5\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_18_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTIE1\[0\] VGND VGND VPWR VPWR TIE1\[0\]/HI TIE1\[0\]/LO sky130_fd_sc_hd__conb_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_31_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV SLICE\[0\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_0_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_1_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[7\].FLOATBUF0\[63\] TIE0\[7\]/LO FBUFENBUF0\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_24_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_7_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.DEC0.ABUF\[0\] A0BUF\[0\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.AND7/A
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_30_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_23_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_16_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_26_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_2_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_2_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_19_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_19_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.DEC1.AND5 SLICE\[3\].RAM8.DEC1.AND7/B SLICE\[3\].RAM8.DEC1.AND7/A
+ SLICE\[3\].RAM8.DEC1.AND7/C SLICE\[3\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC1.AND5/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_12_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_12_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF SLICE\[2\].RAM8.DEC0.AND6/X VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_21_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV SLICE\[1\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_28_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WEBUF\[6\] WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WEBUF\[6\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_21_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_4_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV SLICE\[0\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_23_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[1\] Do0_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF0\[57\]/Z
+ VGND VGND VPWR VPWR Do0[57] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBYTE\[1\].FLOATBUF0\[13\] TIE0\[1\]/LO FBUFENBUF0\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_21_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBYTE\[5\].FLOATBUF0\[44\] TIE0\[5\]/LO FBUFENBUF0\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[1\] BYTE\[2\].FLOATBUF1\[17\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_16_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_32_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[4\].DIODE\[4\] BYTE\[4\].FLOATBUF0\[36\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_18_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[2\] Do1_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF1\[10\]/Z
+ VGND VGND VPWR VPWR Do1[10] sky130_fd_sc_hd__dfxtp_1
Xfill_12_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIODE_A1\[4\] A0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[6\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_1_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_27_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_20_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_20_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_20_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_20_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[5\] Do0_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF0\[29\]/Z
+ VGND VGND VPWR VPWR Do0[29] sky130_fd_sc_hd__dfxtp_1
Xtap_29_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_29_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.DEC1.ABUF\[1\] A1BUF\[1\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC1.AND7/B
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV SLICE\[1\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_33_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_33_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_5_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_5_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfill_10_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XBYTE\[1\].FLOATBUF0\[9\] TIE0\[1\]/LO FBUFENBUF0\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.DEC0.AND2 SLICE\[0\].RAM8.DEC0.AND7/C SLICE\[0\].RAM8.DEC0.AND7/A
+ SLICE\[0\].RAM8.DEC0.AND7/B SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WEBUF\[3\] WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WEBUF\[3\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_25_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_15_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_31_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_31_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfill_0_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[3\].FLOATBUF0\[25\] TIE0\[3\]/LO FBUFENBUF0\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XFBUFENBUF0\[4\] EN0 VGND VGND VPWR VPWR FBUFENBUF0\[4\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XBYTE\[7\].FLOATBUF0\[56\] TIE0\[7\]/LO FBUFENBUF0\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_6_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_7_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XA1BUF\[4\] A1[4] VGND VGND VPWR VPWR DEC1.AND3/A sky130_fd_sc_hd__clkbuf_2
Xtap_30_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF SLICE\[2\].RAM8.DEC0.AND5/X VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_14_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[7\].DIODE\[1\] BYTE\[7\].FLOATBUF1\[57\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV SLICE\[1\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_2_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_2_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[1\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[12\] Di0[12] VGND VGND VPWR VPWR DIBUF\[12\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[0\].FLOATBUF1\[4\] TIE1\[0\]/LO FBUFENBUF1\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_19_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV SLICE\[0\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_2_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.DEC1.AND6 SLICE\[3\].RAM8.DEC1.AND7/A SLICE\[3\].RAM8.DEC1.AND7/B
+ SLICE\[3\].RAM8.DEC1.AND7/C SLICE\[3\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC1.AND6/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_12_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_12_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_14_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[6\].Do_FF\[2\] Do1_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF1\[50\]/Z
+ VGND VGND VPWR VPWR Do1[50] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_28_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[1\] BYTE\[1\].FLOATBUF0\[9\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_4_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_23_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_23_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.Do_CLKBUF\[6\] Do1_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do1_REG.Do_CLKBUF\[6\]/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_11_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[5\] BYTE\[3\].FLOATBUF1\[29\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XTIE0\[6\] VGND VGND VPWR VPWR TIE0\[6\]/HI TIE0\[6\]/LO sky130_fd_sc_hd__conb_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_14_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_8_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_8_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_32_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV SLICE\[2\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[2\] Do0_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF0\[2\]/Z
+ VGND VGND VPWR VPWR Do0[2] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_34_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV SLICE\[1\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_22_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[6\] Do1_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF1\[22\]/Z
+ VGND VGND VPWR VPWR Do1[22] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_12_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_1_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_27_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_20_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_20_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_29_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_17_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_5_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_5_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_5_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDIBUF\[42\] Di0[42] VGND VGND VPWR VPWR DIBUF\[42\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_8_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_10_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.DEC0.AND3 SLICE\[0\].RAM8.DEC0.AND7/C SLICE\[0\].RAM8.DEC0.AND7/B
+ SLICE\[0\].RAM8.DEC0.AND7/A SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[3\].FLOATBUF1\[30\] TIE1\[3\]/LO FBUFENBUF1\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_32_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF SLICE\[2\].RAM8.DEC0.AND4/X VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_25_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[7\].FLOATBUF1\[61\] TIE1\[7\]/LO FBUFENBUF1\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_31_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_31_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_31_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_0_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV SLICE\[1\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.DEC1.ABUF\[2\] A1BUF\[2\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC1.AND7/C
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[6\].DIODE\[1\] BYTE\[6\].FLOATBUF0\[49\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_6_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_7_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_30_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_26_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_26_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_14_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_14_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_2_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_2_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[2\] Do0_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF0\[42\]/Z
+ VGND VGND VPWR VPWR Do0[42] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_12_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.DEC1.AND7 SLICE\[3\].RAM8.DEC1.AND7/A SLICE\[3\].RAM8.DEC1.AND7/B
+ SLICE\[3\].RAM8.DEC1.AND7/C SLICE\[3\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC1.AND7/X
+ sky130_fd_sc_hd__and4_2
Xtap_12_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_12_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[2\] BYTE\[0\].FLOATBUF1\[2\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.DEC1.AND0 SLICE\[1\].RAM8.DEC1.AND7/A SLICE\[1\].RAM8.DEC1.AND7/B
+ SLICE\[1\].RAM8.DEC1.AND7/C SLICE\[1\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC1.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XDo1_REG.OUTREG_BYTE\[7\].Do_FF\[6\] Do1_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF1\[62\]/Z
+ VGND VGND VPWR VPWR Do1[62] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_14_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_25_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[1\].FLOATBUF1\[11\] TIE1\[1\]/LO FBUFENBUF1\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[5\] BYTE\[2\].FLOATBUF0\[21\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV SLICE\[2\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[5\].FLOATBUF1\[42\] TIE1\[5\]/LO FBUFENBUF1\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_0_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV SLICE\[1\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_23_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_23_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_11_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_11_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_14_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_8_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[6\] Do0_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF0\[14\]/Z
+ VGND VGND VPWR VPWR Do0[14] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_26_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_18_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_34_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_22_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_22_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_12_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF SLICE\[2\].RAM8.DEC0.AND3/X VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_1_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_1_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_20_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_20_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_29_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_17_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_17_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV SLICE\[2\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_5_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_5_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_5_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[35\] Di0[35] VGND VGND VPWR VPWR DIBUF\[35\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_8_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.DEC0.AND4 SLICE\[0\].RAM8.DEC0.AND7/A SLICE\[0\].RAM8.DEC0.AND7/B
+ SLICE\[0\].RAM8.DEC0.AND7/C SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[4\].FLOATBUF1\[38\] TIE1\[4\]/LO FBUFENBUF1\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[2\] Di0[2] VGND VGND VPWR VPWR DIBUF\[2\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[5\].DIODE\[2\] BYTE\[5\].FLOATBUF1\[42\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_25_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_18_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_15_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_31_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_31_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_31_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[7\].DIODE\[5\] BYTE\[7\].FLOATBUF0\[61\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WEBUF\[7\] WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WEBUF\[7\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_6_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[4\].Do_FF\[3\] Do1_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF1\[35\]/Z
+ VGND VGND VPWR VPWR Do1[35] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_30_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XFBUFENBUF1\[7\] EN1 VGND VGND VPWR VPWR FBUFENBUF1\[7\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_14_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_14_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_30_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_30_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[3\].FLOATBUF0\[30\] TIE0\[3\]/LO FBUFENBUF0\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[6\] Do0_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF0\[54\]/Z
+ VGND VGND VPWR VPWR Do0[54] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
Xfill_2_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_2_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV SLICE\[2\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[7\].FLOATBUF0\[61\] TIE0\[7\]/LO FBUFENBUF0\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[6\] BYTE\[1\].FLOATBUF1\[14\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV SLICE\[1\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_12_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_12_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.DEC1.AND1 SLICE\[1\].RAM8.DEC1.AND7/C SLICE\[1\].RAM8.DEC1.AND7/B
+ SLICE\[1\].RAM8.DEC1.AND7/A SLICE\[1\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC1.AND1/X
+ sky130_fd_sc_hd__and4bb_2
Xtap_21_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_14_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_25_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_28_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[2\].FLOATBUF1\[19\] TIE1\[2\]/LO FBUFENBUF1\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[7\] Do1_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF1\[7\]/Z
+ VGND VGND VPWR VPWR Do1[7] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_23_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.CLKBUF CLKBUF/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.CLKBUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_11_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF SLICE\[2\].RAM8.DEC0.AND2/X VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_8_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_8_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_26_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_19_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WEBUF\[4\] WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WEBUF\[4\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV SLICE\[3\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_18_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_18_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_34_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_34_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_22_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_22_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV SLICE\[2\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XBYTE\[1\].FLOATBUF0\[11\] TIE0\[1\]/LO FBUFENBUF0\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_5_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBYTE\[5\].FLOATBUF0\[42\] TIE0\[5\]/LO FBUFENBUF0\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_1_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_1_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_20_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_29_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[4\].DIODE\[2\] BYTE\[4\].FLOATBUF0\[34\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_17_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_17_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.DEC0.ABUF\[2\] A0BUF\[2\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.AND7/C
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_5_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[6\].DIODE\[6\] BYTE\[6\].FLOATBUF1\[54\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfill_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[0\] Do1_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF1\[8\]/Z
+ VGND VGND VPWR VPWR Do1[8] sky130_fd_sc_hd__dfxtp_1
Xfill_10_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[28\] Di0[28] VGND VGND VPWR VPWR DIBUF\[28\]/X sky130_fd_sc_hd__clkbuf_16
XDIODE_A1\[2\] A0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.DEC0.AND5 SLICE\[0\].RAM8.DEC0.AND7/B SLICE\[0\].RAM8.DEC0.AND7/A
+ SLICE\[0\].RAM8.DEC0.AND7/C SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_18_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_15_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_15_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_31_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[3\] Do0_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF0\[27\]/Z
+ VGND VGND VPWR VPWR Do0[27] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_2_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_2_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
Xfill_28_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV SLICE\[2\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.Root_CLKBUF CLKBUF/X VGND VGND VPWR VPWR Do1_REG.Root_CLKBUF/X sky130_fd_sc_hd__clkbuf_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[5\].Do_FF\[7\] Do1_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF1\[47\]/Z
+ VGND VGND VPWR VPWR Do1[47] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_7_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WEBUF\[1\] WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WEBUF\[1\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_30_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_23_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_16_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[6\] BYTE\[0\].FLOATBUF0\[6\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_14_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_30_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_30_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_2_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_2_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBYTE\[4\].FLOATBUF0\[38\] TIE0\[4\]/LO FBUFENBUF0\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XFBUFENBUF0\[2\] EN0 VGND VGND VPWR VPWR FBUFENBUF0\[2\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_4_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_12_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_12_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XA1BUF\[2\] A1[2] VGND VGND VPWR VPWR A1BUF\[2\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.DEC1.AND2 SLICE\[1\].RAM8.DEC1.AND7/C SLICE\[1\].RAM8.DEC1.AND7/A
+ SLICE\[1\].RAM8.DEC1.AND7/B SLICE\[1\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC1.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_21_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_14_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_7_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_25_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_8_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF SLICE\[2\].RAM8.DEC0.AND1/X VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_28_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[10\] Di0[10] VGND VGND VPWR VPWR DIBUF\[10\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV SLICE\[3\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_4_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[0\].FLOATBUF1\[2\] TIE1\[0\]/LO FBUFENBUF1\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_0_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_23_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV SLICE\[2\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_11_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_12_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[6\].Do_FF\[0\] Do1_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF1\[48\]/Z
+ VGND VGND VPWR VPWR Do1[48] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_8_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_8_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[58\] Di0[58] VGND VGND VPWR VPWR DIBUF\[58\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_33_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_26_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_18_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_34_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.Do_CLKBUF\[4\] Do1_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do1_REG.Do_CLKBUF\[4\]/X
+ sky130_fd_sc_hd__clkbuf_4
Xfill_22_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_22_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_5_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[2\].FLOATBUF0\[19\] TIE0\[2\]/LO FBUFENBUF0\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[3\] BYTE\[3\].FLOATBUF1\[27\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTIE0\[4\] VGND VGND VPWR VPWR TIE0\[4\]/HI TIE0\[4\]/LO sky130_fd_sc_hd__conb_1
Xfill_12_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_1_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_1_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_31_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[5\].DIODE\[6\] BYTE\[5\].FLOATBUF0\[46\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[0\] Do0_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF0\[0\]/Z
+ VGND VGND VPWR VPWR Do0[0] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_20_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_20_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_29_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_17_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_33_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[6\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[4\] Do1_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF1\[20\]/Z
+ VGND VGND VPWR VPWR Do1[20] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_5_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_5_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV SLICE\[3\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_8_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDEC0.AND0 DEC0.AND3/B DEC0.AND3/A EN0BUF/X VGND VGND VPWR VPWR DEC0.AND0/Y sky130_fd_sc_hd__nor3b_2
XSLICE\[0\].RAM8.DEC0.AND6 SLICE\[0\].RAM8.DEC0.AND7/A SLICE\[0\].RAM8.DEC0.AND7/B
+ SLICE\[0\].RAM8.DEC0.AND7/C SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_15_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[7\] Do0_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF0\[39\]/Z
+ VGND VGND VPWR VPWR Do0[39] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.SEL1BUF SLICE\[3\].RAM8.DEC1.AND7/X VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[7\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_31_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_2_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_28_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_28_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[40\] Di0[40] VGND VGND VPWR VPWR DIBUF\[40\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_6_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_7_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_23_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_16_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_26_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_26_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_14_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_14_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF SLICE\[2\].RAM8.DEC0.AND0/Y VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_30_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_30_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_30_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_2_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.DEC1.ABUF\[0\] A1BUF\[0\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC1.AND7/A
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV SLICE\[3\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_4_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_12_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_12_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV SLICE\[2\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.DEC1.AND3 SLICE\[1\].RAM8.DEC1.AND7/C SLICE\[1\].RAM8.DEC1.AND7/B
+ SLICE\[1\].RAM8.DEC1.AND7/A SLICE\[1\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC1.AND3/X
+ sky130_fd_sc_hd__and4b_2
Xtap_21_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_14_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_25_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_8_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_28_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[0\] Do0_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF0\[40\]/Z
+ VGND VGND VPWR VPWR Do0[40] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_4_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_23_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_23_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_11_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_11_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[0\] BYTE\[0\].FLOATBUF1\[0\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XDo1_REG.OUTREG_BYTE\[7\].Do_FF\[4\] Do1_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF1\[60\]/Z
+ VGND VGND VPWR VPWR Do1[60] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_12_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_5_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_8_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_8_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[3\] BYTE\[2\].FLOATBUF0\[19\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfill_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_19_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[5\].FLOATBUF1\[40\] TIE1\[5\]/LO FBUFENBUF1\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV SLICE\[0\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XBYTE\[6\].FLOATBUF1\[55\] TIE1\[6\]/LO FBUFENBUF1\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[4\].DIODE\[7\] BYTE\[4\].FLOATBUF1\[39\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_22_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_22_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV SLICE\[3\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_12_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_1_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[4\] Do0_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF0\[12\]/Z
+ VGND VGND VPWR VPWR Do0[12] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_31_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_24_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[6\].W.SEL1BUF SLICE\[3\].RAM8.DEC1.AND6/X VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[6\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_20_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_29_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_17_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_33_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_33_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_5_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_8_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_10_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDEC0.AND1 DEC0.AND3/A DEC0.AND3/B EN0BUF/X VGND VGND VPWR VPWR DEC0.AND1/X sky130_fd_sc_hd__and3b_2
XSLICE\[0\].RAM8.DEC0.AND7 SLICE\[0\].RAM8.DEC0.AND7/A SLICE\[0\].RAM8.DEC0.AND7/B
+ SLICE\[0\].RAM8.DEC0.AND7/C SLICE\[0\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_15_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_31_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_0_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_2_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_28_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_28_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV SLICE\[3\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[33\] Di0[33] VGND VGND VPWR VPWR DIBUF\[33\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_6_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_7_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_7_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[4\].FLOATBUF1\[36\] TIE1\[4\]/LO FBUFENBUF1\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[5\].DIODE\[0\] BYTE\[5\].FLOATBUF1\[40\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XDIBUF\[0\] Di0[0] VGND VGND VPWR VPWR DIBUF\[0\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_23_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_26_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_9_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_14_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_14_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_30_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_30_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_30_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_2_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[7\].DIODE\[3\] BYTE\[7\].FLOATBUF0\[59\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WEBUF\[5\] WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WEBUF\[5\]/X
+ sky130_fd_sc_hd__clkbuf_2
Xfill_4_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_12_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF SLICE\[1\].RAM8.DEC0.AND7/X VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XDo1_REG.OUTREG_BYTE\[4\].Do_FF\[1\] Do1_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF1\[33\]/Z
+ VGND VGND VPWR VPWR Do1[33] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.DEC1.AND4 SLICE\[1\].RAM8.DEC1.AND7/A SLICE\[1\].RAM8.DEC1.AND7/B
+ SLICE\[1\].RAM8.DEC1.AND7/C SLICE\[1\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC1.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_21_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_14_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_7_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_25_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFBUFENBUF1\[5\] EN1 VGND VGND VPWR VPWR FBUFENBUF1\[5\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_8_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_8_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[4\] Do0_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF0\[52\]/Z
+ VGND VGND VPWR VPWR Do0[52] sky130_fd_sc_hd__dfxtp_1
Xfill_28_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.DEC0.AND0 SLICE\[3\].RAM8.DEC0.AND7/A SLICE\[3\].RAM8.DEC0.AND7/B
+ SLICE\[3\].RAM8.DEC0.AND7/C SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_4_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV SLICE\[0\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[4\] BYTE\[1\].FLOATBUF1\[12\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_23_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_23_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
Xfill_11_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_11_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV SLICE\[3\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_12_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_5_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[7\] BYTE\[3\].FLOATBUF0\[31\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_8_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_8_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_33_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_26_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.SEL1BUF SLICE\[3\].RAM8.DEC1.AND5/X VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[5\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_19_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.Do_CLKBUF\[6\] Do0_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do0_REG.Do_CLKBUF\[6\]/X
+ sky130_fd_sc_hd__clkbuf_4
XBYTE\[2\].FLOATBUF1\[17\] TIE1\[2\]/LO FBUFENBUF1\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[5\] Do1_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF1\[5\]/Z
+ VGND VGND VPWR VPWR Do1[5] sky130_fd_sc_hd__dfxtp_1
Xtap_18_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[6\].FLOATBUF1\[48\] TIE1\[6\]/LO FBUFENBUF1\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_34_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfill_22_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_22_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_5_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XDIBUF\[63\] Di0[63] VGND VGND VPWR VPWR DIBUF\[63\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_31_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_17_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WEBUF\[2\] WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WEBUF\[2\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_20_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_20_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_29_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_17_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTIE1\[7\] VGND VGND VPWR VPWR TIE1\[7\]/HI TIE1\[7\]/LO sky130_fd_sc_hd__conb_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_33_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_10_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_5_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV SLICE\[0\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDEC0.AND2 DEC0.AND3/B DEC0.AND3/A EN0BUF/X VGND VGND VPWR VPWR DEC0.AND2/X sky130_fd_sc_hd__and3b_2
XBYTE\[5\].FLOATBUF0\[40\] TIE0\[5\]/LO FBUFENBUF0\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XBYTE\[6\].FLOATBUF0\[55\] TIE0\[6\]/LO FBUFENBUF0\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_15_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_31_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_2_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_2_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[4\].DIODE\[0\] BYTE\[4\].FLOATBUF0\[32\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfill_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_28_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.DEC0.ABUF\[0\] A0BUF\[0\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.AND7/A
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[6\].DIODE\[4\] BYTE\[6\].FLOATBUF1\[52\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_6_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[26\] Di0[26] VGND VGND VPWR VPWR DIBUF\[26\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XDIODE_A1\[0\] A0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_7_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF SLICE\[1\].RAM8.DEC0.AND6/X VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_26_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_26_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_9_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_14_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_30_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[1\] Do0_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF0\[25\]/Z
+ VGND VGND VPWR VPWR Do0[25] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_2_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_16_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV SLICE\[0\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[5\].Do_FF\[5\] Do1_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF1\[45\]/Z
+ VGND VGND VPWR VPWR Do1[45] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_4_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_12_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
Xtap_12_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.DEC1.AND5 SLICE\[1\].RAM8.DEC1.AND7/B SLICE\[1\].RAM8.DEC1.AND7/A
+ SLICE\[1\].RAM8.DEC1.AND7/C SLICE\[1\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC1.AND5/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV SLICE\[3\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_21_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_25_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[4\] BYTE\[0\].FLOATBUF0\[4\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_8_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_8_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.CLKBUF CLKBUF/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.CLKBUF/X sky130_fd_sc_hd__clkbuf_2
XBYTE\[4\].FLOATBUF0\[36\] TIE0\[4\]/LO FBUFENBUF0\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.SEL1BUF SLICE\[3\].RAM8.DEC1.AND4/X VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[4\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_28_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XFBUFENBUF0\[0\] EN0 VGND VGND VPWR VPWR FBUFENBUF0\[0\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.DEC0.AND1 SLICE\[3\].RAM8.DEC0.AND7/C SLICE\[3\].RAM8.DEC0.AND7/B
+ SLICE\[3\].RAM8.DEC0.AND7/A SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_23_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XA1BUF\[0\] A1[0] VGND VGND VPWR VPWR A1BUF\[0\]/X sky130_fd_sc_hd__clkbuf_2
Xfill_11_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XEN0BUF EN0 VGND VGND VPWR VPWR EN0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_11_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_12_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_5_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_8_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_19_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_18_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[0\].FLOATBUF1\[0\] TIE1\[0\]/LO FBUFENBUF1\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_18_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV SLICE\[1\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_34_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_22_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_5_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_5_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV SLICE\[0\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[56\] Di0[56] VGND VGND VPWR VPWR DIBUF\[56\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_24_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfill_17_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.DEC1.ABUF\[1\] A1BUF\[1\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC1.AND7/B
+ sky130_fd_sc_hd__clkbuf_2
Xfill_0_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_20_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_17_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo1_REG.Do_CLKBUF\[2\] Do1_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do1_REG.Do_CLKBUF\[2\]/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_10_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[2\].FLOATBUF0\[17\] TIE0\[2\]/LO FBUFENBUF0\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_5_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[1\] BYTE\[3\].FLOATBUF1\[25\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_19_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_5_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XTIE0\[2\] VGND VGND VPWR VPWR TIE0\[2\]/HI TIE0\[2\]/LO sky130_fd_sc_hd__conb_1
Xfill_10_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF SLICE\[1\].RAM8.DEC0.AND5/X VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XDEC0.AND3 DEC0.AND3/A DEC0.AND3/B EN0BUF/X VGND VGND VPWR VPWR DEC0.AND3/X sky130_fd_sc_hd__and3_2
XBYTE\[6\].FLOATBUF0\[48\] TIE0\[6\]/LO FBUFENBUF0\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_15_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_31_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[5\].DIODE\[4\] BYTE\[5\].FLOATBUF0\[44\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_31_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_2_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_28_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[2\] Do1_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF1\[18\]/Z
+ VGND VGND VPWR VPWR Do1[18] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV SLICE\[0\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[19\] Di0[19] VGND VGND VPWR VPWR DIBUF\[19\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_26_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
Xtap_9_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[5\] Do0_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF0\[37\]/Z
+ VGND VGND VPWR VPWR Do0[37] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_14_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_30_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_28_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.SEL1BUF SLICE\[3\].RAM8.DEC1.AND3/X VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[3\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_2_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_2_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_16_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_4_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.DEC1.ENBUF DEC1.AND2/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC1.AND7/D
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.DEC1.AND6 SLICE\[1\].RAM8.DEC1.AND7/A SLICE\[1\].RAM8.DEC1.AND7/B
+ SLICE\[1\].RAM8.DEC1.AND7/C SLICE\[1\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC1.AND6/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_25_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_25_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_8_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_8_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_27_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_28_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.DEC0.AND2 SLICE\[3\].RAM8.DEC0.AND7/C SLICE\[3\].RAM8.DEC0.AND7/A
+ SLICE\[3\].RAM8.DEC0.AND7/B SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV SLICE\[1\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_23_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_23_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_11_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_11_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_12_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV SLICE\[0\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_5_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_13_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_8_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_26_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_19_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_34_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_22_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_5_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_5_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[7\].Do_FF\[2\] Do1_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF1\[58\]/Z
+ VGND VGND VPWR VPWR Do1[58] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF SLICE\[1\].RAM8.DEC0.AND4/X VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_24_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_31_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XWEBUF\[6\] WE0[6] VGND VGND VPWR VPWR WEBUF\[6\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[1\] BYTE\[2\].FLOATBUF0\[17\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_24_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[49\] Di0[49] VGND VGND VPWR VPWR DIBUF\[49\]/X sky130_fd_sc_hd__clkbuf_16
XBYTE\[2\].FLOATBUF1\[22\] TIE1\[2\]/LO FBUFENBUF1\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_17_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_20_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_29_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_29_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[6\].FLOATBUF1\[53\] TIE1\[6\]/LO FBUFENBUF1\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_17_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_17_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDo1_REG.OUTREG_BYTE\[4\].DIODE\[5\] BYTE\[4\].FLOATBUF1\[37\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfill_33_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_10_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_10_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_5_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_19_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_10_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV SLICE\[1\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WEBUF\[6\] WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[6\]/X
+ sky130_fd_sc_hd__clkbuf_2
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[2\] Do0_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF0\[10\]/Z
+ VGND VGND VPWR VPWR Do0[10] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_22_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_2_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_28_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_28_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.SEL1BUF SLICE\[3\].RAM8.DEC1.AND2/X VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[2\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[6\] Do1_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF1\[30\]/Z
+ VGND VGND VPWR VPWR Do1[30] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_21_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_6_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_26_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_14_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_14_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_30_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[0\].FLOATBUF0\[6\] TIE0\[0\]/LO FBUFENBUF0\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_2_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_16_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_32_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV SLICE\[1\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[31\] Di0[31] VGND VGND VPWR VPWR DIBUF\[31\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_4_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[4\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_12_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[4\].FLOATBUF1\[34\] TIE1\[4\]/LO FBUFENBUF1\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.DEC1.AND7 SLICE\[1\].RAM8.DEC1.AND7/A SLICE\[1\].RAM8.DEC1.AND7/B
+ SLICE\[1\].RAM8.DEC1.AND7/C SLICE\[1\].RAM8.DEC1.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC1.AND7/X
+ sky130_fd_sc_hd__and4_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV SLICE\[0\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_7_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_25_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_25_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_8_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_33_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_27_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[7\].DIODE\[1\] BYTE\[7\].FLOATBUF0\[57\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XBYTE\[1\].FLOATBUF1\[8\] TIE1\[1\]/LO FBUFENBUF1\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.DEC0.AND3 SLICE\[3\].RAM8.DEC0.AND7/C SLICE\[3\].RAM8.DEC0.AND7/B
+ SLICE\[3\].RAM8.DEC0.AND7/A SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WEBUF\[3\] WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WEBUF\[3\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_23_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_11_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_12_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_5_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF SLICE\[1\].RAM8.DEC0.AND3/X VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XFBUFENBUF1\[3\] EN1 VGND VGND VPWR VPWR FBUFENBUF1\[3\]/X sky130_fd_sc_hd__clkbuf_2
Xtap_13_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_8_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_8_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[2\] Do0_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF0\[50\]/Z
+ VGND VGND VPWR VPWR Do0[50] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_33_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.DEC0.ENBUF DEC0.AND2/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.AND7/D
+ sky130_fd_sc_hd__clkbuf_2
Xfill_26_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_19_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.DEC0.ABUF\[1\] A0BUF\[1\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.AND7/B
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_18_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[2\] BYTE\[1\].FLOATBUF1\[10\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_34_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_34_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV SLICE\[2\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_22_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_22_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_5_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_5_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_10_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV SLICE\[1\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[5\] BYTE\[3\].FLOATBUF0\[29\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_31_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
Xfill_24_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_17_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.Do_CLKBUF\[4\] Do0_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do0_REG.Do_CLKBUF\[4\]/X
+ sky130_fd_sc_hd__clkbuf_4
Xfill_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_20_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[9\] Di0[9] VGND VGND VPWR VPWR DIBUF\[9\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_29_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[3\] Do1_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF1\[3\]/Z
+ VGND VGND VPWR VPWR Do1[3] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.SEL1BUF SLICE\[3\].RAM8.DEC1.AND1/X VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[1\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_17_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_33_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_10_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_5_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[6\] Do0_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF0\[22\]/Z
+ VGND VGND VPWR VPWR Do0[22] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[61\] Di0[61] VGND VGND VPWR VPWR DIBUF\[61\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_15_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_22_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfill_15_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_31_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WEBUF\[0\] WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WEBUF\[0\]/X
+ sky130_fd_sc_hd__clkbuf_2
Xtap_31_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_2_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XTIE1\[5\] VGND VGND VPWR VPWR TIE1\[5\]/HI TIE1\[5\]/LO sky130_fd_sc_hd__conb_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_21_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[2\].FLOATBUF0\[22\] TIE0\[2\]/LO FBUFENBUF0\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV SLICE\[1\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_6_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[6\].FLOATBUF0\[53\] TIE0\[6\]/LO FBUFENBUF0\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_26_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_14_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_14_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_30_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_16_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XDo1_REG.OUTREG_BYTE\[6\].DIODE\[2\] BYTE\[6\].FLOATBUF1\[50\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_4_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[24\] Di0[24] VGND VGND VPWR VPWR DIBUF\[24\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_14_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_7_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF SLICE\[1\].RAM8.DEC0.AND2/X VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_25_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XA0BUF\[4\] A0[4] VGND VGND VPWR VPWR DEC0.AND3/A sky130_fd_sc_hd__clkbuf_2
Xtap_8_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_33_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_27_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.DEC0.AND4 SLICE\[3\].RAM8.DEC0.AND7/A SLICE\[3\].RAM8.DEC0.AND7/B
+ SLICE\[3\].RAM8.DEC0.AND7/C SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.AND4/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[5\].Do_FF\[3\] Do1_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF1\[43\]/Z
+ VGND VGND VPWR VPWR Do1[43] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_23_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV SLICE\[2\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_11_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_12_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_5_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV SLICE\[1\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[2\] BYTE\[0\].FLOATBUF0\[2\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_13_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[6\] Do0_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF0\[62\]/Z
+ VGND VGND VPWR VPWR Do0[62] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[0\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[4\].FLOATBUF0\[34\] TIE0\[4\]/LO FBUFENBUF0\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_26_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_19_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[6\] BYTE\[2\].FLOATBUF1\[22\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.SEL1BUF SLICE\[3\].RAM8.DEC1.AND0/Y VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[0\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_18_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_0_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_22_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_22_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_5_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_5_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_5_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_3_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_31_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_24_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[7\] Do1_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF1\[15\]/Z
+ VGND VGND VPWR VPWR Do1[15] sky130_fd_sc_hd__dfxtp_1
Xfill_17_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_0_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_0_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[10\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.DEC0.ABUF\[2\] A0BUF\[2\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.AND7/C
+ sky130_fd_sc_hd__clkbuf_2
Xtap_29_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_17_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_17_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_10_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_19_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV SLICE\[2\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XDIBUF\[54\] Di0[54] VGND VGND VPWR VPWR DIBUF\[54\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_22_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_15_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xtap_31_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_2_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_28_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.Do_CLKBUF\[0\] Do1_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do1_REG.Do_CLKBUF\[0\]/X
+ sky130_fd_sc_hd__clkbuf_4
Xtap_21_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XTIE0\[0\] VGND VGND VPWR VPWR TIE0\[0\]/HI TIE0\[0\]/LO sky130_fd_sc_hd__conb_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_26_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF SLICE\[1\].RAM8.DEC0.AND1/X VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_14_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[5\].DIODE\[2\] BYTE\[5\].FLOATBUF0\[42\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfill_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_30_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_30_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[55\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_32_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[7\].DIODE\[6\] BYTE\[7\].FLOATBUF1\[62\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[0\] Do1_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF1\[16\]/Z
+ VGND VGND VPWR VPWR Do1[16] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV SLICE\[2\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XDIBUF\[17\] Di0[17] VGND VGND VPWR VPWR DIBUF\[17\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_7_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[3\] Do0_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF0\[35\]/Z
+ VGND VGND VPWR VPWR Do0[35] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_25_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_25_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV SLICE\[1\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_8_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_33_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_26_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_19_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[6\].Do_FF\[7\] Do1_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF1\[55\]/Z
+ VGND VGND VPWR VPWR Do1[55] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.DEC0.AND5 SLICE\[3\].RAM8.DEC0.AND7/B SLICE\[3\].RAM8.DEC0.AND7/A
+ SLICE\[3\].RAM8.DEC0.AND7/C SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.AND5/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_2_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[6\] BYTE\[1\].FLOATBUF0\[14\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_12_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_5_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_13_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_8_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_26_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_19_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[7\] Do0_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF0\[7\]/Z
+ VGND VGND VPWR VPWR Do0[7] sky130_fd_sc_hd__dfxtp_1
Xfill_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_22_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_5_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV SLICE\[3\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_3_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_24_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV SLICE\[2\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.SEL1BUF SLICE\[2\].RAM8.DEC1.AND7/X VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[7\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_31_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_17_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_0_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_29_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_17_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XDIODE_A0\[4\] A0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XDo1_REG.OUTREG_BYTE\[7\].Do_FF\[0\] Do1_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF1\[56\]/Z
+ VGND VGND VPWR VPWR Do1[56] sky130_fd_sc_hd__dfxtp_1
Xtap_19_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_1_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF SLICE\[1\].RAM8.DEC0.AND0/Y VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XWEBUF\[4\] WE0[4] VGND VGND VPWR VPWR WEBUF\[4\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[47\] Di0[47] VGND VGND VPWR VPWR DIBUF\[47\]/X sky130_fd_sc_hd__clkbuf_16
XBYTE\[2\].FLOATBUF1\[20\] TIE1\[2\]/LO FBUFENBUF1\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_15_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[6\].FLOATBUF1\[51\] TIE1\[6\]/LO FBUFENBUF1\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_2_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_28_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[4\].DIODE\[3\] BYTE\[4\].FLOATBUF1\[35\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV SLICE\[2\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[6\].DIODE\[6\] BYTE\[6\].FLOATBUF0\[54\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WEBUF\[4\] WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[4\]/X
+ sky130_fd_sc_hd__clkbuf_2
Xfill_6_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[0\] Do0_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF0\[8\]/Z
+ VGND VGND VPWR VPWR Do0[8] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_20_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_30_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_28_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[4\] Do1_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF1\[28\]/Z
+ VGND VGND VPWR VPWR Do1[28] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_32_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_4_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[7\] Do0_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF0\[47\]/Z
+ VGND VGND VPWR VPWR Do0[47] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_25_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_25_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_8_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[7\] BYTE\[0\].FLOATBUF1\[7\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_33_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_26_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[0\].FLOATBUF0\[4\] TIE0\[0\]/LO FBUFENBUF0\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_27_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_19_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_27_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.DEC0.AND6 SLICE\[3\].RAM8.DEC0.AND7/A SLICE\[3\].RAM8.DEC0.AND7/B
+ SLICE\[3\].RAM8.DEC0.AND7/C SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.AND6/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_3_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_3_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_2_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[4\].FLOATBUF1\[32\] TIE1\[4\]/LO FBUFENBUF1\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV SLICE\[3\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XBYTE\[5\].FLOATBUF1\[47\] TIE1\[5\]/LO FBUFENBUF1\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_12_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_5_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV SLICE\[2\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_31_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.SEL1BUF SLICE\[2\].RAM8.DEC1.AND6/X VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[6\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_19_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WEBUF\[1\] WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WEBUF\[1\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_5_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_5_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_3_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XFBUFENBUF1\[1\] EN1 VGND VGND VPWR VPWR FBUFENBUF1\[1\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_12_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[0\] Do0_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF0\[48\]/Z
+ VGND VGND VPWR VPWR Do0[48] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_31_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_17_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_9_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[0\] BYTE\[1\].FLOATBUF1\[8\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfill_17_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_10_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_10_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_10_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_19_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_19_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_1_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[3\] BYTE\[3\].FLOATBUF0\[27\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV SLICE\[3\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_22_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_15_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.Do_CLKBUF\[2\] Do0_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do0_REG.Do_CLKBUF\[2\]/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[3\].FLOATBUF1\[28\] TIE1\[3\]/LO FBUFENBUF1\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[7\] Di0[7] VGND VGND VPWR VPWR DIBUF\[7\]/X sky130_fd_sc_hd__clkbuf_16
XDo1_REG.OUTREG_BYTE\[5\].DIODE\[7\] BYTE\[5\].FLOATBUF1\[47\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_2_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[1\] Do1_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF1\[1\]/Z
+ VGND VGND VPWR VPWR Do1[1] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_28_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XBYTE\[7\].FLOATBUF1\[59\] TIE1\[7\]/LO FBUFENBUF1\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[36\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF SLICE\[0\].RAM8.DEC0.AND7/X VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[4\] Do0_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF0\[20\]/Z
+ VGND VGND VPWR VPWR Do0[20] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_6_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_6_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_20_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfill_13_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_28_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_16_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTIE1\[3\] VGND VGND VPWR VPWR TIE1\[3\]/HI TIE1\[3\]/LO sky130_fd_sc_hd__conb_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_32_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_20_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[2\].FLOATBUF0\[20\] TIE0\[2\]/LO FBUFENBUF0\[2\]/X VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_4_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[6\].FLOATBUF0\[51\] TIE0\[6\]/LO FBUFENBUF0\[6\]/X VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV SLICE\[3\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_25_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_8_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_8_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV SLICE\[2\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.SEL1BUF SLICE\[2\].RAM8.DEC1.AND5/X VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[5\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_33_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_26_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_27_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.DEC0.AND7 SLICE\[3\].RAM8.DEC0.AND7/A SLICE\[3\].RAM8.DEC0.AND7/B
+ SLICE\[3\].RAM8.DEC0.AND7/C SLICE\[3\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.AND7/X
+ sky130_fd_sc_hd__and4_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.DEC0.AND0 SLICE\[1\].RAM8.DEC0.AND7/A SLICE\[1\].RAM8.DEC0.AND7/B
+ SLICE\[1\].RAM8.DEC0.AND7/C SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.AND0/Y
+ sky130_fd_sc_hd__nor4b_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_3_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_3_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDo1_REG.OUTREG_BYTE\[6\].DIODE\[0\] BYTE\[6\].FLOATBUF1\[48\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[22\] Di0[22] VGND VGND VPWR VPWR DIBUF\[22\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_12_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_5_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XA0BUF\[2\] A0[2] VGND VGND VPWR VPWR A0BUF\[2\]/X sky130_fd_sc_hd__clkbuf_2
Xtap_13_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_31_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[5\].Do_FF\[1\] Do1_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF1\[41\]/Z
+ VGND VGND VPWR VPWR Do1[41] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_5_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_5_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_10_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_24_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[0\] BYTE\[0\].FLOATBUF0\[0\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[4\] Do0_REG.Do_CLKBUF\[7\]/X BYTE\[7\].FLOATBUF0\[60\]/Z
+ VGND VGND VPWR VPWR Do0[60] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_12_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_12_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV SLICE\[3\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_31_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBYTE\[4\].FLOATBUF0\[32\] TIE0\[4\]/LO FBUFENBUF0\[4\]/X VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_24_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBYTE\[5\].FLOATBUF0\[47\] TIE0\[5\]/LO FBUFENBUF0\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[4\] BYTE\[2\].FLOATBUF1\[20\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_9_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_33_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
Xtap_10_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF SLICE\[0\].RAM8.DEC0.AND6/X VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[4\].DIODE\[7\] BYTE\[4\].FLOATBUF0\[39\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_1_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[32\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_23_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_22_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[5\] Do1_REG.Do_CLKBUF\[1\]/X BYTE\[1\].FLOATBUF1\[13\]/Z
+ VGND VGND VPWR VPWR Do1[13] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_15_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.DEC0.ABUF\[0\] A0BUF\[0\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.AND7/A
+ sky130_fd_sc_hd__clkbuf_2
Xtap_2_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_2_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_28_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_21_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_21_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[21\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_18_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV SLICE\[3\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_6_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_6_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[52\] Di0[52] VGND VGND VPWR VPWR DIBUF\[52\]/X sky130_fd_sc_hd__clkbuf_16
Xfill_20_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_13_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WEBUF\[6\] WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WEBUF\[6\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.SEL1BUF SLICE\[2\].RAM8.DEC1.AND4/X VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[4\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_28_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_20_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_20_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[3\].FLOATBUF0\[28\] TIE0\[3\]/LO FBUFENBUF0\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XFBUFENBUF0\[7\] EN0 VGND VGND VPWR VPWR FBUFENBUF0\[7\]/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XBYTE\[7\].FLOATBUF0\[59\] TIE0\[7\]/LO FBUFENBUF0\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_9_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_8_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_8_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[5\].DIODE\[0\] BYTE\[5\].FLOATBUF0\[40\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_8_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_33_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_27_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_27_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_27_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_15_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_15_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XDo1_REG.OUTREG_BYTE\[7\].DIODE\[4\] BYTE\[7\].FLOATBUF1\[60\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfill_31_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.DEC0.AND1 SLICE\[1\].RAM8.DEC0.AND7/C SLICE\[1\].RAM8.DEC0.AND7/B
+ SLICE\[1\].RAM8.DEC0.AND7/A SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.AND1/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_3_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[15\] Di0[15] VGND VGND VPWR VPWR DIBUF\[15\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[0\].FLOATBUF1\[7\] TIE1\[0\]/LO FBUFENBUF1\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_5_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[1\] Do0_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF0\[33\]/Z
+ VGND VGND VPWR VPWR Do0[33] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_13_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_31_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV SLICE\[3\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[6\].Do_FF\[5\] Do1_REG.Do_CLKBUF\[6\]/X BYTE\[6\].FLOATBUF1\[53\]/Z
+ VGND VGND VPWR VPWR Do1[53] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_0_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_5_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[4\] BYTE\[1\].FLOATBUF0\[12\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF SLICE\[0\].RAM8.DEC0.AND5/X VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
Xtap_10_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
Xtap_3_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.DEC1.ABUF\[1\] A1BUF\[1\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC1.AND7/B
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_12_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_12_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_17_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_0_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_9_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_9_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[5\] Do0_REG.Do_CLKBUF\[0\]/X BYTE\[0\].FLOATBUF0\[5\]/Z
+ VGND VGND VPWR VPWR Do0[5] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_10_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_19_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_19_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_1_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[17\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_23_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_23_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[7\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_22_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV SLICE\[0\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[1\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_15_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.SEL1BUF SLICE\[2\].RAM8.DEC1.AND3/X VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[3\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_2_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIODE_A0\[2\] A0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_21_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[6\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_18_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_6_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XWEBUF\[2\] WE0[2] VGND VGND VPWR VPWR WEBUF\[2\]/X sky130_fd_sc_hd__clkbuf_2
Xfill_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDIBUF\[45\] Di0[45] VGND VGND VPWR VPWR DIBUF\[45\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_13_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_28_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_16_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_16_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[4\].DIODE\[1\] BYTE\[4\].FLOATBUF1\[33\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xtap_32_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_20_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_20_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_3_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[6\].DIODE\[4\] BYTE\[6\].FLOATBUF0\[52\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WEBUF\[2\] WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[2\]/X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\]/X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[62\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_9_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xtap_8_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_33_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV SLICE\[3\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xtap_26_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[6\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_27_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_27_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[2\] Do1_REG.Do_CLKBUF\[3\]/X BYTE\[3\].FLOATBUF1\[26\]/Z
+ VGND VGND VPWR VPWR Do1[26] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_15_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_31_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_31_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.DEC0.AND2 SLICE\[1\].RAM8.DEC0.AND7/C SLICE\[1\].RAM8.DEC0.AND7/A
+ SLICE\[1\].RAM8.DEC0.AND7/B SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.AND2/X
+ sky130_fd_sc_hd__and4bb_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_3_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_3_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_2_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[5\] Do0_REG.Do_CLKBUF\[5\]/X BYTE\[5\].FLOATBUF0\[45\]/Z
+ VGND VGND VPWR VPWR Do0[45] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF SLICE\[0\].RAM8.DEC0.AND4/X VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.CLKBUF/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_13_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[5\] BYTE\[0\].FLOATBUF1\[5\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_31_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[0\].FLOATBUF0\[2\] TIE0\[0\]/LO FBUFENBUF0\[0\]/X VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_17_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_0_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[5\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_26_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[1\].FLOATBUF1\[14\] TIE1\[1\]/LO FBUFENBUF1\[1\]/X VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_0_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[4\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_5_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_5_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XBYTE\[5\].FLOATBUF1\[45\] TIE1\[5\]/LO FBUFENBUF1\[5\]/X VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xtap_3_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_24_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_24_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xfill_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_12_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV SLICE\[0\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[2\].RAM8.WEBUF\[4\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_17_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\]/X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.SEL1BUF SLICE\[2\].RAM8.DEC1.AND2/X VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[2\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
Xfill_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_9_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_34_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_29_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_10_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_10_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[7\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_19_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_19_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_1_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[2\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_23_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_23_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_23_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_6_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_15_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[3\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_2_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\]/X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_21_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_21_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_21_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[5\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[50\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[29\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_18_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_18_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[1\] BYTE\[3\].FLOATBUF0\[25\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\]/X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_6_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_6_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
Xfill_20_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[38\] Di0[38] VGND VGND VPWR VPWR DIBUF\[38\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0_REG.Do_CLKBUF\[0\] Do0_REG.Root_CLKBUF/X VGND VGND VPWR VPWR Do0_REG.Do_CLKBUF\[0\]/X
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XBYTE\[3\].FLOATBUF1\[26\] TIE1\[3\]/LO FBUFENBUF1\[3\]/X VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[58\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDIBUF\[5\] Di0[5] VGND VGND VPWR VPWR DIBUF\[5\]/X sky130_fd_sc_hd__clkbuf_16
XDo1_REG.OUTREG_BYTE\[5\].DIODE\[5\] BYTE\[5\].FLOATBUF1\[45\]/Z VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_28_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF/X
+ SLICE\[0\].RAM8.WEBUF\[1\]/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtap_16_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XBYTE\[7\].FLOATBUF1\[57\] TIE1\[7\]/LO FBUFENBUF1\[7\]/X VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[39\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_32_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV SLICE\[0\].RAM8.WORD\[2\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/CLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\]/X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_20_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_20_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_3_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_29_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\]/X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\]/X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[2\] Do0_REG.Do_CLKBUF\[2\]/X BYTE\[2\].FLOATBUF0\[18\]/Z
+ VGND VGND VPWR VPWR Do0[18] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[18\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF SLICE\[0\].RAM8.DEC0.AND3/X VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[20\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[47\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_9_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDo1_REG.OUTREG_BYTE\[4\].Do_FF\[6\] Do1_REG.Do_CLKBUF\[4\]/X BYTE\[4\].FLOATBUF1\[38\]/Z
+ VGND VGND VPWR VPWR Do1[38] sky130_fd_sc_hd__dfxtp_1
Xtap_33_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[38\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF1\[48\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_26_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_27_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF/X
+ SLICE\[1\].RAM8.WEBUF\[0\]/X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\]/X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\]/Z
+ sky130_fd_sc_hd__ebufn_2
XTIE1\[1\] VGND VGND VPWR VPWR TIE1\[1\]/HI TIE1\[1\]/LO sky130_fd_sc_hd__conb_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\]/X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_15_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[26\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[1\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_31_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfill_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_31_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[0\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[28\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.DEC0.AND3 SLICE\[1\].RAM8.DEC0.AND7/C SLICE\[1\].RAM8.DEC0.AND7/B
+ SLICE\[1\].RAM8.DEC0.AND7/A SLICE\[1\].RAM8.DEC0.AND7/D VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.AND3/X
+ sky130_fd_sc_hd__and4b_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF/X
+ SLICE\[3\].RAM8.WEBUF\[2\]/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND/X
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[7\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xfill_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_3_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_3_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\]/X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_2_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF1\[19\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\]/X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\]/X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\]/X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[46\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\]/X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[56\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[2\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\]/X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_13_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[7\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[9\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF1\[37\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_13_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.DEC0.ABUF\[1\] A0BUF\[1\]/X VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.AND7/B
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[3\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_31_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[15\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_17_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\]/X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF1\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\]/X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xtap_0_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV SLICE\[0\].RAM8.WORD\[6\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
Xfill_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_26_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF1\[27\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[3\].W.SEL1BUF/X
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV/Y sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_9_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.SEL1BUF SLICE\[2\].RAM8.DEC1.AND1/X VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[1\].W.SEL1BUF/X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\]/X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\]/X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\]/X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\]/X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
Xfill_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF1/A
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF1\[45\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF1/A
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\]/Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[20\] Di0[20] VGND VGND VPWR VPWR DIBUF\[20\]/X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[6\].W.CLKBUF/X
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG/CLK sky130_fd_sc_hd__inv_1
Xtap_5_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/CLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND/X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF1\[57\]/Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF1/A
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV/Y VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_5_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1/A
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV/Y VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF1\[8\]/Z
+ sky130_fd_sc_hd__ebufn_2
Xtap_10_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\]/X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG/GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF1/A sky130_fd_sc_hd__dlxtp_1
.ends

