magic
tech sky130B
magscale 1 2
timestamp 1662419308
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 290 1708 99990 98524
<< metal2 >>
rect 2502 99200 2558 100000
rect 3238 99200 3294 100000
rect 3974 99200 4030 100000
rect 4710 99200 4766 100000
rect 5446 99200 5502 100000
rect 6182 99200 6238 100000
rect 6918 99200 6974 100000
rect 7654 99200 7710 100000
rect 8390 99200 8446 100000
rect 9126 99200 9182 100000
rect 9862 99200 9918 100000
rect 10598 99200 10654 100000
rect 11334 99200 11390 100000
rect 12070 99200 12126 100000
rect 12806 99200 12862 100000
rect 13542 99200 13598 100000
rect 14278 99200 14334 100000
rect 15014 99200 15070 100000
rect 15750 99200 15806 100000
rect 16486 99200 16542 100000
rect 17222 99200 17278 100000
rect 17958 99200 18014 100000
rect 18694 99200 18750 100000
rect 19430 99200 19486 100000
rect 20166 99200 20222 100000
rect 20902 99200 20958 100000
rect 21638 99200 21694 100000
rect 22374 99200 22430 100000
rect 23110 99200 23166 100000
rect 23846 99200 23902 100000
rect 24582 99200 24638 100000
rect 25318 99200 25374 100000
rect 26054 99200 26110 100000
rect 26790 99200 26846 100000
rect 27526 99200 27582 100000
rect 28262 99200 28318 100000
rect 28998 99200 29054 100000
rect 29734 99200 29790 100000
rect 30470 99200 30526 100000
rect 31206 99200 31262 100000
rect 31942 99200 31998 100000
rect 32678 99200 32734 100000
rect 33414 99200 33470 100000
rect 34150 99200 34206 100000
rect 34886 99200 34942 100000
rect 35622 99200 35678 100000
rect 36358 99200 36414 100000
rect 37094 99200 37150 100000
rect 37830 99200 37886 100000
rect 38566 99200 38622 100000
rect 39302 99200 39358 100000
rect 40038 99200 40094 100000
rect 40774 99200 40830 100000
rect 41510 99200 41566 100000
rect 42246 99200 42302 100000
rect 42982 99200 43038 100000
rect 43718 99200 43774 100000
rect 44454 99200 44510 100000
rect 45190 99200 45246 100000
rect 45926 99200 45982 100000
rect 46662 99200 46718 100000
rect 47398 99200 47454 100000
rect 48134 99200 48190 100000
rect 48870 99200 48926 100000
rect 49606 99200 49662 100000
rect 50342 99200 50398 100000
rect 51078 99200 51134 100000
rect 51814 99200 51870 100000
rect 52550 99200 52606 100000
rect 53286 99200 53342 100000
rect 54022 99200 54078 100000
rect 54758 99200 54814 100000
rect 55494 99200 55550 100000
rect 56230 99200 56286 100000
rect 56966 99200 57022 100000
rect 57702 99200 57758 100000
rect 58438 99200 58494 100000
rect 59174 99200 59230 100000
rect 59910 99200 59966 100000
rect 60646 99200 60702 100000
rect 61382 99200 61438 100000
rect 62118 99200 62174 100000
rect 62854 99200 62910 100000
rect 63590 99200 63646 100000
rect 64326 99200 64382 100000
rect 65062 99200 65118 100000
rect 65798 99200 65854 100000
rect 66534 99200 66590 100000
rect 67270 99200 67326 100000
rect 68006 99200 68062 100000
rect 68742 99200 68798 100000
rect 69478 99200 69534 100000
rect 70214 99200 70270 100000
rect 70950 99200 71006 100000
rect 71686 99200 71742 100000
rect 72422 99200 72478 100000
rect 73158 99200 73214 100000
rect 73894 99200 73950 100000
rect 74630 99200 74686 100000
rect 75366 99200 75422 100000
rect 76102 99200 76158 100000
rect 76838 99200 76894 100000
rect 77574 99200 77630 100000
rect 78310 99200 78366 100000
rect 79046 99200 79102 100000
rect 79782 99200 79838 100000
rect 80518 99200 80574 100000
rect 81254 99200 81310 100000
rect 81990 99200 82046 100000
rect 82726 99200 82782 100000
rect 83462 99200 83518 100000
rect 84198 99200 84254 100000
rect 84934 99200 84990 100000
rect 85670 99200 85726 100000
rect 86406 99200 86462 100000
rect 87142 99200 87198 100000
rect 87878 99200 87934 100000
rect 88614 99200 88670 100000
rect 89350 99200 89406 100000
rect 90086 99200 90142 100000
rect 90822 99200 90878 100000
rect 91558 99200 91614 100000
rect 92294 99200 92350 100000
rect 93030 99200 93086 100000
rect 93766 99200 93822 100000
rect 94502 99200 94558 100000
rect 95238 99200 95294 100000
rect 95974 99200 96030 100000
rect 96710 99200 96766 100000
rect 97446 99200 97502 100000
rect 3238 0 3294 800
rect 3974 0 4030 800
rect 4710 0 4766 800
rect 5446 0 5502 800
rect 6182 0 6238 800
rect 6918 0 6974 800
rect 7654 0 7710 800
rect 8390 0 8446 800
rect 9126 0 9182 800
rect 9862 0 9918 800
rect 10598 0 10654 800
rect 11334 0 11390 800
rect 12070 0 12126 800
rect 12806 0 12862 800
rect 13542 0 13598 800
rect 14278 0 14334 800
rect 15014 0 15070 800
rect 15750 0 15806 800
rect 16486 0 16542 800
rect 17222 0 17278 800
rect 17958 0 18014 800
rect 18694 0 18750 800
rect 19430 0 19486 800
rect 20166 0 20222 800
rect 20902 0 20958 800
rect 21638 0 21694 800
rect 22374 0 22430 800
rect 23110 0 23166 800
rect 23846 0 23902 800
rect 24582 0 24638 800
rect 25318 0 25374 800
rect 26054 0 26110 800
rect 26790 0 26846 800
rect 27526 0 27582 800
rect 28262 0 28318 800
rect 28998 0 29054 800
rect 29734 0 29790 800
rect 30470 0 30526 800
rect 31206 0 31262 800
rect 31942 0 31998 800
rect 32678 0 32734 800
rect 33414 0 33470 800
rect 34150 0 34206 800
rect 34886 0 34942 800
rect 35622 0 35678 800
rect 36358 0 36414 800
rect 37094 0 37150 800
rect 37830 0 37886 800
rect 38566 0 38622 800
rect 39302 0 39358 800
rect 40038 0 40094 800
rect 40774 0 40830 800
rect 41510 0 41566 800
rect 42246 0 42302 800
rect 42982 0 43038 800
rect 43718 0 43774 800
rect 44454 0 44510 800
rect 45190 0 45246 800
rect 45926 0 45982 800
rect 46662 0 46718 800
rect 47398 0 47454 800
rect 48134 0 48190 800
rect 48870 0 48926 800
rect 49606 0 49662 800
rect 50342 0 50398 800
rect 51078 0 51134 800
rect 51814 0 51870 800
rect 52550 0 52606 800
rect 53286 0 53342 800
rect 54022 0 54078 800
rect 54758 0 54814 800
rect 55494 0 55550 800
rect 56230 0 56286 800
rect 56966 0 57022 800
rect 57702 0 57758 800
rect 58438 0 58494 800
rect 59174 0 59230 800
rect 59910 0 59966 800
rect 60646 0 60702 800
rect 61382 0 61438 800
rect 62118 0 62174 800
rect 62854 0 62910 800
rect 63590 0 63646 800
rect 64326 0 64382 800
rect 65062 0 65118 800
rect 65798 0 65854 800
rect 66534 0 66590 800
rect 67270 0 67326 800
rect 68006 0 68062 800
rect 68742 0 68798 800
rect 69478 0 69534 800
rect 70214 0 70270 800
rect 70950 0 71006 800
rect 71686 0 71742 800
rect 72422 0 72478 800
rect 73158 0 73214 800
rect 73894 0 73950 800
rect 74630 0 74686 800
rect 75366 0 75422 800
rect 76102 0 76158 800
rect 76838 0 76894 800
rect 77574 0 77630 800
rect 78310 0 78366 800
rect 79046 0 79102 800
rect 79782 0 79838 800
rect 80518 0 80574 800
rect 81254 0 81310 800
rect 81990 0 82046 800
rect 82726 0 82782 800
rect 83462 0 83518 800
rect 84198 0 84254 800
rect 84934 0 84990 800
rect 85670 0 85726 800
rect 86406 0 86462 800
rect 87142 0 87198 800
rect 87878 0 87934 800
rect 88614 0 88670 800
rect 89350 0 89406 800
rect 90086 0 90142 800
rect 90822 0 90878 800
rect 91558 0 91614 800
rect 92294 0 92350 800
rect 93030 0 93086 800
rect 93766 0 93822 800
rect 94502 0 94558 800
rect 95238 0 95294 800
rect 95974 0 96030 800
rect 96710 0 96766 800
<< obsm2 >>
rect 202 99144 2446 99362
rect 2614 99144 3182 99362
rect 3350 99144 3918 99362
rect 4086 99144 4654 99362
rect 4822 99144 5390 99362
rect 5558 99144 6126 99362
rect 6294 99144 6862 99362
rect 7030 99144 7598 99362
rect 7766 99144 8334 99362
rect 8502 99144 9070 99362
rect 9238 99144 9806 99362
rect 9974 99144 10542 99362
rect 10710 99144 11278 99362
rect 11446 99144 12014 99362
rect 12182 99144 12750 99362
rect 12918 99144 13486 99362
rect 13654 99144 14222 99362
rect 14390 99144 14958 99362
rect 15126 99144 15694 99362
rect 15862 99144 16430 99362
rect 16598 99144 17166 99362
rect 17334 99144 17902 99362
rect 18070 99144 18638 99362
rect 18806 99144 19374 99362
rect 19542 99144 20110 99362
rect 20278 99144 20846 99362
rect 21014 99144 21582 99362
rect 21750 99144 22318 99362
rect 22486 99144 23054 99362
rect 23222 99144 23790 99362
rect 23958 99144 24526 99362
rect 24694 99144 25262 99362
rect 25430 99144 25998 99362
rect 26166 99144 26734 99362
rect 26902 99144 27470 99362
rect 27638 99144 28206 99362
rect 28374 99144 28942 99362
rect 29110 99144 29678 99362
rect 29846 99144 30414 99362
rect 30582 99144 31150 99362
rect 31318 99144 31886 99362
rect 32054 99144 32622 99362
rect 32790 99144 33358 99362
rect 33526 99144 34094 99362
rect 34262 99144 34830 99362
rect 34998 99144 35566 99362
rect 35734 99144 36302 99362
rect 36470 99144 37038 99362
rect 37206 99144 37774 99362
rect 37942 99144 38510 99362
rect 38678 99144 39246 99362
rect 39414 99144 39982 99362
rect 40150 99144 40718 99362
rect 40886 99144 41454 99362
rect 41622 99144 42190 99362
rect 42358 99144 42926 99362
rect 43094 99144 43662 99362
rect 43830 99144 44398 99362
rect 44566 99144 45134 99362
rect 45302 99144 45870 99362
rect 46038 99144 46606 99362
rect 46774 99144 47342 99362
rect 47510 99144 48078 99362
rect 48246 99144 48814 99362
rect 48982 99144 49550 99362
rect 49718 99144 50286 99362
rect 50454 99144 51022 99362
rect 51190 99144 51758 99362
rect 51926 99144 52494 99362
rect 52662 99144 53230 99362
rect 53398 99144 53966 99362
rect 54134 99144 54702 99362
rect 54870 99144 55438 99362
rect 55606 99144 56174 99362
rect 56342 99144 56910 99362
rect 57078 99144 57646 99362
rect 57814 99144 58382 99362
rect 58550 99144 59118 99362
rect 59286 99144 59854 99362
rect 60022 99144 60590 99362
rect 60758 99144 61326 99362
rect 61494 99144 62062 99362
rect 62230 99144 62798 99362
rect 62966 99144 63534 99362
rect 63702 99144 64270 99362
rect 64438 99144 65006 99362
rect 65174 99144 65742 99362
rect 65910 99144 66478 99362
rect 66646 99144 67214 99362
rect 67382 99144 67950 99362
rect 68118 99144 68686 99362
rect 68854 99144 69422 99362
rect 69590 99144 70158 99362
rect 70326 99144 70894 99362
rect 71062 99144 71630 99362
rect 71798 99144 72366 99362
rect 72534 99144 73102 99362
rect 73270 99144 73838 99362
rect 74006 99144 74574 99362
rect 74742 99144 75310 99362
rect 75478 99144 76046 99362
rect 76214 99144 76782 99362
rect 76950 99144 77518 99362
rect 77686 99144 78254 99362
rect 78422 99144 78990 99362
rect 79158 99144 79726 99362
rect 79894 99144 80462 99362
rect 80630 99144 81198 99362
rect 81366 99144 81934 99362
rect 82102 99144 82670 99362
rect 82838 99144 83406 99362
rect 83574 99144 84142 99362
rect 84310 99144 84878 99362
rect 85046 99144 85614 99362
rect 85782 99144 86350 99362
rect 86518 99144 87086 99362
rect 87254 99144 87822 99362
rect 87990 99144 88558 99362
rect 88726 99144 89294 99362
rect 89462 99144 90030 99362
rect 90198 99144 90766 99362
rect 90934 99144 91502 99362
rect 91670 99144 92238 99362
rect 92406 99144 92974 99362
rect 93142 99144 93710 99362
rect 93878 99144 94446 99362
rect 94614 99144 95182 99362
rect 95350 99144 95918 99362
rect 96086 99144 96654 99362
rect 96822 99144 97390 99362
rect 97558 99144 99986 99362
rect 202 856 99986 99144
rect 202 734 3182 856
rect 3350 734 3918 856
rect 4086 734 4654 856
rect 4822 734 5390 856
rect 5558 734 6126 856
rect 6294 734 6862 856
rect 7030 734 7598 856
rect 7766 734 8334 856
rect 8502 734 9070 856
rect 9238 734 9806 856
rect 9974 734 10542 856
rect 10710 734 11278 856
rect 11446 734 12014 856
rect 12182 734 12750 856
rect 12918 734 13486 856
rect 13654 734 14222 856
rect 14390 734 14958 856
rect 15126 734 15694 856
rect 15862 734 16430 856
rect 16598 734 17166 856
rect 17334 734 17902 856
rect 18070 734 18638 856
rect 18806 734 19374 856
rect 19542 734 20110 856
rect 20278 734 20846 856
rect 21014 734 21582 856
rect 21750 734 22318 856
rect 22486 734 23054 856
rect 23222 734 23790 856
rect 23958 734 24526 856
rect 24694 734 25262 856
rect 25430 734 25998 856
rect 26166 734 26734 856
rect 26902 734 27470 856
rect 27638 734 28206 856
rect 28374 734 28942 856
rect 29110 734 29678 856
rect 29846 734 30414 856
rect 30582 734 31150 856
rect 31318 734 31886 856
rect 32054 734 32622 856
rect 32790 734 33358 856
rect 33526 734 34094 856
rect 34262 734 34830 856
rect 34998 734 35566 856
rect 35734 734 36302 856
rect 36470 734 37038 856
rect 37206 734 37774 856
rect 37942 734 38510 856
rect 38678 734 39246 856
rect 39414 734 39982 856
rect 40150 734 40718 856
rect 40886 734 41454 856
rect 41622 734 42190 856
rect 42358 734 42926 856
rect 43094 734 43662 856
rect 43830 734 44398 856
rect 44566 734 45134 856
rect 45302 734 45870 856
rect 46038 734 46606 856
rect 46774 734 47342 856
rect 47510 734 48078 856
rect 48246 734 48814 856
rect 48982 734 49550 856
rect 49718 734 50286 856
rect 50454 734 51022 856
rect 51190 734 51758 856
rect 51926 734 52494 856
rect 52662 734 53230 856
rect 53398 734 53966 856
rect 54134 734 54702 856
rect 54870 734 55438 856
rect 55606 734 56174 856
rect 56342 734 56910 856
rect 57078 734 57646 856
rect 57814 734 58382 856
rect 58550 734 59118 856
rect 59286 734 59854 856
rect 60022 734 60590 856
rect 60758 734 61326 856
rect 61494 734 62062 856
rect 62230 734 62798 856
rect 62966 734 63534 856
rect 63702 734 64270 856
rect 64438 734 65006 856
rect 65174 734 65742 856
rect 65910 734 66478 856
rect 66646 734 67214 856
rect 67382 734 67950 856
rect 68118 734 68686 856
rect 68854 734 69422 856
rect 69590 734 70158 856
rect 70326 734 70894 856
rect 71062 734 71630 856
rect 71798 734 72366 856
rect 72534 734 73102 856
rect 73270 734 73838 856
rect 74006 734 74574 856
rect 74742 734 75310 856
rect 75478 734 76046 856
rect 76214 734 76782 856
rect 76950 734 77518 856
rect 77686 734 78254 856
rect 78422 734 78990 856
rect 79158 734 79726 856
rect 79894 734 80462 856
rect 80630 734 81198 856
rect 81366 734 81934 856
rect 82102 734 82670 856
rect 82838 734 83406 856
rect 83574 734 84142 856
rect 84310 734 84878 856
rect 85046 734 85614 856
rect 85782 734 86350 856
rect 86518 734 87086 856
rect 87254 734 87822 856
rect 87990 734 88558 856
rect 88726 734 89294 856
rect 89462 734 90030 856
rect 90198 734 90766 856
rect 90934 734 91502 856
rect 91670 734 92238 856
rect 92406 734 92974 856
rect 93142 734 93710 856
rect 93878 734 94446 856
rect 94614 734 95182 856
rect 95350 734 95918 856
rect 96086 734 96654 856
rect 96822 734 99986 856
<< metal3 >>
rect 99200 93032 100000 93152
rect 99200 92352 100000 92472
rect 99200 91672 100000 91792
rect 99200 90992 100000 91112
rect 99200 90312 100000 90432
rect 99200 89632 100000 89752
rect 99200 88952 100000 89072
rect 99200 88272 100000 88392
rect 99200 87592 100000 87712
rect 99200 86912 100000 87032
rect 99200 86232 100000 86352
rect 99200 85552 100000 85672
rect 99200 84872 100000 84992
rect 99200 84192 100000 84312
rect 99200 83512 100000 83632
rect 99200 82832 100000 82952
rect 99200 82152 100000 82272
rect 99200 81472 100000 81592
rect 99200 80792 100000 80912
rect 99200 80112 100000 80232
rect 99200 79432 100000 79552
rect 99200 78752 100000 78872
rect 99200 78072 100000 78192
rect 99200 77392 100000 77512
rect 99200 76712 100000 76832
rect 99200 76032 100000 76152
rect 99200 75352 100000 75472
rect 99200 74672 100000 74792
rect 99200 73992 100000 74112
rect 99200 73312 100000 73432
rect 99200 72632 100000 72752
rect 99200 71952 100000 72072
rect 99200 71272 100000 71392
rect 99200 70592 100000 70712
rect 99200 69912 100000 70032
rect 99200 69232 100000 69352
rect 99200 68552 100000 68672
rect 99200 67872 100000 67992
rect 99200 67192 100000 67312
rect 99200 66512 100000 66632
rect 99200 65832 100000 65952
rect 99200 65152 100000 65272
rect 99200 64472 100000 64592
rect 99200 63792 100000 63912
rect 99200 63112 100000 63232
rect 99200 62432 100000 62552
rect 99200 61752 100000 61872
rect 99200 61072 100000 61192
rect 99200 60392 100000 60512
rect 99200 59712 100000 59832
rect 99200 59032 100000 59152
rect 99200 58352 100000 58472
rect 99200 57672 100000 57792
rect 99200 56992 100000 57112
rect 99200 56312 100000 56432
rect 99200 55632 100000 55752
rect 99200 54952 100000 55072
rect 99200 54272 100000 54392
rect 99200 53592 100000 53712
rect 99200 52912 100000 53032
rect 99200 52232 100000 52352
rect 99200 51552 100000 51672
rect 99200 50872 100000 50992
rect 99200 50192 100000 50312
rect 99200 49512 100000 49632
rect 99200 48832 100000 48952
rect 99200 48152 100000 48272
rect 99200 47472 100000 47592
rect 99200 46792 100000 46912
rect 99200 46112 100000 46232
rect 99200 45432 100000 45552
rect 99200 44752 100000 44872
rect 99200 44072 100000 44192
rect 99200 43392 100000 43512
rect 99200 42712 100000 42832
rect 99200 42032 100000 42152
rect 99200 41352 100000 41472
rect 99200 40672 100000 40792
rect 99200 39992 100000 40112
rect 99200 39312 100000 39432
rect 99200 38632 100000 38752
rect 99200 37952 100000 38072
rect 99200 37272 100000 37392
rect 99200 36592 100000 36712
rect 99200 35912 100000 36032
rect 99200 35232 100000 35352
rect 99200 34552 100000 34672
rect 99200 33872 100000 33992
rect 99200 33192 100000 33312
rect 99200 32512 100000 32632
rect 99200 31832 100000 31952
rect 99200 31152 100000 31272
rect 99200 30472 100000 30592
rect 99200 29792 100000 29912
rect 99200 29112 100000 29232
rect 99200 28432 100000 28552
rect 99200 27752 100000 27872
rect 99200 27072 100000 27192
rect 99200 26392 100000 26512
rect 99200 25712 100000 25832
rect 99200 25032 100000 25152
rect 99200 24352 100000 24472
rect 99200 23672 100000 23792
rect 99200 22992 100000 23112
rect 99200 22312 100000 22432
rect 99200 21632 100000 21752
rect 99200 20952 100000 21072
rect 99200 20272 100000 20392
rect 99200 19592 100000 19712
rect 99200 18912 100000 19032
rect 99200 18232 100000 18352
rect 99200 17552 100000 17672
rect 99200 16872 100000 16992
rect 99200 16192 100000 16312
rect 99200 15512 100000 15632
rect 99200 14832 100000 14952
rect 99200 14152 100000 14272
rect 99200 13472 100000 13592
rect 99200 12792 100000 12912
rect 99200 12112 100000 12232
rect 99200 11432 100000 11552
rect 99200 10752 100000 10872
rect 99200 10072 100000 10192
rect 99200 9392 100000 9512
rect 99200 8712 100000 8832
rect 99200 8032 100000 8152
rect 99200 7352 100000 7472
rect 99200 6672 100000 6792
<< obsm3 >>
rect 197 93232 99991 98836
rect 197 92952 99120 93232
rect 197 92552 99991 92952
rect 197 92272 99120 92552
rect 197 91872 99991 92272
rect 197 91592 99120 91872
rect 197 91192 99991 91592
rect 197 90912 99120 91192
rect 197 90512 99991 90912
rect 197 90232 99120 90512
rect 197 89832 99991 90232
rect 197 89552 99120 89832
rect 197 89152 99991 89552
rect 197 88872 99120 89152
rect 197 88472 99991 88872
rect 197 88192 99120 88472
rect 197 87792 99991 88192
rect 197 87512 99120 87792
rect 197 87112 99991 87512
rect 197 86832 99120 87112
rect 197 86432 99991 86832
rect 197 86152 99120 86432
rect 197 85752 99991 86152
rect 197 85472 99120 85752
rect 197 85072 99991 85472
rect 197 84792 99120 85072
rect 197 84392 99991 84792
rect 197 84112 99120 84392
rect 197 83712 99991 84112
rect 197 83432 99120 83712
rect 197 83032 99991 83432
rect 197 82752 99120 83032
rect 197 82352 99991 82752
rect 197 82072 99120 82352
rect 197 81672 99991 82072
rect 197 81392 99120 81672
rect 197 80992 99991 81392
rect 197 80712 99120 80992
rect 197 80312 99991 80712
rect 197 80032 99120 80312
rect 197 79632 99991 80032
rect 197 79352 99120 79632
rect 197 78952 99991 79352
rect 197 78672 99120 78952
rect 197 78272 99991 78672
rect 197 77992 99120 78272
rect 197 77592 99991 77992
rect 197 77312 99120 77592
rect 197 76912 99991 77312
rect 197 76632 99120 76912
rect 197 76232 99991 76632
rect 197 75952 99120 76232
rect 197 75552 99991 75952
rect 197 75272 99120 75552
rect 197 74872 99991 75272
rect 197 74592 99120 74872
rect 197 74192 99991 74592
rect 197 73912 99120 74192
rect 197 73512 99991 73912
rect 197 73232 99120 73512
rect 197 72832 99991 73232
rect 197 72552 99120 72832
rect 197 72152 99991 72552
rect 197 71872 99120 72152
rect 197 71472 99991 71872
rect 197 71192 99120 71472
rect 197 70792 99991 71192
rect 197 70512 99120 70792
rect 197 70112 99991 70512
rect 197 69832 99120 70112
rect 197 69432 99991 69832
rect 197 69152 99120 69432
rect 197 68752 99991 69152
rect 197 68472 99120 68752
rect 197 68072 99991 68472
rect 197 67792 99120 68072
rect 197 67392 99991 67792
rect 197 67112 99120 67392
rect 197 66712 99991 67112
rect 197 66432 99120 66712
rect 197 66032 99991 66432
rect 197 65752 99120 66032
rect 197 65352 99991 65752
rect 197 65072 99120 65352
rect 197 64672 99991 65072
rect 197 64392 99120 64672
rect 197 63992 99991 64392
rect 197 63712 99120 63992
rect 197 63312 99991 63712
rect 197 63032 99120 63312
rect 197 62632 99991 63032
rect 197 62352 99120 62632
rect 197 61952 99991 62352
rect 197 61672 99120 61952
rect 197 61272 99991 61672
rect 197 60992 99120 61272
rect 197 60592 99991 60992
rect 197 60312 99120 60592
rect 197 59912 99991 60312
rect 197 59632 99120 59912
rect 197 59232 99991 59632
rect 197 58952 99120 59232
rect 197 58552 99991 58952
rect 197 58272 99120 58552
rect 197 57872 99991 58272
rect 197 57592 99120 57872
rect 197 57192 99991 57592
rect 197 56912 99120 57192
rect 197 56512 99991 56912
rect 197 56232 99120 56512
rect 197 55832 99991 56232
rect 197 55552 99120 55832
rect 197 55152 99991 55552
rect 197 54872 99120 55152
rect 197 54472 99991 54872
rect 197 54192 99120 54472
rect 197 53792 99991 54192
rect 197 53512 99120 53792
rect 197 53112 99991 53512
rect 197 52832 99120 53112
rect 197 52432 99991 52832
rect 197 52152 99120 52432
rect 197 51752 99991 52152
rect 197 51472 99120 51752
rect 197 51072 99991 51472
rect 197 50792 99120 51072
rect 197 50392 99991 50792
rect 197 50112 99120 50392
rect 197 49712 99991 50112
rect 197 49432 99120 49712
rect 197 49032 99991 49432
rect 197 48752 99120 49032
rect 197 48352 99991 48752
rect 197 48072 99120 48352
rect 197 47672 99991 48072
rect 197 47392 99120 47672
rect 197 46992 99991 47392
rect 197 46712 99120 46992
rect 197 46312 99991 46712
rect 197 46032 99120 46312
rect 197 45632 99991 46032
rect 197 45352 99120 45632
rect 197 44952 99991 45352
rect 197 44672 99120 44952
rect 197 44272 99991 44672
rect 197 43992 99120 44272
rect 197 43592 99991 43992
rect 197 43312 99120 43592
rect 197 42912 99991 43312
rect 197 42632 99120 42912
rect 197 42232 99991 42632
rect 197 41952 99120 42232
rect 197 41552 99991 41952
rect 197 41272 99120 41552
rect 197 40872 99991 41272
rect 197 40592 99120 40872
rect 197 40192 99991 40592
rect 197 39912 99120 40192
rect 197 39512 99991 39912
rect 197 39232 99120 39512
rect 197 38832 99991 39232
rect 197 38552 99120 38832
rect 197 38152 99991 38552
rect 197 37872 99120 38152
rect 197 37472 99991 37872
rect 197 37192 99120 37472
rect 197 36792 99991 37192
rect 197 36512 99120 36792
rect 197 36112 99991 36512
rect 197 35832 99120 36112
rect 197 35432 99991 35832
rect 197 35152 99120 35432
rect 197 34752 99991 35152
rect 197 34472 99120 34752
rect 197 34072 99991 34472
rect 197 33792 99120 34072
rect 197 33392 99991 33792
rect 197 33112 99120 33392
rect 197 32712 99991 33112
rect 197 32432 99120 32712
rect 197 32032 99991 32432
rect 197 31752 99120 32032
rect 197 31352 99991 31752
rect 197 31072 99120 31352
rect 197 30672 99991 31072
rect 197 30392 99120 30672
rect 197 29992 99991 30392
rect 197 29712 99120 29992
rect 197 29312 99991 29712
rect 197 29032 99120 29312
rect 197 28632 99991 29032
rect 197 28352 99120 28632
rect 197 27952 99991 28352
rect 197 27672 99120 27952
rect 197 27272 99991 27672
rect 197 26992 99120 27272
rect 197 26592 99991 26992
rect 197 26312 99120 26592
rect 197 25912 99991 26312
rect 197 25632 99120 25912
rect 197 25232 99991 25632
rect 197 24952 99120 25232
rect 197 24552 99991 24952
rect 197 24272 99120 24552
rect 197 23872 99991 24272
rect 197 23592 99120 23872
rect 197 23192 99991 23592
rect 197 22912 99120 23192
rect 197 22512 99991 22912
rect 197 22232 99120 22512
rect 197 21832 99991 22232
rect 197 21552 99120 21832
rect 197 21152 99991 21552
rect 197 20872 99120 21152
rect 197 20472 99991 20872
rect 197 20192 99120 20472
rect 197 19792 99991 20192
rect 197 19512 99120 19792
rect 197 19112 99991 19512
rect 197 18832 99120 19112
rect 197 18432 99991 18832
rect 197 18152 99120 18432
rect 197 17752 99991 18152
rect 197 17472 99120 17752
rect 197 17072 99991 17472
rect 197 16792 99120 17072
rect 197 16392 99991 16792
rect 197 16112 99120 16392
rect 197 15712 99991 16112
rect 197 15432 99120 15712
rect 197 15032 99991 15432
rect 197 14752 99120 15032
rect 197 14352 99991 14752
rect 197 14072 99120 14352
rect 197 13672 99991 14072
rect 197 13392 99120 13672
rect 197 12992 99991 13392
rect 197 12712 99120 12992
rect 197 12312 99991 12712
rect 197 12032 99120 12312
rect 197 11632 99991 12032
rect 197 11352 99120 11632
rect 197 10952 99991 11352
rect 197 10672 99120 10952
rect 197 10272 99991 10672
rect 197 9992 99120 10272
rect 197 9592 99991 9992
rect 197 9312 99120 9592
rect 197 8912 99991 9312
rect 197 8632 99120 8912
rect 197 8232 99991 8632
rect 197 7952 99120 8232
rect 197 7552 99991 7952
rect 197 7272 99120 7552
rect 197 6872 99991 7272
rect 197 6592 99120 6872
rect 197 1395 99991 6592
<< metal4 >>
rect 1794 2128 2414 97424
rect 19794 2128 20414 97424
rect 37794 2128 38414 97424
rect 55794 2128 56414 97424
rect 73794 2128 74414 97424
rect 91794 2128 92414 97424
<< obsm4 >>
rect 427 97504 98565 98837
rect 427 2048 1714 97504
rect 2494 2048 19714 97504
rect 20494 2048 37714 97504
rect 38494 2048 55714 97504
rect 56494 2048 73714 97504
rect 74494 2048 91714 97504
rect 92494 2048 98565 97504
rect 427 1395 98565 2048
<< labels >>
rlabel metal4 s 19794 2128 20414 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 55794 2128 56414 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 91794 2128 92414 97424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1794 2128 2414 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 37794 2128 38414 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 73794 2128 74414 97424 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 99200 6672 100000 6792 6 a[0]
port 3 nsew signal input
rlabel metal3 s 99200 13472 100000 13592 6 a[10]
port 4 nsew signal input
rlabel metal3 s 99200 14152 100000 14272 6 a[11]
port 5 nsew signal input
rlabel metal3 s 99200 14832 100000 14952 6 a[12]
port 6 nsew signal input
rlabel metal3 s 99200 15512 100000 15632 6 a[13]
port 7 nsew signal input
rlabel metal3 s 99200 16192 100000 16312 6 a[14]
port 8 nsew signal input
rlabel metal3 s 99200 16872 100000 16992 6 a[15]
port 9 nsew signal input
rlabel metal3 s 99200 17552 100000 17672 6 a[16]
port 10 nsew signal input
rlabel metal3 s 99200 18232 100000 18352 6 a[17]
port 11 nsew signal input
rlabel metal3 s 99200 18912 100000 19032 6 a[18]
port 12 nsew signal input
rlabel metal3 s 99200 19592 100000 19712 6 a[19]
port 13 nsew signal input
rlabel metal3 s 99200 7352 100000 7472 6 a[1]
port 14 nsew signal input
rlabel metal3 s 99200 20272 100000 20392 6 a[20]
port 15 nsew signal input
rlabel metal3 s 99200 20952 100000 21072 6 a[21]
port 16 nsew signal input
rlabel metal3 s 99200 21632 100000 21752 6 a[22]
port 17 nsew signal input
rlabel metal3 s 99200 22312 100000 22432 6 a[23]
port 18 nsew signal input
rlabel metal3 s 99200 22992 100000 23112 6 a[24]
port 19 nsew signal input
rlabel metal3 s 99200 23672 100000 23792 6 a[25]
port 20 nsew signal input
rlabel metal3 s 99200 24352 100000 24472 6 a[26]
port 21 nsew signal input
rlabel metal3 s 99200 25032 100000 25152 6 a[27]
port 22 nsew signal input
rlabel metal3 s 99200 25712 100000 25832 6 a[28]
port 23 nsew signal input
rlabel metal3 s 99200 26392 100000 26512 6 a[29]
port 24 nsew signal input
rlabel metal3 s 99200 8032 100000 8152 6 a[2]
port 25 nsew signal input
rlabel metal3 s 99200 27072 100000 27192 6 a[30]
port 26 nsew signal input
rlabel metal3 s 99200 27752 100000 27872 6 a[31]
port 27 nsew signal input
rlabel metal3 s 99200 28432 100000 28552 6 a[32]
port 28 nsew signal input
rlabel metal3 s 99200 29112 100000 29232 6 a[33]
port 29 nsew signal input
rlabel metal3 s 99200 29792 100000 29912 6 a[34]
port 30 nsew signal input
rlabel metal3 s 99200 30472 100000 30592 6 a[35]
port 31 nsew signal input
rlabel metal3 s 99200 31152 100000 31272 6 a[36]
port 32 nsew signal input
rlabel metal3 s 99200 31832 100000 31952 6 a[37]
port 33 nsew signal input
rlabel metal3 s 99200 32512 100000 32632 6 a[38]
port 34 nsew signal input
rlabel metal3 s 99200 33192 100000 33312 6 a[39]
port 35 nsew signal input
rlabel metal3 s 99200 8712 100000 8832 6 a[3]
port 36 nsew signal input
rlabel metal3 s 99200 33872 100000 33992 6 a[40]
port 37 nsew signal input
rlabel metal3 s 99200 34552 100000 34672 6 a[41]
port 38 nsew signal input
rlabel metal3 s 99200 35232 100000 35352 6 a[42]
port 39 nsew signal input
rlabel metal3 s 99200 35912 100000 36032 6 a[43]
port 40 nsew signal input
rlabel metal3 s 99200 36592 100000 36712 6 a[44]
port 41 nsew signal input
rlabel metal3 s 99200 37272 100000 37392 6 a[45]
port 42 nsew signal input
rlabel metal3 s 99200 37952 100000 38072 6 a[46]
port 43 nsew signal input
rlabel metal3 s 99200 38632 100000 38752 6 a[47]
port 44 nsew signal input
rlabel metal3 s 99200 39312 100000 39432 6 a[48]
port 45 nsew signal input
rlabel metal3 s 99200 39992 100000 40112 6 a[49]
port 46 nsew signal input
rlabel metal3 s 99200 9392 100000 9512 6 a[4]
port 47 nsew signal input
rlabel metal3 s 99200 40672 100000 40792 6 a[50]
port 48 nsew signal input
rlabel metal3 s 99200 41352 100000 41472 6 a[51]
port 49 nsew signal input
rlabel metal3 s 99200 42032 100000 42152 6 a[52]
port 50 nsew signal input
rlabel metal3 s 99200 42712 100000 42832 6 a[53]
port 51 nsew signal input
rlabel metal3 s 99200 43392 100000 43512 6 a[54]
port 52 nsew signal input
rlabel metal3 s 99200 44072 100000 44192 6 a[55]
port 53 nsew signal input
rlabel metal3 s 99200 44752 100000 44872 6 a[56]
port 54 nsew signal input
rlabel metal3 s 99200 45432 100000 45552 6 a[57]
port 55 nsew signal input
rlabel metal3 s 99200 46112 100000 46232 6 a[58]
port 56 nsew signal input
rlabel metal3 s 99200 46792 100000 46912 6 a[59]
port 57 nsew signal input
rlabel metal3 s 99200 10072 100000 10192 6 a[5]
port 58 nsew signal input
rlabel metal3 s 99200 47472 100000 47592 6 a[60]
port 59 nsew signal input
rlabel metal3 s 99200 48152 100000 48272 6 a[61]
port 60 nsew signal input
rlabel metal3 s 99200 48832 100000 48952 6 a[62]
port 61 nsew signal input
rlabel metal3 s 99200 49512 100000 49632 6 a[63]
port 62 nsew signal input
rlabel metal3 s 99200 10752 100000 10872 6 a[6]
port 63 nsew signal input
rlabel metal3 s 99200 11432 100000 11552 6 a[7]
port 64 nsew signal input
rlabel metal3 s 99200 12112 100000 12232 6 a[8]
port 65 nsew signal input
rlabel metal3 s 99200 12792 100000 12912 6 a[9]
port 66 nsew signal input
rlabel metal3 s 99200 50192 100000 50312 6 b[0]
port 67 nsew signal input
rlabel metal3 s 99200 56992 100000 57112 6 b[10]
port 68 nsew signal input
rlabel metal3 s 99200 57672 100000 57792 6 b[11]
port 69 nsew signal input
rlabel metal3 s 99200 58352 100000 58472 6 b[12]
port 70 nsew signal input
rlabel metal3 s 99200 59032 100000 59152 6 b[13]
port 71 nsew signal input
rlabel metal3 s 99200 59712 100000 59832 6 b[14]
port 72 nsew signal input
rlabel metal3 s 99200 60392 100000 60512 6 b[15]
port 73 nsew signal input
rlabel metal3 s 99200 61072 100000 61192 6 b[16]
port 74 nsew signal input
rlabel metal3 s 99200 61752 100000 61872 6 b[17]
port 75 nsew signal input
rlabel metal3 s 99200 62432 100000 62552 6 b[18]
port 76 nsew signal input
rlabel metal3 s 99200 63112 100000 63232 6 b[19]
port 77 nsew signal input
rlabel metal3 s 99200 50872 100000 50992 6 b[1]
port 78 nsew signal input
rlabel metal3 s 99200 63792 100000 63912 6 b[20]
port 79 nsew signal input
rlabel metal3 s 99200 64472 100000 64592 6 b[21]
port 80 nsew signal input
rlabel metal3 s 99200 65152 100000 65272 6 b[22]
port 81 nsew signal input
rlabel metal3 s 99200 65832 100000 65952 6 b[23]
port 82 nsew signal input
rlabel metal3 s 99200 66512 100000 66632 6 b[24]
port 83 nsew signal input
rlabel metal3 s 99200 67192 100000 67312 6 b[25]
port 84 nsew signal input
rlabel metal3 s 99200 67872 100000 67992 6 b[26]
port 85 nsew signal input
rlabel metal3 s 99200 68552 100000 68672 6 b[27]
port 86 nsew signal input
rlabel metal3 s 99200 69232 100000 69352 6 b[28]
port 87 nsew signal input
rlabel metal3 s 99200 69912 100000 70032 6 b[29]
port 88 nsew signal input
rlabel metal3 s 99200 51552 100000 51672 6 b[2]
port 89 nsew signal input
rlabel metal3 s 99200 70592 100000 70712 6 b[30]
port 90 nsew signal input
rlabel metal3 s 99200 71272 100000 71392 6 b[31]
port 91 nsew signal input
rlabel metal3 s 99200 71952 100000 72072 6 b[32]
port 92 nsew signal input
rlabel metal3 s 99200 72632 100000 72752 6 b[33]
port 93 nsew signal input
rlabel metal3 s 99200 73312 100000 73432 6 b[34]
port 94 nsew signal input
rlabel metal3 s 99200 73992 100000 74112 6 b[35]
port 95 nsew signal input
rlabel metal3 s 99200 74672 100000 74792 6 b[36]
port 96 nsew signal input
rlabel metal3 s 99200 75352 100000 75472 6 b[37]
port 97 nsew signal input
rlabel metal3 s 99200 76032 100000 76152 6 b[38]
port 98 nsew signal input
rlabel metal3 s 99200 76712 100000 76832 6 b[39]
port 99 nsew signal input
rlabel metal3 s 99200 52232 100000 52352 6 b[3]
port 100 nsew signal input
rlabel metal3 s 99200 77392 100000 77512 6 b[40]
port 101 nsew signal input
rlabel metal3 s 99200 78072 100000 78192 6 b[41]
port 102 nsew signal input
rlabel metal3 s 99200 78752 100000 78872 6 b[42]
port 103 nsew signal input
rlabel metal3 s 99200 79432 100000 79552 6 b[43]
port 104 nsew signal input
rlabel metal3 s 99200 80112 100000 80232 6 b[44]
port 105 nsew signal input
rlabel metal3 s 99200 80792 100000 80912 6 b[45]
port 106 nsew signal input
rlabel metal3 s 99200 81472 100000 81592 6 b[46]
port 107 nsew signal input
rlabel metal3 s 99200 82152 100000 82272 6 b[47]
port 108 nsew signal input
rlabel metal3 s 99200 82832 100000 82952 6 b[48]
port 109 nsew signal input
rlabel metal3 s 99200 83512 100000 83632 6 b[49]
port 110 nsew signal input
rlabel metal3 s 99200 52912 100000 53032 6 b[4]
port 111 nsew signal input
rlabel metal3 s 99200 84192 100000 84312 6 b[50]
port 112 nsew signal input
rlabel metal3 s 99200 84872 100000 84992 6 b[51]
port 113 nsew signal input
rlabel metal3 s 99200 85552 100000 85672 6 b[52]
port 114 nsew signal input
rlabel metal3 s 99200 86232 100000 86352 6 b[53]
port 115 nsew signal input
rlabel metal3 s 99200 86912 100000 87032 6 b[54]
port 116 nsew signal input
rlabel metal3 s 99200 87592 100000 87712 6 b[55]
port 117 nsew signal input
rlabel metal3 s 99200 88272 100000 88392 6 b[56]
port 118 nsew signal input
rlabel metal3 s 99200 88952 100000 89072 6 b[57]
port 119 nsew signal input
rlabel metal3 s 99200 89632 100000 89752 6 b[58]
port 120 nsew signal input
rlabel metal3 s 99200 90312 100000 90432 6 b[59]
port 121 nsew signal input
rlabel metal3 s 99200 53592 100000 53712 6 b[5]
port 122 nsew signal input
rlabel metal3 s 99200 90992 100000 91112 6 b[60]
port 123 nsew signal input
rlabel metal3 s 99200 91672 100000 91792 6 b[61]
port 124 nsew signal input
rlabel metal3 s 99200 92352 100000 92472 6 b[62]
port 125 nsew signal input
rlabel metal3 s 99200 93032 100000 93152 6 b[63]
port 126 nsew signal input
rlabel metal3 s 99200 54272 100000 54392 6 b[6]
port 127 nsew signal input
rlabel metal3 s 99200 54952 100000 55072 6 b[7]
port 128 nsew signal input
rlabel metal3 s 99200 55632 100000 55752 6 b[8]
port 129 nsew signal input
rlabel metal3 s 99200 56312 100000 56432 6 b[9]
port 130 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 c[0]
port 131 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 c[100]
port 132 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 c[101]
port 133 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 c[102]
port 134 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 c[103]
port 135 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 c[104]
port 136 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 c[105]
port 137 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 c[106]
port 138 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 c[107]
port 139 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 c[108]
port 140 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 c[109]
port 141 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 c[10]
port 142 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 c[110]
port 143 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 c[111]
port 144 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 c[112]
port 145 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 c[113]
port 146 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 c[114]
port 147 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 c[115]
port 148 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 c[116]
port 149 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 c[117]
port 150 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 c[118]
port 151 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 c[119]
port 152 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 c[11]
port 153 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 c[120]
port 154 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 c[121]
port 155 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 c[122]
port 156 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 c[123]
port 157 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 c[124]
port 158 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 c[125]
port 159 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 c[126]
port 160 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 c[127]
port 161 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 c[12]
port 162 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 c[13]
port 163 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 c[14]
port 164 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 c[15]
port 165 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 c[16]
port 166 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 c[17]
port 167 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 c[18]
port 168 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 c[19]
port 169 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 c[1]
port 170 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 c[20]
port 171 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 c[21]
port 172 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 c[22]
port 173 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 c[23]
port 174 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 c[24]
port 175 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 c[25]
port 176 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 c[26]
port 177 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 c[27]
port 178 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 c[28]
port 179 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 c[29]
port 180 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 c[2]
port 181 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 c[30]
port 182 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 c[31]
port 183 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 c[32]
port 184 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 c[33]
port 185 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 c[34]
port 186 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 c[35]
port 187 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 c[36]
port 188 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 c[37]
port 189 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 c[38]
port 190 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 c[39]
port 191 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 c[3]
port 192 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 c[40]
port 193 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 c[41]
port 194 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 c[42]
port 195 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 c[43]
port 196 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 c[44]
port 197 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 c[45]
port 198 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 c[46]
port 199 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 c[47]
port 200 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 c[48]
port 201 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 c[49]
port 202 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 c[4]
port 203 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 c[50]
port 204 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 c[51]
port 205 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 c[52]
port 206 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 c[53]
port 207 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 c[54]
port 208 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 c[55]
port 209 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 c[56]
port 210 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 c[57]
port 211 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 c[58]
port 212 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 c[59]
port 213 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 c[5]
port 214 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 c[60]
port 215 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 c[61]
port 216 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 c[62]
port 217 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 c[63]
port 218 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 c[64]
port 219 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 c[65]
port 220 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 c[66]
port 221 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 c[67]
port 222 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 c[68]
port 223 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 c[69]
port 224 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 c[6]
port 225 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 c[70]
port 226 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 c[71]
port 227 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 c[72]
port 228 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 c[73]
port 229 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 c[74]
port 230 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 c[75]
port 231 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 c[76]
port 232 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 c[77]
port 233 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 c[78]
port 234 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 c[79]
port 235 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 c[7]
port 236 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 c[80]
port 237 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 c[81]
port 238 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 c[82]
port 239 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 c[83]
port 240 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 c[84]
port 241 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 c[85]
port 242 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 c[86]
port 243 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 c[87]
port 244 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 c[88]
port 245 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 c[89]
port 246 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 c[8]
port 247 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 c[90]
port 248 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 c[91]
port 249 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 c[92]
port 250 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 c[93]
port 251 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 c[94]
port 252 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 c[95]
port 253 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 c[96]
port 254 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 c[97]
port 255 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 c[98]
port 256 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 c[99]
port 257 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 c[9]
port 258 nsew signal input
rlabel metal2 s 97446 99200 97502 100000 6 clk
port 259 nsew signal input
rlabel metal2 s 2502 99200 2558 100000 6 o[0]
port 260 nsew signal output
rlabel metal2 s 76102 99200 76158 100000 6 o[100]
port 261 nsew signal output
rlabel metal2 s 76838 99200 76894 100000 6 o[101]
port 262 nsew signal output
rlabel metal2 s 77574 99200 77630 100000 6 o[102]
port 263 nsew signal output
rlabel metal2 s 78310 99200 78366 100000 6 o[103]
port 264 nsew signal output
rlabel metal2 s 79046 99200 79102 100000 6 o[104]
port 265 nsew signal output
rlabel metal2 s 79782 99200 79838 100000 6 o[105]
port 266 nsew signal output
rlabel metal2 s 80518 99200 80574 100000 6 o[106]
port 267 nsew signal output
rlabel metal2 s 81254 99200 81310 100000 6 o[107]
port 268 nsew signal output
rlabel metal2 s 81990 99200 82046 100000 6 o[108]
port 269 nsew signal output
rlabel metal2 s 82726 99200 82782 100000 6 o[109]
port 270 nsew signal output
rlabel metal2 s 9862 99200 9918 100000 6 o[10]
port 271 nsew signal output
rlabel metal2 s 83462 99200 83518 100000 6 o[110]
port 272 nsew signal output
rlabel metal2 s 84198 99200 84254 100000 6 o[111]
port 273 nsew signal output
rlabel metal2 s 84934 99200 84990 100000 6 o[112]
port 274 nsew signal output
rlabel metal2 s 85670 99200 85726 100000 6 o[113]
port 275 nsew signal output
rlabel metal2 s 86406 99200 86462 100000 6 o[114]
port 276 nsew signal output
rlabel metal2 s 87142 99200 87198 100000 6 o[115]
port 277 nsew signal output
rlabel metal2 s 87878 99200 87934 100000 6 o[116]
port 278 nsew signal output
rlabel metal2 s 88614 99200 88670 100000 6 o[117]
port 279 nsew signal output
rlabel metal2 s 89350 99200 89406 100000 6 o[118]
port 280 nsew signal output
rlabel metal2 s 90086 99200 90142 100000 6 o[119]
port 281 nsew signal output
rlabel metal2 s 10598 99200 10654 100000 6 o[11]
port 282 nsew signal output
rlabel metal2 s 90822 99200 90878 100000 6 o[120]
port 283 nsew signal output
rlabel metal2 s 91558 99200 91614 100000 6 o[121]
port 284 nsew signal output
rlabel metal2 s 92294 99200 92350 100000 6 o[122]
port 285 nsew signal output
rlabel metal2 s 93030 99200 93086 100000 6 o[123]
port 286 nsew signal output
rlabel metal2 s 93766 99200 93822 100000 6 o[124]
port 287 nsew signal output
rlabel metal2 s 94502 99200 94558 100000 6 o[125]
port 288 nsew signal output
rlabel metal2 s 95238 99200 95294 100000 6 o[126]
port 289 nsew signal output
rlabel metal2 s 95974 99200 96030 100000 6 o[127]
port 290 nsew signal output
rlabel metal2 s 11334 99200 11390 100000 6 o[12]
port 291 nsew signal output
rlabel metal2 s 12070 99200 12126 100000 6 o[13]
port 292 nsew signal output
rlabel metal2 s 12806 99200 12862 100000 6 o[14]
port 293 nsew signal output
rlabel metal2 s 13542 99200 13598 100000 6 o[15]
port 294 nsew signal output
rlabel metal2 s 14278 99200 14334 100000 6 o[16]
port 295 nsew signal output
rlabel metal2 s 15014 99200 15070 100000 6 o[17]
port 296 nsew signal output
rlabel metal2 s 15750 99200 15806 100000 6 o[18]
port 297 nsew signal output
rlabel metal2 s 16486 99200 16542 100000 6 o[19]
port 298 nsew signal output
rlabel metal2 s 3238 99200 3294 100000 6 o[1]
port 299 nsew signal output
rlabel metal2 s 17222 99200 17278 100000 6 o[20]
port 300 nsew signal output
rlabel metal2 s 17958 99200 18014 100000 6 o[21]
port 301 nsew signal output
rlabel metal2 s 18694 99200 18750 100000 6 o[22]
port 302 nsew signal output
rlabel metal2 s 19430 99200 19486 100000 6 o[23]
port 303 nsew signal output
rlabel metal2 s 20166 99200 20222 100000 6 o[24]
port 304 nsew signal output
rlabel metal2 s 20902 99200 20958 100000 6 o[25]
port 305 nsew signal output
rlabel metal2 s 21638 99200 21694 100000 6 o[26]
port 306 nsew signal output
rlabel metal2 s 22374 99200 22430 100000 6 o[27]
port 307 nsew signal output
rlabel metal2 s 23110 99200 23166 100000 6 o[28]
port 308 nsew signal output
rlabel metal2 s 23846 99200 23902 100000 6 o[29]
port 309 nsew signal output
rlabel metal2 s 3974 99200 4030 100000 6 o[2]
port 310 nsew signal output
rlabel metal2 s 24582 99200 24638 100000 6 o[30]
port 311 nsew signal output
rlabel metal2 s 25318 99200 25374 100000 6 o[31]
port 312 nsew signal output
rlabel metal2 s 26054 99200 26110 100000 6 o[32]
port 313 nsew signal output
rlabel metal2 s 26790 99200 26846 100000 6 o[33]
port 314 nsew signal output
rlabel metal2 s 27526 99200 27582 100000 6 o[34]
port 315 nsew signal output
rlabel metal2 s 28262 99200 28318 100000 6 o[35]
port 316 nsew signal output
rlabel metal2 s 28998 99200 29054 100000 6 o[36]
port 317 nsew signal output
rlabel metal2 s 29734 99200 29790 100000 6 o[37]
port 318 nsew signal output
rlabel metal2 s 30470 99200 30526 100000 6 o[38]
port 319 nsew signal output
rlabel metal2 s 31206 99200 31262 100000 6 o[39]
port 320 nsew signal output
rlabel metal2 s 4710 99200 4766 100000 6 o[3]
port 321 nsew signal output
rlabel metal2 s 31942 99200 31998 100000 6 o[40]
port 322 nsew signal output
rlabel metal2 s 32678 99200 32734 100000 6 o[41]
port 323 nsew signal output
rlabel metal2 s 33414 99200 33470 100000 6 o[42]
port 324 nsew signal output
rlabel metal2 s 34150 99200 34206 100000 6 o[43]
port 325 nsew signal output
rlabel metal2 s 34886 99200 34942 100000 6 o[44]
port 326 nsew signal output
rlabel metal2 s 35622 99200 35678 100000 6 o[45]
port 327 nsew signal output
rlabel metal2 s 36358 99200 36414 100000 6 o[46]
port 328 nsew signal output
rlabel metal2 s 37094 99200 37150 100000 6 o[47]
port 329 nsew signal output
rlabel metal2 s 37830 99200 37886 100000 6 o[48]
port 330 nsew signal output
rlabel metal2 s 38566 99200 38622 100000 6 o[49]
port 331 nsew signal output
rlabel metal2 s 5446 99200 5502 100000 6 o[4]
port 332 nsew signal output
rlabel metal2 s 39302 99200 39358 100000 6 o[50]
port 333 nsew signal output
rlabel metal2 s 40038 99200 40094 100000 6 o[51]
port 334 nsew signal output
rlabel metal2 s 40774 99200 40830 100000 6 o[52]
port 335 nsew signal output
rlabel metal2 s 41510 99200 41566 100000 6 o[53]
port 336 nsew signal output
rlabel metal2 s 42246 99200 42302 100000 6 o[54]
port 337 nsew signal output
rlabel metal2 s 42982 99200 43038 100000 6 o[55]
port 338 nsew signal output
rlabel metal2 s 43718 99200 43774 100000 6 o[56]
port 339 nsew signal output
rlabel metal2 s 44454 99200 44510 100000 6 o[57]
port 340 nsew signal output
rlabel metal2 s 45190 99200 45246 100000 6 o[58]
port 341 nsew signal output
rlabel metal2 s 45926 99200 45982 100000 6 o[59]
port 342 nsew signal output
rlabel metal2 s 6182 99200 6238 100000 6 o[5]
port 343 nsew signal output
rlabel metal2 s 46662 99200 46718 100000 6 o[60]
port 344 nsew signal output
rlabel metal2 s 47398 99200 47454 100000 6 o[61]
port 345 nsew signal output
rlabel metal2 s 48134 99200 48190 100000 6 o[62]
port 346 nsew signal output
rlabel metal2 s 48870 99200 48926 100000 6 o[63]
port 347 nsew signal output
rlabel metal2 s 49606 99200 49662 100000 6 o[64]
port 348 nsew signal output
rlabel metal2 s 50342 99200 50398 100000 6 o[65]
port 349 nsew signal output
rlabel metal2 s 51078 99200 51134 100000 6 o[66]
port 350 nsew signal output
rlabel metal2 s 51814 99200 51870 100000 6 o[67]
port 351 nsew signal output
rlabel metal2 s 52550 99200 52606 100000 6 o[68]
port 352 nsew signal output
rlabel metal2 s 53286 99200 53342 100000 6 o[69]
port 353 nsew signal output
rlabel metal2 s 6918 99200 6974 100000 6 o[6]
port 354 nsew signal output
rlabel metal2 s 54022 99200 54078 100000 6 o[70]
port 355 nsew signal output
rlabel metal2 s 54758 99200 54814 100000 6 o[71]
port 356 nsew signal output
rlabel metal2 s 55494 99200 55550 100000 6 o[72]
port 357 nsew signal output
rlabel metal2 s 56230 99200 56286 100000 6 o[73]
port 358 nsew signal output
rlabel metal2 s 56966 99200 57022 100000 6 o[74]
port 359 nsew signal output
rlabel metal2 s 57702 99200 57758 100000 6 o[75]
port 360 nsew signal output
rlabel metal2 s 58438 99200 58494 100000 6 o[76]
port 361 nsew signal output
rlabel metal2 s 59174 99200 59230 100000 6 o[77]
port 362 nsew signal output
rlabel metal2 s 59910 99200 59966 100000 6 o[78]
port 363 nsew signal output
rlabel metal2 s 60646 99200 60702 100000 6 o[79]
port 364 nsew signal output
rlabel metal2 s 7654 99200 7710 100000 6 o[7]
port 365 nsew signal output
rlabel metal2 s 61382 99200 61438 100000 6 o[80]
port 366 nsew signal output
rlabel metal2 s 62118 99200 62174 100000 6 o[81]
port 367 nsew signal output
rlabel metal2 s 62854 99200 62910 100000 6 o[82]
port 368 nsew signal output
rlabel metal2 s 63590 99200 63646 100000 6 o[83]
port 369 nsew signal output
rlabel metal2 s 64326 99200 64382 100000 6 o[84]
port 370 nsew signal output
rlabel metal2 s 65062 99200 65118 100000 6 o[85]
port 371 nsew signal output
rlabel metal2 s 65798 99200 65854 100000 6 o[86]
port 372 nsew signal output
rlabel metal2 s 66534 99200 66590 100000 6 o[87]
port 373 nsew signal output
rlabel metal2 s 67270 99200 67326 100000 6 o[88]
port 374 nsew signal output
rlabel metal2 s 68006 99200 68062 100000 6 o[89]
port 375 nsew signal output
rlabel metal2 s 8390 99200 8446 100000 6 o[8]
port 376 nsew signal output
rlabel metal2 s 68742 99200 68798 100000 6 o[90]
port 377 nsew signal output
rlabel metal2 s 69478 99200 69534 100000 6 o[91]
port 378 nsew signal output
rlabel metal2 s 70214 99200 70270 100000 6 o[92]
port 379 nsew signal output
rlabel metal2 s 70950 99200 71006 100000 6 o[93]
port 380 nsew signal output
rlabel metal2 s 71686 99200 71742 100000 6 o[94]
port 381 nsew signal output
rlabel metal2 s 72422 99200 72478 100000 6 o[95]
port 382 nsew signal output
rlabel metal2 s 73158 99200 73214 100000 6 o[96]
port 383 nsew signal output
rlabel metal2 s 73894 99200 73950 100000 6 o[97]
port 384 nsew signal output
rlabel metal2 s 74630 99200 74686 100000 6 o[98]
port 385 nsew signal output
rlabel metal2 s 75366 99200 75422 100000 6 o[99]
port 386 nsew signal output
rlabel metal2 s 9126 99200 9182 100000 6 o[9]
port 387 nsew signal output
rlabel metal2 s 96710 99200 96766 100000 6 rst
port 388 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 35817042
string GDS_FILE /scratch/mpw7/caravel_user_project/openlane/multiply_add_64x64/runs/22_09_06_08_57/results/signoff/multiply_add_64x64.magic.gds
string GDS_START 295336
<< end >>

