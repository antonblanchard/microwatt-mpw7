magic
tech sky130A
magscale 1 2
timestamp 1670231968
<< obsli1 >>
rect 4048 20111 313444 177361
<< obsm1 >>
rect 658 76 314902 197464
<< metal2 >>
rect 5078 197072 5134 197472
rect 9954 197072 10010 197472
rect 14830 197072 14886 197472
rect 19706 197072 19762 197472
rect 24582 197072 24638 197472
rect 29458 197072 29514 197472
rect 34334 197072 34390 197472
rect 39210 197072 39266 197472
rect 44086 197072 44142 197472
rect 48962 197072 49018 197472
rect 53838 197072 53894 197472
rect 58714 197072 58770 197472
rect 63590 197072 63646 197472
rect 68466 197072 68522 197472
rect 73342 197072 73398 197472
rect 78218 197072 78274 197472
rect 83094 197072 83150 197472
rect 87970 197072 88026 197472
rect 92846 197072 92902 197472
rect 97722 197072 97778 197472
rect 102598 197072 102654 197472
rect 107474 197072 107530 197472
rect 112350 197072 112406 197472
rect 117226 197072 117282 197472
rect 122102 197072 122158 197472
rect 126978 197072 127034 197472
rect 131854 197072 131910 197472
rect 136730 197072 136786 197472
rect 141606 197072 141662 197472
rect 146482 197072 146538 197472
rect 151358 197072 151414 197472
rect 156234 197072 156290 197472
rect 161110 197072 161166 197472
rect 165986 197072 166042 197472
rect 170862 197072 170918 197472
rect 175738 197072 175794 197472
rect 180614 197072 180670 197472
rect 185490 197072 185546 197472
rect 190366 197072 190422 197472
rect 195242 197072 195298 197472
rect 200118 197072 200174 197472
rect 204994 197072 205050 197472
rect 209870 197072 209926 197472
rect 214746 197072 214802 197472
rect 219622 197072 219678 197472
rect 224498 197072 224554 197472
rect 229374 197072 229430 197472
rect 234250 197072 234306 197472
rect 239126 197072 239182 197472
rect 244002 197072 244058 197472
rect 248878 197072 248934 197472
rect 253754 197072 253810 197472
rect 258630 197072 258686 197472
rect 263506 197072 263562 197472
rect 268382 197072 268438 197472
rect 273258 197072 273314 197472
rect 278134 197072 278190 197472
rect 283010 197072 283066 197472
rect 287886 197072 287942 197472
rect 292762 197072 292818 197472
rect 297638 197072 297694 197472
rect 302514 197072 302570 197472
rect 307390 197072 307446 197472
rect 312266 197072 312322 197472
rect 5078 0 5134 400
rect 9954 0 10010 400
rect 14830 0 14886 400
rect 19706 0 19762 400
rect 24582 0 24638 400
rect 29458 0 29514 400
rect 34334 0 34390 400
rect 39210 0 39266 400
rect 44086 0 44142 400
rect 48962 0 49018 400
rect 53838 0 53894 400
rect 58714 0 58770 400
rect 63590 0 63646 400
rect 68466 0 68522 400
rect 73342 0 73398 400
rect 78218 0 78274 400
rect 83094 0 83150 400
rect 87970 0 88026 400
rect 92846 0 92902 400
rect 97722 0 97778 400
rect 102598 0 102654 400
rect 107474 0 107530 400
rect 112350 0 112406 400
rect 117226 0 117282 400
rect 122102 0 122158 400
rect 126978 0 127034 400
rect 131854 0 131910 400
rect 136730 0 136786 400
rect 141606 0 141662 400
rect 146482 0 146538 400
rect 151358 0 151414 400
rect 156234 0 156290 400
rect 161110 0 161166 400
rect 165986 0 166042 400
rect 170862 0 170918 400
rect 175738 0 175794 400
rect 180614 0 180670 400
rect 185490 0 185546 400
rect 190366 0 190422 400
rect 195242 0 195298 400
rect 200118 0 200174 400
rect 204994 0 205050 400
rect 209870 0 209926 400
rect 214746 0 214802 400
rect 219622 0 219678 400
rect 224498 0 224554 400
rect 229374 0 229430 400
rect 234250 0 234306 400
rect 239126 0 239182 400
rect 244002 0 244058 400
rect 248878 0 248934 400
rect 253754 0 253810 400
rect 258630 0 258686 400
rect 263506 0 263562 400
rect 268382 0 268438 400
rect 273258 0 273314 400
rect 278134 0 278190 400
rect 283010 0 283066 400
rect 287886 0 287942 400
rect 292762 0 292818 400
rect 297638 0 297694 400
rect 302514 0 302570 400
rect 307390 0 307446 400
rect 312266 0 312322 400
<< obsm2 >>
rect 664 197016 5022 197470
rect 5190 197016 9898 197470
rect 10066 197016 14774 197470
rect 14942 197016 19650 197470
rect 19818 197016 24526 197470
rect 24694 197016 29402 197470
rect 29570 197016 34278 197470
rect 34446 197016 39154 197470
rect 39322 197016 44030 197470
rect 44198 197016 48906 197470
rect 49074 197016 53782 197470
rect 53950 197016 58658 197470
rect 58826 197016 63534 197470
rect 63702 197016 68410 197470
rect 68578 197016 73286 197470
rect 73454 197016 78162 197470
rect 78330 197016 83038 197470
rect 83206 197016 87914 197470
rect 88082 197016 92790 197470
rect 92958 197016 97666 197470
rect 97834 197016 102542 197470
rect 102710 197016 107418 197470
rect 107586 197016 112294 197470
rect 112462 197016 117170 197470
rect 117338 197016 122046 197470
rect 122214 197016 126922 197470
rect 127090 197016 131798 197470
rect 131966 197016 136674 197470
rect 136842 197016 141550 197470
rect 141718 197016 146426 197470
rect 146594 197016 151302 197470
rect 151470 197016 156178 197470
rect 156346 197016 161054 197470
rect 161222 197016 165930 197470
rect 166098 197016 170806 197470
rect 170974 197016 175682 197470
rect 175850 197016 180558 197470
rect 180726 197016 185434 197470
rect 185602 197016 190310 197470
rect 190478 197016 195186 197470
rect 195354 197016 200062 197470
rect 200230 197016 204938 197470
rect 205106 197016 209814 197470
rect 209982 197016 214690 197470
rect 214858 197016 219566 197470
rect 219734 197016 224442 197470
rect 224610 197016 229318 197470
rect 229486 197016 234194 197470
rect 234362 197016 239070 197470
rect 239238 197016 243946 197470
rect 244114 197016 248822 197470
rect 248990 197016 253698 197470
rect 253866 197016 258574 197470
rect 258742 197016 263450 197470
rect 263618 197016 268326 197470
rect 268494 197016 273202 197470
rect 273370 197016 278078 197470
rect 278246 197016 282954 197470
rect 283122 197016 287830 197470
rect 287998 197016 292706 197470
rect 292874 197016 297582 197470
rect 297750 197016 302458 197470
rect 302626 197016 307334 197470
rect 307502 197016 312210 197470
rect 312378 197016 314896 197470
rect 664 456 314896 197016
rect 664 70 5022 456
rect 5190 70 9898 456
rect 10066 70 14774 456
rect 14942 70 19650 456
rect 19818 70 24526 456
rect 24694 70 29402 456
rect 29570 70 34278 456
rect 34446 70 39154 456
rect 39322 70 44030 456
rect 44198 70 48906 456
rect 49074 70 53782 456
rect 53950 70 58658 456
rect 58826 70 63534 456
rect 63702 70 68410 456
rect 68578 70 73286 456
rect 73454 70 78162 456
rect 78330 70 83038 456
rect 83206 70 87914 456
rect 88082 70 92790 456
rect 92958 70 97666 456
rect 97834 70 102542 456
rect 102710 70 107418 456
rect 107586 70 112294 456
rect 112462 70 117170 456
rect 117338 70 122046 456
rect 122214 70 126922 456
rect 127090 70 131798 456
rect 131966 70 136674 456
rect 136842 70 141550 456
rect 141718 70 146426 456
rect 146594 70 151302 456
rect 151470 70 156178 456
rect 156346 70 161054 456
rect 161222 70 165930 456
rect 166098 70 170806 456
rect 170974 70 175682 456
rect 175850 70 180558 456
rect 180726 70 185434 456
rect 185602 70 190310 456
rect 190478 70 195186 456
rect 195354 70 200062 456
rect 200230 70 204938 456
rect 205106 70 209814 456
rect 209982 70 214690 456
rect 214858 70 219566 456
rect 219734 70 224442 456
rect 224610 70 229318 456
rect 229486 70 234194 456
rect 234362 70 239070 456
rect 239238 70 243946 456
rect 244114 70 248822 456
rect 248990 70 253698 456
rect 253866 70 258574 456
rect 258742 70 263450 456
rect 263618 70 268326 456
rect 268494 70 273202 456
rect 273370 70 278078 456
rect 278246 70 282954 456
rect 283122 70 287830 456
rect 287998 70 292706 456
rect 292874 70 297582 456
rect 297750 70 302458 456
rect 302626 70 307334 456
rect 307502 70 312210 456
rect 312378 70 314896 456
<< metal3 >>
rect 317092 191088 317492 191208
rect 317092 180208 317492 180328
rect 317092 169328 317492 169448
rect 317092 158448 317492 158568
rect 317092 147568 317492 147688
rect 317092 136688 317492 136808
rect 317092 125808 317492 125928
rect 317092 114928 317492 115048
rect 317092 104048 317492 104168
rect 0 98608 400 98728
rect 317092 93168 317492 93288
rect 317092 82288 317492 82408
rect 317092 71408 317492 71528
rect 317092 60528 317492 60648
rect 317092 49648 317492 49768
rect 317092 38768 317492 38888
rect 317092 27888 317492 28008
rect 317092 17008 317492 17128
rect 317092 6128 317492 6248
<< obsm3 >>
rect 400 191288 317092 197437
rect 400 191008 317012 191288
rect 400 180408 317092 191008
rect 400 180128 317012 180408
rect 400 169528 317092 180128
rect 400 169248 317012 169528
rect 400 158648 317092 169248
rect 400 158368 317012 158648
rect 400 147768 317092 158368
rect 400 147488 317012 147768
rect 400 136888 317092 147488
rect 400 136608 317012 136888
rect 400 126008 317092 136608
rect 400 125728 317012 126008
rect 400 115128 317092 125728
rect 400 114848 317012 115128
rect 400 104248 317092 114848
rect 400 103968 317012 104248
rect 400 98808 317092 103968
rect 480 98528 317092 98808
rect 400 93368 317092 98528
rect 400 93088 317012 93368
rect 400 82488 317092 93088
rect 400 82208 317012 82488
rect 400 71608 317092 82208
rect 400 71328 317012 71608
rect 400 60728 317092 71328
rect 400 60448 317012 60728
rect 400 49848 317092 60448
rect 400 49568 317012 49848
rect 400 38968 317092 49568
rect 400 38688 317012 38968
rect 400 28088 317092 38688
rect 400 27808 317012 28088
rect 400 17208 317092 27808
rect 400 16928 317012 17208
rect 400 6328 317092 16928
rect 400 6048 317012 6328
rect 400 171 317092 6048
<< metal4 >>
rect 4738 20080 5358 177392
rect 22738 20080 23358 177392
rect 40738 20080 41358 177392
rect 58738 20080 59358 177392
rect 76738 20080 77358 177392
rect 94738 20080 95358 177392
rect 112738 20080 113358 177392
rect 130738 20080 131358 177392
rect 148738 20080 149358 177392
rect 166738 20080 167358 177392
rect 184738 20080 185358 177392
rect 202738 20080 203358 177392
rect 220738 20080 221358 177392
rect 238738 20080 239358 177392
rect 256738 20080 257358 177392
rect 274738 20080 275358 177392
rect 292738 20080 293358 177392
rect 310738 20080 311358 177392
<< obsm4 >>
rect 8523 177472 314029 197437
rect 8523 20000 22658 177472
rect 23438 20000 40658 177472
rect 41438 20000 58658 177472
rect 59438 20000 76658 177472
rect 77438 20000 94658 177472
rect 95438 20000 112658 177472
rect 113438 20000 130658 177472
rect 131438 20000 148658 177472
rect 149438 20000 166658 177472
rect 167438 20000 184658 177472
rect 185438 20000 202658 177472
rect 203438 20000 220658 177472
rect 221438 20000 238658 177472
rect 239438 20000 256658 177472
rect 257438 20000 274658 177472
rect 275438 20000 292658 177472
rect 293438 20000 310658 177472
rect 311438 20000 314029 177472
rect 8523 171 314029 20000
<< labels >>
rlabel metal3 s 317092 104048 317492 104168 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 317092 114928 317492 115048 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 317092 125808 317492 125928 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 317092 136688 317492 136808 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 317092 147568 317492 147688 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 317092 158448 317492 158568 6 A0[5]
port 6 nsew signal input
rlabel metal3 s 317092 169328 317492 169448 6 A0[6]
port 7 nsew signal input
rlabel metal3 s 317092 180208 317492 180328 6 A0[7]
port 8 nsew signal input
rlabel metal3 s 317092 191088 317492 191208 6 A0[8]
port 9 nsew signal input
rlabel metal3 s 0 98608 400 98728 6 CLK
port 10 nsew signal input
rlabel metal2 s 5078 0 5134 400 6 Di0[0]
port 11 nsew signal input
rlabel metal2 s 53838 0 53894 400 6 Di0[10]
port 12 nsew signal input
rlabel metal2 s 58714 0 58770 400 6 Di0[11]
port 13 nsew signal input
rlabel metal2 s 63590 0 63646 400 6 Di0[12]
port 14 nsew signal input
rlabel metal2 s 68466 0 68522 400 6 Di0[13]
port 15 nsew signal input
rlabel metal2 s 73342 0 73398 400 6 Di0[14]
port 16 nsew signal input
rlabel metal2 s 78218 0 78274 400 6 Di0[15]
port 17 nsew signal input
rlabel metal2 s 83094 0 83150 400 6 Di0[16]
port 18 nsew signal input
rlabel metal2 s 87970 0 88026 400 6 Di0[17]
port 19 nsew signal input
rlabel metal2 s 92846 0 92902 400 6 Di0[18]
port 20 nsew signal input
rlabel metal2 s 97722 0 97778 400 6 Di0[19]
port 21 nsew signal input
rlabel metal2 s 9954 0 10010 400 6 Di0[1]
port 22 nsew signal input
rlabel metal2 s 102598 0 102654 400 6 Di0[20]
port 23 nsew signal input
rlabel metal2 s 107474 0 107530 400 6 Di0[21]
port 24 nsew signal input
rlabel metal2 s 112350 0 112406 400 6 Di0[22]
port 25 nsew signal input
rlabel metal2 s 117226 0 117282 400 6 Di0[23]
port 26 nsew signal input
rlabel metal2 s 122102 0 122158 400 6 Di0[24]
port 27 nsew signal input
rlabel metal2 s 126978 0 127034 400 6 Di0[25]
port 28 nsew signal input
rlabel metal2 s 131854 0 131910 400 6 Di0[26]
port 29 nsew signal input
rlabel metal2 s 136730 0 136786 400 6 Di0[27]
port 30 nsew signal input
rlabel metal2 s 141606 0 141662 400 6 Di0[28]
port 31 nsew signal input
rlabel metal2 s 146482 0 146538 400 6 Di0[29]
port 32 nsew signal input
rlabel metal2 s 14830 0 14886 400 6 Di0[2]
port 33 nsew signal input
rlabel metal2 s 151358 0 151414 400 6 Di0[30]
port 34 nsew signal input
rlabel metal2 s 156234 0 156290 400 6 Di0[31]
port 35 nsew signal input
rlabel metal2 s 161110 0 161166 400 6 Di0[32]
port 36 nsew signal input
rlabel metal2 s 165986 0 166042 400 6 Di0[33]
port 37 nsew signal input
rlabel metal2 s 170862 0 170918 400 6 Di0[34]
port 38 nsew signal input
rlabel metal2 s 175738 0 175794 400 6 Di0[35]
port 39 nsew signal input
rlabel metal2 s 180614 0 180670 400 6 Di0[36]
port 40 nsew signal input
rlabel metal2 s 185490 0 185546 400 6 Di0[37]
port 41 nsew signal input
rlabel metal2 s 190366 0 190422 400 6 Di0[38]
port 42 nsew signal input
rlabel metal2 s 195242 0 195298 400 6 Di0[39]
port 43 nsew signal input
rlabel metal2 s 19706 0 19762 400 6 Di0[3]
port 44 nsew signal input
rlabel metal2 s 200118 0 200174 400 6 Di0[40]
port 45 nsew signal input
rlabel metal2 s 204994 0 205050 400 6 Di0[41]
port 46 nsew signal input
rlabel metal2 s 209870 0 209926 400 6 Di0[42]
port 47 nsew signal input
rlabel metal2 s 214746 0 214802 400 6 Di0[43]
port 48 nsew signal input
rlabel metal2 s 219622 0 219678 400 6 Di0[44]
port 49 nsew signal input
rlabel metal2 s 224498 0 224554 400 6 Di0[45]
port 50 nsew signal input
rlabel metal2 s 229374 0 229430 400 6 Di0[46]
port 51 nsew signal input
rlabel metal2 s 234250 0 234306 400 6 Di0[47]
port 52 nsew signal input
rlabel metal2 s 239126 0 239182 400 6 Di0[48]
port 53 nsew signal input
rlabel metal2 s 244002 0 244058 400 6 Di0[49]
port 54 nsew signal input
rlabel metal2 s 24582 0 24638 400 6 Di0[4]
port 55 nsew signal input
rlabel metal2 s 248878 0 248934 400 6 Di0[50]
port 56 nsew signal input
rlabel metal2 s 253754 0 253810 400 6 Di0[51]
port 57 nsew signal input
rlabel metal2 s 258630 0 258686 400 6 Di0[52]
port 58 nsew signal input
rlabel metal2 s 263506 0 263562 400 6 Di0[53]
port 59 nsew signal input
rlabel metal2 s 268382 0 268438 400 6 Di0[54]
port 60 nsew signal input
rlabel metal2 s 273258 0 273314 400 6 Di0[55]
port 61 nsew signal input
rlabel metal2 s 278134 0 278190 400 6 Di0[56]
port 62 nsew signal input
rlabel metal2 s 283010 0 283066 400 6 Di0[57]
port 63 nsew signal input
rlabel metal2 s 287886 0 287942 400 6 Di0[58]
port 64 nsew signal input
rlabel metal2 s 292762 0 292818 400 6 Di0[59]
port 65 nsew signal input
rlabel metal2 s 29458 0 29514 400 6 Di0[5]
port 66 nsew signal input
rlabel metal2 s 297638 0 297694 400 6 Di0[60]
port 67 nsew signal input
rlabel metal2 s 302514 0 302570 400 6 Di0[61]
port 68 nsew signal input
rlabel metal2 s 307390 0 307446 400 6 Di0[62]
port 69 nsew signal input
rlabel metal2 s 312266 0 312322 400 6 Di0[63]
port 70 nsew signal input
rlabel metal2 s 34334 0 34390 400 6 Di0[6]
port 71 nsew signal input
rlabel metal2 s 39210 0 39266 400 6 Di0[7]
port 72 nsew signal input
rlabel metal2 s 44086 0 44142 400 6 Di0[8]
port 73 nsew signal input
rlabel metal2 s 48962 0 49018 400 6 Di0[9]
port 74 nsew signal input
rlabel metal2 s 5078 197072 5134 197472 6 Do0[0]
port 75 nsew signal output
rlabel metal2 s 53838 197072 53894 197472 6 Do0[10]
port 76 nsew signal output
rlabel metal2 s 58714 197072 58770 197472 6 Do0[11]
port 77 nsew signal output
rlabel metal2 s 63590 197072 63646 197472 6 Do0[12]
port 78 nsew signal output
rlabel metal2 s 68466 197072 68522 197472 6 Do0[13]
port 79 nsew signal output
rlabel metal2 s 73342 197072 73398 197472 6 Do0[14]
port 80 nsew signal output
rlabel metal2 s 78218 197072 78274 197472 6 Do0[15]
port 81 nsew signal output
rlabel metal2 s 83094 197072 83150 197472 6 Do0[16]
port 82 nsew signal output
rlabel metal2 s 87970 197072 88026 197472 6 Do0[17]
port 83 nsew signal output
rlabel metal2 s 92846 197072 92902 197472 6 Do0[18]
port 84 nsew signal output
rlabel metal2 s 97722 197072 97778 197472 6 Do0[19]
port 85 nsew signal output
rlabel metal2 s 9954 197072 10010 197472 6 Do0[1]
port 86 nsew signal output
rlabel metal2 s 102598 197072 102654 197472 6 Do0[20]
port 87 nsew signal output
rlabel metal2 s 107474 197072 107530 197472 6 Do0[21]
port 88 nsew signal output
rlabel metal2 s 112350 197072 112406 197472 6 Do0[22]
port 89 nsew signal output
rlabel metal2 s 117226 197072 117282 197472 6 Do0[23]
port 90 nsew signal output
rlabel metal2 s 122102 197072 122158 197472 6 Do0[24]
port 91 nsew signal output
rlabel metal2 s 126978 197072 127034 197472 6 Do0[25]
port 92 nsew signal output
rlabel metal2 s 131854 197072 131910 197472 6 Do0[26]
port 93 nsew signal output
rlabel metal2 s 136730 197072 136786 197472 6 Do0[27]
port 94 nsew signal output
rlabel metal2 s 141606 197072 141662 197472 6 Do0[28]
port 95 nsew signal output
rlabel metal2 s 146482 197072 146538 197472 6 Do0[29]
port 96 nsew signal output
rlabel metal2 s 14830 197072 14886 197472 6 Do0[2]
port 97 nsew signal output
rlabel metal2 s 151358 197072 151414 197472 6 Do0[30]
port 98 nsew signal output
rlabel metal2 s 156234 197072 156290 197472 6 Do0[31]
port 99 nsew signal output
rlabel metal2 s 161110 197072 161166 197472 6 Do0[32]
port 100 nsew signal output
rlabel metal2 s 165986 197072 166042 197472 6 Do0[33]
port 101 nsew signal output
rlabel metal2 s 170862 197072 170918 197472 6 Do0[34]
port 102 nsew signal output
rlabel metal2 s 175738 197072 175794 197472 6 Do0[35]
port 103 nsew signal output
rlabel metal2 s 180614 197072 180670 197472 6 Do0[36]
port 104 nsew signal output
rlabel metal2 s 185490 197072 185546 197472 6 Do0[37]
port 105 nsew signal output
rlabel metal2 s 190366 197072 190422 197472 6 Do0[38]
port 106 nsew signal output
rlabel metal2 s 195242 197072 195298 197472 6 Do0[39]
port 107 nsew signal output
rlabel metal2 s 19706 197072 19762 197472 6 Do0[3]
port 108 nsew signal output
rlabel metal2 s 200118 197072 200174 197472 6 Do0[40]
port 109 nsew signal output
rlabel metal2 s 204994 197072 205050 197472 6 Do0[41]
port 110 nsew signal output
rlabel metal2 s 209870 197072 209926 197472 6 Do0[42]
port 111 nsew signal output
rlabel metal2 s 214746 197072 214802 197472 6 Do0[43]
port 112 nsew signal output
rlabel metal2 s 219622 197072 219678 197472 6 Do0[44]
port 113 nsew signal output
rlabel metal2 s 224498 197072 224554 197472 6 Do0[45]
port 114 nsew signal output
rlabel metal2 s 229374 197072 229430 197472 6 Do0[46]
port 115 nsew signal output
rlabel metal2 s 234250 197072 234306 197472 6 Do0[47]
port 116 nsew signal output
rlabel metal2 s 239126 197072 239182 197472 6 Do0[48]
port 117 nsew signal output
rlabel metal2 s 244002 197072 244058 197472 6 Do0[49]
port 118 nsew signal output
rlabel metal2 s 24582 197072 24638 197472 6 Do0[4]
port 119 nsew signal output
rlabel metal2 s 248878 197072 248934 197472 6 Do0[50]
port 120 nsew signal output
rlabel metal2 s 253754 197072 253810 197472 6 Do0[51]
port 121 nsew signal output
rlabel metal2 s 258630 197072 258686 197472 6 Do0[52]
port 122 nsew signal output
rlabel metal2 s 263506 197072 263562 197472 6 Do0[53]
port 123 nsew signal output
rlabel metal2 s 268382 197072 268438 197472 6 Do0[54]
port 124 nsew signal output
rlabel metal2 s 273258 197072 273314 197472 6 Do0[55]
port 125 nsew signal output
rlabel metal2 s 278134 197072 278190 197472 6 Do0[56]
port 126 nsew signal output
rlabel metal2 s 283010 197072 283066 197472 6 Do0[57]
port 127 nsew signal output
rlabel metal2 s 287886 197072 287942 197472 6 Do0[58]
port 128 nsew signal output
rlabel metal2 s 292762 197072 292818 197472 6 Do0[59]
port 129 nsew signal output
rlabel metal2 s 29458 197072 29514 197472 6 Do0[5]
port 130 nsew signal output
rlabel metal2 s 297638 197072 297694 197472 6 Do0[60]
port 131 nsew signal output
rlabel metal2 s 302514 197072 302570 197472 6 Do0[61]
port 132 nsew signal output
rlabel metal2 s 307390 197072 307446 197472 6 Do0[62]
port 133 nsew signal output
rlabel metal2 s 312266 197072 312322 197472 6 Do0[63]
port 134 nsew signal output
rlabel metal2 s 34334 197072 34390 197472 6 Do0[6]
port 135 nsew signal output
rlabel metal2 s 39210 197072 39266 197472 6 Do0[7]
port 136 nsew signal output
rlabel metal2 s 44086 197072 44142 197472 6 Do0[8]
port 137 nsew signal output
rlabel metal2 s 48962 197072 49018 197472 6 Do0[9]
port 138 nsew signal output
rlabel metal3 s 317092 6128 317492 6248 6 EN0
port 139 nsew signal input
rlabel metal4 s 22738 20080 23358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 58738 20080 59358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 94738 20080 95358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 130738 20080 131358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 166738 20080 167358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 202738 20080 203358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 238738 20080 239358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 274738 20080 275358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 310738 20080 311358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 4738 20080 5358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 40738 20080 41358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 76738 20080 77358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 112738 20080 113358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 148738 20080 149358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 184738 20080 185358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 220738 20080 221358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 256738 20080 257358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 292738 20080 293358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal3 s 317092 17008 317492 17128 6 WE0[0]
port 142 nsew signal input
rlabel metal3 s 317092 27888 317492 28008 6 WE0[1]
port 143 nsew signal input
rlabel metal3 s 317092 38768 317492 38888 6 WE0[2]
port 144 nsew signal input
rlabel metal3 s 317092 49648 317492 49768 6 WE0[3]
port 145 nsew signal input
rlabel metal3 s 317092 60528 317492 60648 6 WE0[4]
port 146 nsew signal input
rlabel metal3 s 317092 71408 317492 71528 6 WE0[5]
port 147 nsew signal input
rlabel metal3 s 317092 82288 317492 82408 6 WE0[6]
port 148 nsew signal input
rlabel metal3 s 317092 93168 317492 93288 6 WE0[7]
port 149 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 317492 197472
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 189301874
string GDS_FILE /mnt/dffram/build/512x64_DEFAULT/openlane/runs/RUN_2022.12.05_07.28.55/results/signoff/RAM512.magic.gds
string GDS_START 165654
<< end >>

