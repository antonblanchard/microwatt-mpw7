// This is the unpowered netlist.
module multiply_add_64x64 (clk,
    rst,
    a,
    b,
    c,
    o);
 input clk;
 input rst;
 input [63:0] a;
 input [63:0] b;
 input [127:0] c;
 output [127:0] o;

 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire clknet_leaf_0_clk;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire booth_b0_m0;
 wire booth_b0_m1;
 wire booth_b0_m10;
 wire booth_b0_m11;
 wire booth_b0_m12;
 wire booth_b0_m13;
 wire booth_b0_m14;
 wire booth_b0_m15;
 wire booth_b0_m16;
 wire booth_b0_m17;
 wire booth_b0_m18;
 wire booth_b0_m19;
 wire booth_b0_m2;
 wire booth_b0_m20;
 wire booth_b0_m21;
 wire booth_b0_m22;
 wire booth_b0_m23;
 wire booth_b0_m24;
 wire booth_b0_m25;
 wire booth_b0_m26;
 wire booth_b0_m27;
 wire booth_b0_m28;
 wire booth_b0_m29;
 wire booth_b0_m3;
 wire booth_b0_m30;
 wire booth_b0_m31;
 wire booth_b0_m32;
 wire booth_b0_m33;
 wire booth_b0_m34;
 wire booth_b0_m35;
 wire booth_b0_m36;
 wire booth_b0_m37;
 wire booth_b0_m38;
 wire booth_b0_m39;
 wire booth_b0_m4;
 wire booth_b0_m40;
 wire booth_b0_m41;
 wire booth_b0_m42;
 wire booth_b0_m43;
 wire booth_b0_m44;
 wire booth_b0_m45;
 wire booth_b0_m46;
 wire booth_b0_m47;
 wire booth_b0_m48;
 wire booth_b0_m49;
 wire booth_b0_m5;
 wire booth_b0_m50;
 wire booth_b0_m51;
 wire booth_b0_m52;
 wire booth_b0_m53;
 wire booth_b0_m54;
 wire booth_b0_m55;
 wire booth_b0_m56;
 wire booth_b0_m57;
 wire booth_b0_m58;
 wire booth_b0_m59;
 wire booth_b0_m6;
 wire booth_b0_m60;
 wire booth_b0_m61;
 wire booth_b0_m62;
 wire booth_b0_m63;
 wire booth_b0_m64;
 wire booth_b0_m7;
 wire booth_b0_m8;
 wire booth_b0_m9;
 wire booth_b10_m0;
 wire booth_b10_m1;
 wire booth_b10_m10;
 wire booth_b10_m11;
 wire booth_b10_m12;
 wire booth_b10_m13;
 wire booth_b10_m14;
 wire booth_b10_m15;
 wire booth_b10_m16;
 wire booth_b10_m17;
 wire booth_b10_m18;
 wire booth_b10_m19;
 wire booth_b10_m2;
 wire booth_b10_m20;
 wire booth_b10_m21;
 wire booth_b10_m22;
 wire booth_b10_m23;
 wire booth_b10_m24;
 wire booth_b10_m25;
 wire booth_b10_m26;
 wire booth_b10_m27;
 wire booth_b10_m28;
 wire booth_b10_m29;
 wire booth_b10_m3;
 wire booth_b10_m30;
 wire booth_b10_m31;
 wire booth_b10_m32;
 wire booth_b10_m33;
 wire booth_b10_m34;
 wire booth_b10_m35;
 wire booth_b10_m36;
 wire booth_b10_m37;
 wire booth_b10_m38;
 wire booth_b10_m39;
 wire booth_b10_m4;
 wire booth_b10_m40;
 wire booth_b10_m41;
 wire booth_b10_m42;
 wire booth_b10_m43;
 wire booth_b10_m44;
 wire booth_b10_m45;
 wire booth_b10_m46;
 wire booth_b10_m47;
 wire booth_b10_m48;
 wire booth_b10_m49;
 wire booth_b10_m5;
 wire booth_b10_m50;
 wire booth_b10_m51;
 wire booth_b10_m52;
 wire booth_b10_m53;
 wire booth_b10_m54;
 wire booth_b10_m55;
 wire booth_b10_m56;
 wire booth_b10_m57;
 wire booth_b10_m58;
 wire booth_b10_m59;
 wire booth_b10_m6;
 wire booth_b10_m60;
 wire booth_b10_m61;
 wire booth_b10_m62;
 wire booth_b10_m63;
 wire booth_b10_m64;
 wire booth_b10_m7;
 wire booth_b10_m8;
 wire booth_b10_m9;
 wire booth_b12_m0;
 wire booth_b12_m1;
 wire booth_b12_m10;
 wire booth_b12_m11;
 wire booth_b12_m12;
 wire booth_b12_m13;
 wire booth_b12_m14;
 wire booth_b12_m15;
 wire booth_b12_m16;
 wire booth_b12_m17;
 wire booth_b12_m18;
 wire booth_b12_m19;
 wire booth_b12_m2;
 wire booth_b12_m20;
 wire booth_b12_m21;
 wire booth_b12_m22;
 wire booth_b12_m23;
 wire booth_b12_m24;
 wire booth_b12_m25;
 wire booth_b12_m26;
 wire booth_b12_m27;
 wire booth_b12_m28;
 wire booth_b12_m29;
 wire booth_b12_m3;
 wire booth_b12_m30;
 wire booth_b12_m31;
 wire booth_b12_m32;
 wire booth_b12_m33;
 wire booth_b12_m34;
 wire booth_b12_m35;
 wire booth_b12_m36;
 wire booth_b12_m37;
 wire booth_b12_m38;
 wire booth_b12_m39;
 wire booth_b12_m4;
 wire booth_b12_m40;
 wire booth_b12_m41;
 wire booth_b12_m42;
 wire booth_b12_m43;
 wire booth_b12_m44;
 wire booth_b12_m45;
 wire booth_b12_m46;
 wire booth_b12_m47;
 wire booth_b12_m48;
 wire booth_b12_m49;
 wire booth_b12_m5;
 wire booth_b12_m50;
 wire booth_b12_m51;
 wire booth_b12_m52;
 wire booth_b12_m53;
 wire booth_b12_m54;
 wire booth_b12_m55;
 wire booth_b12_m56;
 wire booth_b12_m57;
 wire booth_b12_m58;
 wire booth_b12_m59;
 wire booth_b12_m6;
 wire booth_b12_m60;
 wire booth_b12_m61;
 wire booth_b12_m62;
 wire booth_b12_m63;
 wire booth_b12_m64;
 wire booth_b12_m7;
 wire booth_b12_m8;
 wire booth_b12_m9;
 wire booth_b14_m0;
 wire booth_b14_m1;
 wire booth_b14_m10;
 wire booth_b14_m11;
 wire booth_b14_m12;
 wire booth_b14_m13;
 wire booth_b14_m14;
 wire booth_b14_m15;
 wire booth_b14_m16;
 wire booth_b14_m17;
 wire booth_b14_m18;
 wire booth_b14_m19;
 wire booth_b14_m2;
 wire booth_b14_m20;
 wire booth_b14_m21;
 wire booth_b14_m22;
 wire booth_b14_m23;
 wire booth_b14_m24;
 wire booth_b14_m25;
 wire booth_b14_m26;
 wire booth_b14_m27;
 wire booth_b14_m28;
 wire booth_b14_m29;
 wire booth_b14_m3;
 wire booth_b14_m30;
 wire booth_b14_m31;
 wire booth_b14_m32;
 wire booth_b14_m33;
 wire booth_b14_m34;
 wire booth_b14_m35;
 wire booth_b14_m36;
 wire booth_b14_m37;
 wire booth_b14_m38;
 wire booth_b14_m39;
 wire booth_b14_m4;
 wire booth_b14_m40;
 wire booth_b14_m41;
 wire booth_b14_m42;
 wire booth_b14_m43;
 wire booth_b14_m44;
 wire booth_b14_m45;
 wire booth_b14_m46;
 wire booth_b14_m47;
 wire booth_b14_m48;
 wire booth_b14_m49;
 wire booth_b14_m5;
 wire booth_b14_m50;
 wire booth_b14_m51;
 wire booth_b14_m52;
 wire booth_b14_m53;
 wire booth_b14_m54;
 wire booth_b14_m55;
 wire booth_b14_m56;
 wire booth_b14_m57;
 wire booth_b14_m58;
 wire booth_b14_m59;
 wire booth_b14_m6;
 wire booth_b14_m60;
 wire booth_b14_m61;
 wire booth_b14_m62;
 wire booth_b14_m63;
 wire booth_b14_m64;
 wire booth_b14_m7;
 wire booth_b14_m8;
 wire booth_b14_m9;
 wire booth_b16_m0;
 wire booth_b16_m1;
 wire booth_b16_m10;
 wire booth_b16_m11;
 wire booth_b16_m12;
 wire booth_b16_m13;
 wire booth_b16_m14;
 wire booth_b16_m15;
 wire booth_b16_m16;
 wire booth_b16_m17;
 wire booth_b16_m18;
 wire booth_b16_m19;
 wire booth_b16_m2;
 wire booth_b16_m20;
 wire booth_b16_m21;
 wire booth_b16_m22;
 wire booth_b16_m23;
 wire booth_b16_m24;
 wire booth_b16_m25;
 wire booth_b16_m26;
 wire booth_b16_m27;
 wire booth_b16_m28;
 wire booth_b16_m29;
 wire booth_b16_m3;
 wire booth_b16_m30;
 wire booth_b16_m31;
 wire booth_b16_m32;
 wire booth_b16_m33;
 wire booth_b16_m34;
 wire booth_b16_m35;
 wire booth_b16_m36;
 wire booth_b16_m37;
 wire booth_b16_m38;
 wire booth_b16_m39;
 wire booth_b16_m4;
 wire booth_b16_m40;
 wire booth_b16_m41;
 wire booth_b16_m42;
 wire booth_b16_m43;
 wire booth_b16_m44;
 wire booth_b16_m45;
 wire booth_b16_m46;
 wire booth_b16_m47;
 wire booth_b16_m48;
 wire booth_b16_m49;
 wire booth_b16_m5;
 wire booth_b16_m50;
 wire booth_b16_m51;
 wire booth_b16_m52;
 wire booth_b16_m53;
 wire booth_b16_m54;
 wire booth_b16_m55;
 wire booth_b16_m56;
 wire booth_b16_m57;
 wire booth_b16_m58;
 wire booth_b16_m59;
 wire booth_b16_m6;
 wire booth_b16_m60;
 wire booth_b16_m61;
 wire booth_b16_m62;
 wire booth_b16_m63;
 wire booth_b16_m64;
 wire booth_b16_m7;
 wire booth_b16_m8;
 wire booth_b16_m9;
 wire booth_b18_m0;
 wire booth_b18_m1;
 wire booth_b18_m10;
 wire booth_b18_m11;
 wire booth_b18_m12;
 wire booth_b18_m13;
 wire booth_b18_m14;
 wire booth_b18_m15;
 wire booth_b18_m16;
 wire booth_b18_m17;
 wire booth_b18_m18;
 wire booth_b18_m19;
 wire booth_b18_m2;
 wire booth_b18_m20;
 wire booth_b18_m21;
 wire booth_b18_m22;
 wire booth_b18_m23;
 wire booth_b18_m24;
 wire booth_b18_m25;
 wire booth_b18_m26;
 wire booth_b18_m27;
 wire booth_b18_m28;
 wire booth_b18_m29;
 wire booth_b18_m3;
 wire booth_b18_m30;
 wire booth_b18_m31;
 wire booth_b18_m32;
 wire booth_b18_m33;
 wire booth_b18_m34;
 wire booth_b18_m35;
 wire booth_b18_m36;
 wire booth_b18_m37;
 wire booth_b18_m38;
 wire booth_b18_m39;
 wire booth_b18_m4;
 wire booth_b18_m40;
 wire booth_b18_m41;
 wire booth_b18_m42;
 wire booth_b18_m43;
 wire booth_b18_m44;
 wire booth_b18_m45;
 wire booth_b18_m46;
 wire booth_b18_m47;
 wire booth_b18_m48;
 wire booth_b18_m49;
 wire booth_b18_m5;
 wire booth_b18_m50;
 wire booth_b18_m51;
 wire booth_b18_m52;
 wire booth_b18_m53;
 wire booth_b18_m54;
 wire booth_b18_m55;
 wire booth_b18_m56;
 wire booth_b18_m57;
 wire booth_b18_m58;
 wire booth_b18_m59;
 wire booth_b18_m6;
 wire booth_b18_m60;
 wire booth_b18_m61;
 wire booth_b18_m62;
 wire booth_b18_m63;
 wire booth_b18_m64;
 wire booth_b18_m7;
 wire booth_b18_m8;
 wire booth_b18_m9;
 wire booth_b20_m0;
 wire booth_b20_m1;
 wire booth_b20_m10;
 wire booth_b20_m11;
 wire booth_b20_m12;
 wire booth_b20_m13;
 wire booth_b20_m14;
 wire booth_b20_m15;
 wire booth_b20_m16;
 wire booth_b20_m17;
 wire booth_b20_m18;
 wire booth_b20_m19;
 wire booth_b20_m2;
 wire booth_b20_m20;
 wire booth_b20_m21;
 wire booth_b20_m22;
 wire booth_b20_m23;
 wire booth_b20_m24;
 wire booth_b20_m25;
 wire booth_b20_m26;
 wire booth_b20_m27;
 wire booth_b20_m28;
 wire booth_b20_m29;
 wire booth_b20_m3;
 wire booth_b20_m30;
 wire booth_b20_m31;
 wire booth_b20_m32;
 wire booth_b20_m33;
 wire booth_b20_m34;
 wire booth_b20_m35;
 wire booth_b20_m36;
 wire booth_b20_m37;
 wire booth_b20_m38;
 wire booth_b20_m39;
 wire booth_b20_m4;
 wire booth_b20_m40;
 wire booth_b20_m41;
 wire booth_b20_m42;
 wire booth_b20_m43;
 wire booth_b20_m44;
 wire booth_b20_m45;
 wire booth_b20_m46;
 wire booth_b20_m47;
 wire booth_b20_m48;
 wire booth_b20_m49;
 wire booth_b20_m5;
 wire booth_b20_m50;
 wire booth_b20_m51;
 wire booth_b20_m52;
 wire booth_b20_m53;
 wire booth_b20_m54;
 wire booth_b20_m55;
 wire booth_b20_m56;
 wire booth_b20_m57;
 wire booth_b20_m58;
 wire booth_b20_m59;
 wire booth_b20_m6;
 wire booth_b20_m60;
 wire booth_b20_m61;
 wire booth_b20_m62;
 wire booth_b20_m63;
 wire booth_b20_m64;
 wire booth_b20_m7;
 wire booth_b20_m8;
 wire booth_b20_m9;
 wire booth_b22_m0;
 wire booth_b22_m1;
 wire booth_b22_m10;
 wire booth_b22_m11;
 wire booth_b22_m12;
 wire booth_b22_m13;
 wire booth_b22_m14;
 wire booth_b22_m15;
 wire booth_b22_m16;
 wire booth_b22_m17;
 wire booth_b22_m18;
 wire booth_b22_m19;
 wire booth_b22_m2;
 wire booth_b22_m20;
 wire booth_b22_m21;
 wire booth_b22_m22;
 wire booth_b22_m23;
 wire booth_b22_m24;
 wire booth_b22_m25;
 wire booth_b22_m26;
 wire booth_b22_m27;
 wire booth_b22_m28;
 wire booth_b22_m29;
 wire booth_b22_m3;
 wire booth_b22_m30;
 wire booth_b22_m31;
 wire booth_b22_m32;
 wire booth_b22_m33;
 wire booth_b22_m34;
 wire booth_b22_m35;
 wire booth_b22_m36;
 wire booth_b22_m37;
 wire booth_b22_m38;
 wire booth_b22_m39;
 wire booth_b22_m4;
 wire booth_b22_m40;
 wire booth_b22_m41;
 wire booth_b22_m42;
 wire booth_b22_m43;
 wire booth_b22_m44;
 wire booth_b22_m45;
 wire booth_b22_m46;
 wire booth_b22_m47;
 wire booth_b22_m48;
 wire booth_b22_m49;
 wire booth_b22_m5;
 wire booth_b22_m50;
 wire booth_b22_m51;
 wire booth_b22_m52;
 wire booth_b22_m53;
 wire booth_b22_m54;
 wire booth_b22_m55;
 wire booth_b22_m56;
 wire booth_b22_m57;
 wire booth_b22_m58;
 wire booth_b22_m59;
 wire booth_b22_m6;
 wire booth_b22_m60;
 wire booth_b22_m61;
 wire booth_b22_m62;
 wire booth_b22_m63;
 wire booth_b22_m64;
 wire booth_b22_m7;
 wire booth_b22_m8;
 wire booth_b22_m9;
 wire booth_b24_m0;
 wire booth_b24_m1;
 wire booth_b24_m10;
 wire booth_b24_m11;
 wire booth_b24_m12;
 wire booth_b24_m13;
 wire booth_b24_m14;
 wire booth_b24_m15;
 wire booth_b24_m16;
 wire booth_b24_m17;
 wire booth_b24_m18;
 wire booth_b24_m19;
 wire booth_b24_m2;
 wire booth_b24_m20;
 wire booth_b24_m21;
 wire booth_b24_m22;
 wire booth_b24_m23;
 wire booth_b24_m24;
 wire booth_b24_m25;
 wire booth_b24_m26;
 wire booth_b24_m27;
 wire booth_b24_m28;
 wire booth_b24_m29;
 wire booth_b24_m3;
 wire booth_b24_m30;
 wire booth_b24_m31;
 wire booth_b24_m32;
 wire booth_b24_m33;
 wire booth_b24_m34;
 wire booth_b24_m35;
 wire booth_b24_m36;
 wire booth_b24_m37;
 wire booth_b24_m38;
 wire booth_b24_m39;
 wire booth_b24_m4;
 wire booth_b24_m40;
 wire booth_b24_m41;
 wire booth_b24_m42;
 wire booth_b24_m43;
 wire booth_b24_m44;
 wire booth_b24_m45;
 wire booth_b24_m46;
 wire booth_b24_m47;
 wire booth_b24_m48;
 wire booth_b24_m49;
 wire booth_b24_m5;
 wire booth_b24_m50;
 wire booth_b24_m51;
 wire booth_b24_m52;
 wire booth_b24_m53;
 wire booth_b24_m54;
 wire booth_b24_m55;
 wire booth_b24_m56;
 wire booth_b24_m57;
 wire booth_b24_m58;
 wire booth_b24_m59;
 wire booth_b24_m6;
 wire booth_b24_m60;
 wire booth_b24_m61;
 wire booth_b24_m62;
 wire booth_b24_m63;
 wire booth_b24_m64;
 wire booth_b24_m7;
 wire booth_b24_m8;
 wire booth_b24_m9;
 wire booth_b26_m0;
 wire booth_b26_m1;
 wire booth_b26_m10;
 wire booth_b26_m11;
 wire booth_b26_m12;
 wire booth_b26_m13;
 wire booth_b26_m14;
 wire booth_b26_m15;
 wire booth_b26_m16;
 wire booth_b26_m17;
 wire booth_b26_m18;
 wire booth_b26_m19;
 wire booth_b26_m2;
 wire booth_b26_m20;
 wire booth_b26_m21;
 wire booth_b26_m22;
 wire booth_b26_m23;
 wire booth_b26_m24;
 wire booth_b26_m25;
 wire booth_b26_m26;
 wire booth_b26_m27;
 wire booth_b26_m28;
 wire booth_b26_m29;
 wire booth_b26_m3;
 wire booth_b26_m30;
 wire booth_b26_m31;
 wire booth_b26_m32;
 wire booth_b26_m33;
 wire booth_b26_m34;
 wire booth_b26_m35;
 wire booth_b26_m36;
 wire booth_b26_m37;
 wire booth_b26_m38;
 wire booth_b26_m39;
 wire booth_b26_m4;
 wire booth_b26_m40;
 wire booth_b26_m41;
 wire booth_b26_m42;
 wire booth_b26_m43;
 wire booth_b26_m44;
 wire booth_b26_m45;
 wire booth_b26_m46;
 wire booth_b26_m47;
 wire booth_b26_m48;
 wire booth_b26_m49;
 wire booth_b26_m5;
 wire booth_b26_m50;
 wire booth_b26_m51;
 wire booth_b26_m52;
 wire booth_b26_m53;
 wire booth_b26_m54;
 wire booth_b26_m55;
 wire booth_b26_m56;
 wire booth_b26_m57;
 wire booth_b26_m58;
 wire booth_b26_m59;
 wire booth_b26_m6;
 wire booth_b26_m60;
 wire booth_b26_m61;
 wire booth_b26_m62;
 wire booth_b26_m63;
 wire booth_b26_m64;
 wire booth_b26_m7;
 wire booth_b26_m8;
 wire booth_b26_m9;
 wire booth_b28_m0;
 wire booth_b28_m1;
 wire booth_b28_m10;
 wire booth_b28_m11;
 wire booth_b28_m12;
 wire booth_b28_m13;
 wire booth_b28_m14;
 wire booth_b28_m15;
 wire booth_b28_m16;
 wire booth_b28_m17;
 wire booth_b28_m18;
 wire booth_b28_m19;
 wire booth_b28_m2;
 wire booth_b28_m20;
 wire booth_b28_m21;
 wire booth_b28_m22;
 wire booth_b28_m23;
 wire booth_b28_m24;
 wire booth_b28_m25;
 wire booth_b28_m26;
 wire booth_b28_m27;
 wire booth_b28_m28;
 wire booth_b28_m29;
 wire booth_b28_m3;
 wire booth_b28_m30;
 wire booth_b28_m31;
 wire booth_b28_m32;
 wire booth_b28_m33;
 wire booth_b28_m34;
 wire booth_b28_m35;
 wire booth_b28_m36;
 wire booth_b28_m37;
 wire booth_b28_m38;
 wire booth_b28_m39;
 wire booth_b28_m4;
 wire booth_b28_m40;
 wire booth_b28_m41;
 wire booth_b28_m42;
 wire booth_b28_m43;
 wire booth_b28_m44;
 wire booth_b28_m45;
 wire booth_b28_m46;
 wire booth_b28_m47;
 wire booth_b28_m48;
 wire booth_b28_m49;
 wire booth_b28_m5;
 wire booth_b28_m50;
 wire booth_b28_m51;
 wire booth_b28_m52;
 wire booth_b28_m53;
 wire booth_b28_m54;
 wire booth_b28_m55;
 wire booth_b28_m56;
 wire booth_b28_m57;
 wire booth_b28_m58;
 wire booth_b28_m59;
 wire booth_b28_m6;
 wire booth_b28_m60;
 wire booth_b28_m61;
 wire booth_b28_m62;
 wire booth_b28_m63;
 wire booth_b28_m64;
 wire booth_b28_m7;
 wire booth_b28_m8;
 wire booth_b28_m9;
 wire booth_b2_m0;
 wire booth_b2_m1;
 wire booth_b2_m10;
 wire booth_b2_m11;
 wire booth_b2_m12;
 wire booth_b2_m13;
 wire booth_b2_m14;
 wire booth_b2_m15;
 wire booth_b2_m16;
 wire booth_b2_m17;
 wire booth_b2_m18;
 wire booth_b2_m19;
 wire booth_b2_m2;
 wire booth_b2_m20;
 wire booth_b2_m21;
 wire booth_b2_m22;
 wire booth_b2_m23;
 wire booth_b2_m24;
 wire booth_b2_m25;
 wire booth_b2_m26;
 wire booth_b2_m27;
 wire booth_b2_m28;
 wire booth_b2_m29;
 wire booth_b2_m3;
 wire booth_b2_m30;
 wire booth_b2_m31;
 wire booth_b2_m32;
 wire booth_b2_m33;
 wire booth_b2_m34;
 wire booth_b2_m35;
 wire booth_b2_m36;
 wire booth_b2_m37;
 wire booth_b2_m38;
 wire booth_b2_m39;
 wire booth_b2_m4;
 wire booth_b2_m40;
 wire booth_b2_m41;
 wire booth_b2_m42;
 wire booth_b2_m43;
 wire booth_b2_m44;
 wire booth_b2_m45;
 wire booth_b2_m46;
 wire booth_b2_m47;
 wire booth_b2_m48;
 wire booth_b2_m49;
 wire booth_b2_m5;
 wire booth_b2_m50;
 wire booth_b2_m51;
 wire booth_b2_m52;
 wire booth_b2_m53;
 wire booth_b2_m54;
 wire booth_b2_m55;
 wire booth_b2_m56;
 wire booth_b2_m57;
 wire booth_b2_m58;
 wire booth_b2_m59;
 wire booth_b2_m6;
 wire booth_b2_m60;
 wire booth_b2_m61;
 wire booth_b2_m62;
 wire booth_b2_m63;
 wire booth_b2_m64;
 wire booth_b2_m7;
 wire booth_b2_m8;
 wire booth_b2_m9;
 wire booth_b30_m0;
 wire booth_b30_m1;
 wire booth_b30_m10;
 wire booth_b30_m11;
 wire booth_b30_m12;
 wire booth_b30_m13;
 wire booth_b30_m14;
 wire booth_b30_m15;
 wire booth_b30_m16;
 wire booth_b30_m17;
 wire booth_b30_m18;
 wire booth_b30_m19;
 wire booth_b30_m2;
 wire booth_b30_m20;
 wire booth_b30_m21;
 wire booth_b30_m22;
 wire booth_b30_m23;
 wire booth_b30_m24;
 wire booth_b30_m25;
 wire booth_b30_m26;
 wire booth_b30_m27;
 wire booth_b30_m28;
 wire booth_b30_m29;
 wire booth_b30_m3;
 wire booth_b30_m30;
 wire booth_b30_m31;
 wire booth_b30_m32;
 wire booth_b30_m33;
 wire booth_b30_m34;
 wire booth_b30_m35;
 wire booth_b30_m36;
 wire booth_b30_m37;
 wire booth_b30_m38;
 wire booth_b30_m39;
 wire booth_b30_m4;
 wire booth_b30_m40;
 wire booth_b30_m41;
 wire booth_b30_m42;
 wire booth_b30_m43;
 wire booth_b30_m44;
 wire booth_b30_m45;
 wire booth_b30_m46;
 wire booth_b30_m47;
 wire booth_b30_m48;
 wire booth_b30_m49;
 wire booth_b30_m5;
 wire booth_b30_m50;
 wire booth_b30_m51;
 wire booth_b30_m52;
 wire booth_b30_m53;
 wire booth_b30_m54;
 wire booth_b30_m55;
 wire booth_b30_m56;
 wire booth_b30_m57;
 wire booth_b30_m58;
 wire booth_b30_m59;
 wire booth_b30_m6;
 wire booth_b30_m60;
 wire booth_b30_m61;
 wire booth_b30_m62;
 wire booth_b30_m63;
 wire booth_b30_m64;
 wire booth_b30_m7;
 wire booth_b30_m8;
 wire booth_b30_m9;
 wire booth_b32_m0;
 wire booth_b32_m1;
 wire booth_b32_m10;
 wire booth_b32_m11;
 wire booth_b32_m12;
 wire booth_b32_m13;
 wire booth_b32_m14;
 wire booth_b32_m15;
 wire booth_b32_m16;
 wire booth_b32_m17;
 wire booth_b32_m18;
 wire booth_b32_m19;
 wire booth_b32_m2;
 wire booth_b32_m20;
 wire booth_b32_m21;
 wire booth_b32_m22;
 wire booth_b32_m23;
 wire booth_b32_m24;
 wire booth_b32_m25;
 wire booth_b32_m26;
 wire booth_b32_m27;
 wire booth_b32_m28;
 wire booth_b32_m29;
 wire booth_b32_m3;
 wire booth_b32_m30;
 wire booth_b32_m31;
 wire booth_b32_m32;
 wire booth_b32_m33;
 wire booth_b32_m34;
 wire booth_b32_m35;
 wire booth_b32_m36;
 wire booth_b32_m37;
 wire booth_b32_m38;
 wire booth_b32_m39;
 wire booth_b32_m4;
 wire booth_b32_m40;
 wire booth_b32_m41;
 wire booth_b32_m42;
 wire booth_b32_m43;
 wire booth_b32_m44;
 wire booth_b32_m45;
 wire booth_b32_m46;
 wire booth_b32_m47;
 wire booth_b32_m48;
 wire booth_b32_m49;
 wire booth_b32_m5;
 wire booth_b32_m50;
 wire booth_b32_m51;
 wire booth_b32_m52;
 wire booth_b32_m53;
 wire booth_b32_m54;
 wire booth_b32_m55;
 wire booth_b32_m56;
 wire booth_b32_m57;
 wire booth_b32_m58;
 wire booth_b32_m59;
 wire booth_b32_m6;
 wire booth_b32_m60;
 wire booth_b32_m61;
 wire booth_b32_m62;
 wire booth_b32_m63;
 wire booth_b32_m64;
 wire booth_b32_m7;
 wire booth_b32_m8;
 wire booth_b32_m9;
 wire booth_b34_m0;
 wire booth_b34_m1;
 wire booth_b34_m10;
 wire booth_b34_m11;
 wire booth_b34_m12;
 wire booth_b34_m13;
 wire booth_b34_m14;
 wire booth_b34_m15;
 wire booth_b34_m16;
 wire booth_b34_m17;
 wire booth_b34_m18;
 wire booth_b34_m19;
 wire booth_b34_m2;
 wire booth_b34_m20;
 wire booth_b34_m21;
 wire booth_b34_m22;
 wire booth_b34_m23;
 wire booth_b34_m24;
 wire booth_b34_m25;
 wire booth_b34_m26;
 wire booth_b34_m27;
 wire booth_b34_m28;
 wire booth_b34_m29;
 wire booth_b34_m3;
 wire booth_b34_m30;
 wire booth_b34_m31;
 wire booth_b34_m32;
 wire booth_b34_m33;
 wire booth_b34_m34;
 wire booth_b34_m35;
 wire booth_b34_m36;
 wire booth_b34_m37;
 wire booth_b34_m38;
 wire booth_b34_m39;
 wire booth_b34_m4;
 wire booth_b34_m40;
 wire booth_b34_m41;
 wire booth_b34_m42;
 wire booth_b34_m43;
 wire booth_b34_m44;
 wire booth_b34_m45;
 wire booth_b34_m46;
 wire booth_b34_m47;
 wire booth_b34_m48;
 wire booth_b34_m49;
 wire booth_b34_m5;
 wire booth_b34_m50;
 wire booth_b34_m51;
 wire booth_b34_m52;
 wire booth_b34_m53;
 wire booth_b34_m54;
 wire booth_b34_m55;
 wire booth_b34_m56;
 wire booth_b34_m57;
 wire booth_b34_m58;
 wire booth_b34_m59;
 wire booth_b34_m6;
 wire booth_b34_m60;
 wire booth_b34_m61;
 wire booth_b34_m62;
 wire booth_b34_m63;
 wire booth_b34_m64;
 wire booth_b34_m7;
 wire booth_b34_m8;
 wire booth_b34_m9;
 wire booth_b36_m0;
 wire booth_b36_m1;
 wire booth_b36_m10;
 wire booth_b36_m11;
 wire booth_b36_m12;
 wire booth_b36_m13;
 wire booth_b36_m14;
 wire booth_b36_m15;
 wire booth_b36_m16;
 wire booth_b36_m17;
 wire booth_b36_m18;
 wire booth_b36_m19;
 wire booth_b36_m2;
 wire booth_b36_m20;
 wire booth_b36_m21;
 wire booth_b36_m22;
 wire booth_b36_m23;
 wire booth_b36_m24;
 wire booth_b36_m25;
 wire booth_b36_m26;
 wire booth_b36_m27;
 wire booth_b36_m28;
 wire booth_b36_m29;
 wire booth_b36_m3;
 wire booth_b36_m30;
 wire booth_b36_m31;
 wire booth_b36_m32;
 wire booth_b36_m33;
 wire booth_b36_m34;
 wire booth_b36_m35;
 wire booth_b36_m36;
 wire booth_b36_m37;
 wire booth_b36_m38;
 wire booth_b36_m39;
 wire booth_b36_m4;
 wire booth_b36_m40;
 wire booth_b36_m41;
 wire booth_b36_m42;
 wire booth_b36_m43;
 wire booth_b36_m44;
 wire booth_b36_m45;
 wire booth_b36_m46;
 wire booth_b36_m47;
 wire booth_b36_m48;
 wire booth_b36_m49;
 wire booth_b36_m5;
 wire booth_b36_m50;
 wire booth_b36_m51;
 wire booth_b36_m52;
 wire booth_b36_m53;
 wire booth_b36_m54;
 wire booth_b36_m55;
 wire booth_b36_m56;
 wire booth_b36_m57;
 wire booth_b36_m58;
 wire booth_b36_m59;
 wire booth_b36_m6;
 wire booth_b36_m60;
 wire booth_b36_m61;
 wire booth_b36_m62;
 wire booth_b36_m63;
 wire booth_b36_m64;
 wire booth_b36_m7;
 wire booth_b36_m8;
 wire booth_b36_m9;
 wire booth_b38_m0;
 wire booth_b38_m1;
 wire booth_b38_m10;
 wire booth_b38_m11;
 wire booth_b38_m12;
 wire booth_b38_m13;
 wire booth_b38_m14;
 wire booth_b38_m15;
 wire booth_b38_m16;
 wire booth_b38_m17;
 wire booth_b38_m18;
 wire booth_b38_m19;
 wire booth_b38_m2;
 wire booth_b38_m20;
 wire booth_b38_m21;
 wire booth_b38_m22;
 wire booth_b38_m23;
 wire booth_b38_m24;
 wire booth_b38_m25;
 wire booth_b38_m26;
 wire booth_b38_m27;
 wire booth_b38_m28;
 wire booth_b38_m29;
 wire booth_b38_m3;
 wire booth_b38_m30;
 wire booth_b38_m31;
 wire booth_b38_m32;
 wire booth_b38_m33;
 wire booth_b38_m34;
 wire booth_b38_m35;
 wire booth_b38_m36;
 wire booth_b38_m37;
 wire booth_b38_m38;
 wire booth_b38_m39;
 wire booth_b38_m4;
 wire booth_b38_m40;
 wire booth_b38_m41;
 wire booth_b38_m42;
 wire booth_b38_m43;
 wire booth_b38_m44;
 wire booth_b38_m45;
 wire booth_b38_m46;
 wire booth_b38_m47;
 wire booth_b38_m48;
 wire booth_b38_m49;
 wire booth_b38_m5;
 wire booth_b38_m50;
 wire booth_b38_m51;
 wire booth_b38_m52;
 wire booth_b38_m53;
 wire booth_b38_m54;
 wire booth_b38_m55;
 wire booth_b38_m56;
 wire booth_b38_m57;
 wire booth_b38_m58;
 wire booth_b38_m59;
 wire booth_b38_m6;
 wire booth_b38_m60;
 wire booth_b38_m61;
 wire booth_b38_m62;
 wire booth_b38_m63;
 wire booth_b38_m64;
 wire booth_b38_m7;
 wire booth_b38_m8;
 wire booth_b38_m9;
 wire booth_b40_m0;
 wire booth_b40_m1;
 wire booth_b40_m10;
 wire booth_b40_m11;
 wire booth_b40_m12;
 wire booth_b40_m13;
 wire booth_b40_m14;
 wire booth_b40_m15;
 wire booth_b40_m16;
 wire booth_b40_m17;
 wire booth_b40_m18;
 wire booth_b40_m19;
 wire booth_b40_m2;
 wire booth_b40_m20;
 wire booth_b40_m21;
 wire booth_b40_m22;
 wire booth_b40_m23;
 wire booth_b40_m24;
 wire booth_b40_m25;
 wire booth_b40_m26;
 wire booth_b40_m27;
 wire booth_b40_m28;
 wire booth_b40_m29;
 wire booth_b40_m3;
 wire booth_b40_m30;
 wire booth_b40_m31;
 wire booth_b40_m32;
 wire booth_b40_m33;
 wire booth_b40_m34;
 wire booth_b40_m35;
 wire booth_b40_m36;
 wire booth_b40_m37;
 wire booth_b40_m38;
 wire booth_b40_m39;
 wire booth_b40_m4;
 wire booth_b40_m40;
 wire booth_b40_m41;
 wire booth_b40_m42;
 wire booth_b40_m43;
 wire booth_b40_m44;
 wire booth_b40_m45;
 wire booth_b40_m46;
 wire booth_b40_m47;
 wire booth_b40_m48;
 wire booth_b40_m49;
 wire booth_b40_m5;
 wire booth_b40_m50;
 wire booth_b40_m51;
 wire booth_b40_m52;
 wire booth_b40_m53;
 wire booth_b40_m54;
 wire booth_b40_m55;
 wire booth_b40_m56;
 wire booth_b40_m57;
 wire booth_b40_m58;
 wire booth_b40_m59;
 wire booth_b40_m6;
 wire booth_b40_m60;
 wire booth_b40_m61;
 wire booth_b40_m62;
 wire booth_b40_m63;
 wire booth_b40_m64;
 wire booth_b40_m7;
 wire booth_b40_m8;
 wire booth_b40_m9;
 wire booth_b42_m0;
 wire booth_b42_m1;
 wire booth_b42_m10;
 wire booth_b42_m11;
 wire booth_b42_m12;
 wire booth_b42_m13;
 wire booth_b42_m14;
 wire booth_b42_m15;
 wire booth_b42_m16;
 wire booth_b42_m17;
 wire booth_b42_m18;
 wire booth_b42_m19;
 wire booth_b42_m2;
 wire booth_b42_m20;
 wire booth_b42_m21;
 wire booth_b42_m22;
 wire booth_b42_m23;
 wire booth_b42_m24;
 wire booth_b42_m25;
 wire booth_b42_m26;
 wire booth_b42_m27;
 wire booth_b42_m28;
 wire booth_b42_m29;
 wire booth_b42_m3;
 wire booth_b42_m30;
 wire booth_b42_m31;
 wire booth_b42_m32;
 wire booth_b42_m33;
 wire booth_b42_m34;
 wire booth_b42_m35;
 wire booth_b42_m36;
 wire booth_b42_m37;
 wire booth_b42_m38;
 wire booth_b42_m39;
 wire booth_b42_m4;
 wire booth_b42_m40;
 wire booth_b42_m41;
 wire booth_b42_m42;
 wire booth_b42_m43;
 wire booth_b42_m44;
 wire booth_b42_m45;
 wire booth_b42_m46;
 wire booth_b42_m47;
 wire booth_b42_m48;
 wire booth_b42_m49;
 wire booth_b42_m5;
 wire booth_b42_m50;
 wire booth_b42_m51;
 wire booth_b42_m52;
 wire booth_b42_m53;
 wire booth_b42_m54;
 wire booth_b42_m55;
 wire booth_b42_m56;
 wire booth_b42_m57;
 wire booth_b42_m58;
 wire booth_b42_m59;
 wire booth_b42_m6;
 wire booth_b42_m60;
 wire booth_b42_m61;
 wire booth_b42_m62;
 wire booth_b42_m63;
 wire booth_b42_m64;
 wire booth_b42_m7;
 wire booth_b42_m8;
 wire booth_b42_m9;
 wire booth_b44_m0;
 wire booth_b44_m1;
 wire booth_b44_m10;
 wire booth_b44_m11;
 wire booth_b44_m12;
 wire booth_b44_m13;
 wire booth_b44_m14;
 wire booth_b44_m15;
 wire booth_b44_m16;
 wire booth_b44_m17;
 wire booth_b44_m18;
 wire booth_b44_m19;
 wire booth_b44_m2;
 wire booth_b44_m20;
 wire booth_b44_m21;
 wire booth_b44_m22;
 wire booth_b44_m23;
 wire booth_b44_m24;
 wire booth_b44_m25;
 wire booth_b44_m26;
 wire booth_b44_m27;
 wire booth_b44_m28;
 wire booth_b44_m29;
 wire booth_b44_m3;
 wire booth_b44_m30;
 wire booth_b44_m31;
 wire booth_b44_m32;
 wire booth_b44_m33;
 wire booth_b44_m34;
 wire booth_b44_m35;
 wire booth_b44_m36;
 wire booth_b44_m37;
 wire booth_b44_m38;
 wire booth_b44_m39;
 wire booth_b44_m4;
 wire booth_b44_m40;
 wire booth_b44_m41;
 wire booth_b44_m42;
 wire booth_b44_m43;
 wire booth_b44_m44;
 wire booth_b44_m45;
 wire booth_b44_m46;
 wire booth_b44_m47;
 wire booth_b44_m48;
 wire booth_b44_m49;
 wire booth_b44_m5;
 wire booth_b44_m50;
 wire booth_b44_m51;
 wire booth_b44_m52;
 wire booth_b44_m53;
 wire booth_b44_m54;
 wire booth_b44_m55;
 wire booth_b44_m56;
 wire booth_b44_m57;
 wire booth_b44_m58;
 wire booth_b44_m59;
 wire booth_b44_m6;
 wire booth_b44_m60;
 wire booth_b44_m61;
 wire booth_b44_m62;
 wire booth_b44_m63;
 wire booth_b44_m64;
 wire booth_b44_m7;
 wire booth_b44_m8;
 wire booth_b44_m9;
 wire booth_b46_m0;
 wire booth_b46_m1;
 wire booth_b46_m10;
 wire booth_b46_m11;
 wire booth_b46_m12;
 wire booth_b46_m13;
 wire booth_b46_m14;
 wire booth_b46_m15;
 wire booth_b46_m16;
 wire booth_b46_m17;
 wire booth_b46_m18;
 wire booth_b46_m19;
 wire booth_b46_m2;
 wire booth_b46_m20;
 wire booth_b46_m21;
 wire booth_b46_m22;
 wire booth_b46_m23;
 wire booth_b46_m24;
 wire booth_b46_m25;
 wire booth_b46_m26;
 wire booth_b46_m27;
 wire booth_b46_m28;
 wire booth_b46_m29;
 wire booth_b46_m3;
 wire booth_b46_m30;
 wire booth_b46_m31;
 wire booth_b46_m32;
 wire booth_b46_m33;
 wire booth_b46_m34;
 wire booth_b46_m35;
 wire booth_b46_m36;
 wire booth_b46_m37;
 wire booth_b46_m38;
 wire booth_b46_m39;
 wire booth_b46_m4;
 wire booth_b46_m40;
 wire booth_b46_m41;
 wire booth_b46_m42;
 wire booth_b46_m43;
 wire booth_b46_m44;
 wire booth_b46_m45;
 wire booth_b46_m46;
 wire booth_b46_m47;
 wire booth_b46_m48;
 wire booth_b46_m49;
 wire booth_b46_m5;
 wire booth_b46_m50;
 wire booth_b46_m51;
 wire booth_b46_m52;
 wire booth_b46_m53;
 wire booth_b46_m54;
 wire booth_b46_m55;
 wire booth_b46_m56;
 wire booth_b46_m57;
 wire booth_b46_m58;
 wire booth_b46_m59;
 wire booth_b46_m6;
 wire booth_b46_m60;
 wire booth_b46_m61;
 wire booth_b46_m62;
 wire booth_b46_m63;
 wire booth_b46_m64;
 wire booth_b46_m7;
 wire booth_b46_m8;
 wire booth_b46_m9;
 wire booth_b48_m0;
 wire booth_b48_m1;
 wire booth_b48_m10;
 wire booth_b48_m11;
 wire booth_b48_m12;
 wire booth_b48_m13;
 wire booth_b48_m14;
 wire booth_b48_m15;
 wire booth_b48_m16;
 wire booth_b48_m17;
 wire booth_b48_m18;
 wire booth_b48_m19;
 wire booth_b48_m2;
 wire booth_b48_m20;
 wire booth_b48_m21;
 wire booth_b48_m22;
 wire booth_b48_m23;
 wire booth_b48_m24;
 wire booth_b48_m25;
 wire booth_b48_m26;
 wire booth_b48_m27;
 wire booth_b48_m28;
 wire booth_b48_m29;
 wire booth_b48_m3;
 wire booth_b48_m30;
 wire booth_b48_m31;
 wire booth_b48_m32;
 wire booth_b48_m33;
 wire booth_b48_m34;
 wire booth_b48_m35;
 wire booth_b48_m36;
 wire booth_b48_m37;
 wire booth_b48_m38;
 wire booth_b48_m39;
 wire booth_b48_m4;
 wire booth_b48_m40;
 wire booth_b48_m41;
 wire booth_b48_m42;
 wire booth_b48_m43;
 wire booth_b48_m44;
 wire booth_b48_m45;
 wire booth_b48_m46;
 wire booth_b48_m47;
 wire booth_b48_m48;
 wire booth_b48_m49;
 wire booth_b48_m5;
 wire booth_b48_m50;
 wire booth_b48_m51;
 wire booth_b48_m52;
 wire booth_b48_m53;
 wire booth_b48_m54;
 wire booth_b48_m55;
 wire booth_b48_m56;
 wire booth_b48_m57;
 wire booth_b48_m58;
 wire booth_b48_m59;
 wire booth_b48_m6;
 wire booth_b48_m60;
 wire booth_b48_m61;
 wire booth_b48_m62;
 wire booth_b48_m63;
 wire booth_b48_m64;
 wire booth_b48_m7;
 wire booth_b48_m8;
 wire booth_b48_m9;
 wire booth_b4_m0;
 wire booth_b4_m1;
 wire booth_b4_m10;
 wire booth_b4_m11;
 wire booth_b4_m12;
 wire booth_b4_m13;
 wire booth_b4_m14;
 wire booth_b4_m15;
 wire booth_b4_m16;
 wire booth_b4_m17;
 wire booth_b4_m18;
 wire booth_b4_m19;
 wire booth_b4_m2;
 wire booth_b4_m20;
 wire booth_b4_m21;
 wire booth_b4_m22;
 wire booth_b4_m23;
 wire booth_b4_m24;
 wire booth_b4_m25;
 wire booth_b4_m26;
 wire booth_b4_m27;
 wire booth_b4_m28;
 wire booth_b4_m29;
 wire booth_b4_m3;
 wire booth_b4_m30;
 wire booth_b4_m31;
 wire booth_b4_m32;
 wire booth_b4_m33;
 wire booth_b4_m34;
 wire booth_b4_m35;
 wire booth_b4_m36;
 wire booth_b4_m37;
 wire booth_b4_m38;
 wire booth_b4_m39;
 wire booth_b4_m4;
 wire booth_b4_m40;
 wire booth_b4_m41;
 wire booth_b4_m42;
 wire booth_b4_m43;
 wire booth_b4_m44;
 wire booth_b4_m45;
 wire booth_b4_m46;
 wire booth_b4_m47;
 wire booth_b4_m48;
 wire booth_b4_m49;
 wire booth_b4_m5;
 wire booth_b4_m50;
 wire booth_b4_m51;
 wire booth_b4_m52;
 wire booth_b4_m53;
 wire booth_b4_m54;
 wire booth_b4_m55;
 wire booth_b4_m56;
 wire booth_b4_m57;
 wire booth_b4_m58;
 wire booth_b4_m59;
 wire booth_b4_m6;
 wire booth_b4_m60;
 wire booth_b4_m61;
 wire booth_b4_m62;
 wire booth_b4_m63;
 wire booth_b4_m64;
 wire booth_b4_m7;
 wire booth_b4_m8;
 wire booth_b4_m9;
 wire booth_b50_m0;
 wire booth_b50_m1;
 wire booth_b50_m10;
 wire booth_b50_m11;
 wire booth_b50_m12;
 wire booth_b50_m13;
 wire booth_b50_m14;
 wire booth_b50_m15;
 wire booth_b50_m16;
 wire booth_b50_m17;
 wire booth_b50_m18;
 wire booth_b50_m19;
 wire booth_b50_m2;
 wire booth_b50_m20;
 wire booth_b50_m21;
 wire booth_b50_m22;
 wire booth_b50_m23;
 wire booth_b50_m24;
 wire booth_b50_m25;
 wire booth_b50_m26;
 wire booth_b50_m27;
 wire booth_b50_m28;
 wire booth_b50_m29;
 wire booth_b50_m3;
 wire booth_b50_m30;
 wire booth_b50_m31;
 wire booth_b50_m32;
 wire booth_b50_m33;
 wire booth_b50_m34;
 wire booth_b50_m35;
 wire booth_b50_m36;
 wire booth_b50_m37;
 wire booth_b50_m38;
 wire booth_b50_m39;
 wire booth_b50_m4;
 wire booth_b50_m40;
 wire booth_b50_m41;
 wire booth_b50_m42;
 wire booth_b50_m43;
 wire booth_b50_m44;
 wire booth_b50_m45;
 wire booth_b50_m46;
 wire booth_b50_m47;
 wire booth_b50_m48;
 wire booth_b50_m49;
 wire booth_b50_m5;
 wire booth_b50_m50;
 wire booth_b50_m51;
 wire booth_b50_m52;
 wire booth_b50_m53;
 wire booth_b50_m54;
 wire booth_b50_m55;
 wire booth_b50_m56;
 wire booth_b50_m57;
 wire booth_b50_m58;
 wire booth_b50_m59;
 wire booth_b50_m6;
 wire booth_b50_m60;
 wire booth_b50_m61;
 wire booth_b50_m62;
 wire booth_b50_m63;
 wire booth_b50_m64;
 wire booth_b50_m7;
 wire booth_b50_m8;
 wire booth_b50_m9;
 wire booth_b52_m0;
 wire booth_b52_m1;
 wire booth_b52_m10;
 wire booth_b52_m11;
 wire booth_b52_m12;
 wire booth_b52_m13;
 wire booth_b52_m14;
 wire booth_b52_m15;
 wire booth_b52_m16;
 wire booth_b52_m17;
 wire booth_b52_m18;
 wire booth_b52_m19;
 wire booth_b52_m2;
 wire booth_b52_m20;
 wire booth_b52_m21;
 wire booth_b52_m22;
 wire booth_b52_m23;
 wire booth_b52_m24;
 wire booth_b52_m25;
 wire booth_b52_m26;
 wire booth_b52_m27;
 wire booth_b52_m28;
 wire booth_b52_m29;
 wire booth_b52_m3;
 wire booth_b52_m30;
 wire booth_b52_m31;
 wire booth_b52_m32;
 wire booth_b52_m33;
 wire booth_b52_m34;
 wire booth_b52_m35;
 wire booth_b52_m36;
 wire booth_b52_m37;
 wire booth_b52_m38;
 wire booth_b52_m39;
 wire booth_b52_m4;
 wire booth_b52_m40;
 wire booth_b52_m41;
 wire booth_b52_m42;
 wire booth_b52_m43;
 wire booth_b52_m44;
 wire booth_b52_m45;
 wire booth_b52_m46;
 wire booth_b52_m47;
 wire booth_b52_m48;
 wire booth_b52_m49;
 wire booth_b52_m5;
 wire booth_b52_m50;
 wire booth_b52_m51;
 wire booth_b52_m52;
 wire booth_b52_m53;
 wire booth_b52_m54;
 wire booth_b52_m55;
 wire booth_b52_m56;
 wire booth_b52_m57;
 wire booth_b52_m58;
 wire booth_b52_m59;
 wire booth_b52_m6;
 wire booth_b52_m60;
 wire booth_b52_m61;
 wire booth_b52_m62;
 wire booth_b52_m63;
 wire booth_b52_m64;
 wire booth_b52_m7;
 wire booth_b52_m8;
 wire booth_b52_m9;
 wire booth_b54_m0;
 wire booth_b54_m1;
 wire booth_b54_m10;
 wire booth_b54_m11;
 wire booth_b54_m12;
 wire booth_b54_m13;
 wire booth_b54_m14;
 wire booth_b54_m15;
 wire booth_b54_m16;
 wire booth_b54_m17;
 wire booth_b54_m18;
 wire booth_b54_m19;
 wire booth_b54_m2;
 wire booth_b54_m20;
 wire booth_b54_m21;
 wire booth_b54_m22;
 wire booth_b54_m23;
 wire booth_b54_m24;
 wire booth_b54_m25;
 wire booth_b54_m26;
 wire booth_b54_m27;
 wire booth_b54_m28;
 wire booth_b54_m29;
 wire booth_b54_m3;
 wire booth_b54_m30;
 wire booth_b54_m31;
 wire booth_b54_m32;
 wire booth_b54_m33;
 wire booth_b54_m34;
 wire booth_b54_m35;
 wire booth_b54_m36;
 wire booth_b54_m37;
 wire booth_b54_m38;
 wire booth_b54_m39;
 wire booth_b54_m4;
 wire booth_b54_m40;
 wire booth_b54_m41;
 wire booth_b54_m42;
 wire booth_b54_m43;
 wire booth_b54_m44;
 wire booth_b54_m45;
 wire booth_b54_m46;
 wire booth_b54_m47;
 wire booth_b54_m48;
 wire booth_b54_m49;
 wire booth_b54_m5;
 wire booth_b54_m50;
 wire booth_b54_m51;
 wire booth_b54_m52;
 wire booth_b54_m53;
 wire booth_b54_m54;
 wire booth_b54_m55;
 wire booth_b54_m56;
 wire booth_b54_m57;
 wire booth_b54_m58;
 wire booth_b54_m59;
 wire booth_b54_m6;
 wire booth_b54_m60;
 wire booth_b54_m61;
 wire booth_b54_m62;
 wire booth_b54_m63;
 wire booth_b54_m64;
 wire booth_b54_m7;
 wire booth_b54_m8;
 wire booth_b54_m9;
 wire booth_b56_m0;
 wire booth_b56_m1;
 wire booth_b56_m10;
 wire booth_b56_m11;
 wire booth_b56_m12;
 wire booth_b56_m13;
 wire booth_b56_m14;
 wire booth_b56_m15;
 wire booth_b56_m16;
 wire booth_b56_m17;
 wire booth_b56_m18;
 wire booth_b56_m19;
 wire booth_b56_m2;
 wire booth_b56_m20;
 wire booth_b56_m21;
 wire booth_b56_m22;
 wire booth_b56_m23;
 wire booth_b56_m24;
 wire booth_b56_m25;
 wire booth_b56_m26;
 wire booth_b56_m27;
 wire booth_b56_m28;
 wire booth_b56_m29;
 wire booth_b56_m3;
 wire booth_b56_m30;
 wire booth_b56_m31;
 wire booth_b56_m32;
 wire booth_b56_m33;
 wire booth_b56_m34;
 wire booth_b56_m35;
 wire booth_b56_m36;
 wire booth_b56_m37;
 wire booth_b56_m38;
 wire booth_b56_m39;
 wire booth_b56_m4;
 wire booth_b56_m40;
 wire booth_b56_m41;
 wire booth_b56_m42;
 wire booth_b56_m43;
 wire booth_b56_m44;
 wire booth_b56_m45;
 wire booth_b56_m46;
 wire booth_b56_m47;
 wire booth_b56_m48;
 wire booth_b56_m49;
 wire booth_b56_m5;
 wire booth_b56_m50;
 wire booth_b56_m51;
 wire booth_b56_m52;
 wire booth_b56_m53;
 wire booth_b56_m54;
 wire booth_b56_m55;
 wire booth_b56_m56;
 wire booth_b56_m57;
 wire booth_b56_m58;
 wire booth_b56_m59;
 wire booth_b56_m6;
 wire booth_b56_m60;
 wire booth_b56_m61;
 wire booth_b56_m62;
 wire booth_b56_m63;
 wire booth_b56_m64;
 wire booth_b56_m7;
 wire booth_b56_m8;
 wire booth_b56_m9;
 wire booth_b58_m0;
 wire booth_b58_m1;
 wire booth_b58_m10;
 wire booth_b58_m11;
 wire booth_b58_m12;
 wire booth_b58_m13;
 wire booth_b58_m14;
 wire booth_b58_m15;
 wire booth_b58_m16;
 wire booth_b58_m17;
 wire booth_b58_m18;
 wire booth_b58_m19;
 wire booth_b58_m2;
 wire booth_b58_m20;
 wire booth_b58_m21;
 wire booth_b58_m22;
 wire booth_b58_m23;
 wire booth_b58_m24;
 wire booth_b58_m25;
 wire booth_b58_m26;
 wire booth_b58_m27;
 wire booth_b58_m28;
 wire booth_b58_m29;
 wire booth_b58_m3;
 wire booth_b58_m30;
 wire booth_b58_m31;
 wire booth_b58_m32;
 wire booth_b58_m33;
 wire booth_b58_m34;
 wire booth_b58_m35;
 wire booth_b58_m36;
 wire booth_b58_m37;
 wire booth_b58_m38;
 wire booth_b58_m39;
 wire booth_b58_m4;
 wire booth_b58_m40;
 wire booth_b58_m41;
 wire booth_b58_m42;
 wire booth_b58_m43;
 wire booth_b58_m44;
 wire booth_b58_m45;
 wire booth_b58_m46;
 wire booth_b58_m47;
 wire booth_b58_m48;
 wire booth_b58_m49;
 wire booth_b58_m5;
 wire booth_b58_m50;
 wire booth_b58_m51;
 wire booth_b58_m52;
 wire booth_b58_m53;
 wire booth_b58_m54;
 wire booth_b58_m55;
 wire booth_b58_m56;
 wire booth_b58_m57;
 wire booth_b58_m58;
 wire booth_b58_m59;
 wire booth_b58_m6;
 wire booth_b58_m60;
 wire booth_b58_m61;
 wire booth_b58_m62;
 wire booth_b58_m63;
 wire booth_b58_m64;
 wire booth_b58_m7;
 wire booth_b58_m8;
 wire booth_b58_m9;
 wire booth_b60_m0;
 wire booth_b60_m1;
 wire booth_b60_m10;
 wire booth_b60_m11;
 wire booth_b60_m12;
 wire booth_b60_m13;
 wire booth_b60_m14;
 wire booth_b60_m15;
 wire booth_b60_m16;
 wire booth_b60_m17;
 wire booth_b60_m18;
 wire booth_b60_m19;
 wire booth_b60_m2;
 wire booth_b60_m20;
 wire booth_b60_m21;
 wire booth_b60_m22;
 wire booth_b60_m23;
 wire booth_b60_m24;
 wire booth_b60_m25;
 wire booth_b60_m26;
 wire booth_b60_m27;
 wire booth_b60_m28;
 wire booth_b60_m29;
 wire booth_b60_m3;
 wire booth_b60_m30;
 wire booth_b60_m31;
 wire booth_b60_m32;
 wire booth_b60_m33;
 wire booth_b60_m34;
 wire booth_b60_m35;
 wire booth_b60_m36;
 wire booth_b60_m37;
 wire booth_b60_m38;
 wire booth_b60_m39;
 wire booth_b60_m4;
 wire booth_b60_m40;
 wire booth_b60_m41;
 wire booth_b60_m42;
 wire booth_b60_m43;
 wire booth_b60_m44;
 wire booth_b60_m45;
 wire booth_b60_m46;
 wire booth_b60_m47;
 wire booth_b60_m48;
 wire booth_b60_m49;
 wire booth_b60_m5;
 wire booth_b60_m50;
 wire booth_b60_m51;
 wire booth_b60_m52;
 wire booth_b60_m53;
 wire booth_b60_m54;
 wire booth_b60_m55;
 wire booth_b60_m56;
 wire booth_b60_m57;
 wire booth_b60_m58;
 wire booth_b60_m59;
 wire booth_b60_m6;
 wire booth_b60_m60;
 wire booth_b60_m61;
 wire booth_b60_m62;
 wire booth_b60_m63;
 wire booth_b60_m64;
 wire booth_b60_m7;
 wire booth_b60_m8;
 wire booth_b60_m9;
 wire booth_b62_m0;
 wire booth_b62_m1;
 wire booth_b62_m10;
 wire booth_b62_m11;
 wire booth_b62_m12;
 wire booth_b62_m13;
 wire booth_b62_m14;
 wire booth_b62_m15;
 wire booth_b62_m16;
 wire booth_b62_m17;
 wire booth_b62_m18;
 wire booth_b62_m19;
 wire booth_b62_m2;
 wire booth_b62_m20;
 wire booth_b62_m21;
 wire booth_b62_m22;
 wire booth_b62_m23;
 wire booth_b62_m24;
 wire booth_b62_m25;
 wire booth_b62_m26;
 wire booth_b62_m27;
 wire booth_b62_m28;
 wire booth_b62_m29;
 wire booth_b62_m3;
 wire booth_b62_m30;
 wire booth_b62_m31;
 wire booth_b62_m32;
 wire booth_b62_m33;
 wire booth_b62_m34;
 wire booth_b62_m35;
 wire booth_b62_m36;
 wire booth_b62_m37;
 wire booth_b62_m38;
 wire booth_b62_m39;
 wire booth_b62_m4;
 wire booth_b62_m40;
 wire booth_b62_m41;
 wire booth_b62_m42;
 wire booth_b62_m43;
 wire booth_b62_m44;
 wire booth_b62_m45;
 wire booth_b62_m46;
 wire booth_b62_m47;
 wire booth_b62_m48;
 wire booth_b62_m49;
 wire booth_b62_m5;
 wire booth_b62_m50;
 wire booth_b62_m51;
 wire booth_b62_m52;
 wire booth_b62_m53;
 wire booth_b62_m54;
 wire booth_b62_m55;
 wire booth_b62_m56;
 wire booth_b62_m57;
 wire booth_b62_m58;
 wire booth_b62_m59;
 wire booth_b62_m6;
 wire booth_b62_m60;
 wire booth_b62_m61;
 wire booth_b62_m62;
 wire booth_b62_m63;
 wire booth_b62_m64;
 wire booth_b62_m7;
 wire booth_b62_m8;
 wire booth_b62_m9;
 wire booth_b64_m0;
 wire booth_b64_m1;
 wire booth_b64_m10;
 wire booth_b64_m11;
 wire booth_b64_m12;
 wire booth_b64_m13;
 wire booth_b64_m14;
 wire booth_b64_m15;
 wire booth_b64_m16;
 wire booth_b64_m17;
 wire booth_b64_m18;
 wire booth_b64_m19;
 wire booth_b64_m2;
 wire booth_b64_m20;
 wire booth_b64_m21;
 wire booth_b64_m22;
 wire booth_b64_m23;
 wire booth_b64_m24;
 wire booth_b64_m25;
 wire booth_b64_m26;
 wire booth_b64_m27;
 wire booth_b64_m28;
 wire booth_b64_m29;
 wire booth_b64_m3;
 wire booth_b64_m30;
 wire booth_b64_m31;
 wire booth_b64_m32;
 wire booth_b64_m33;
 wire booth_b64_m34;
 wire booth_b64_m35;
 wire booth_b64_m36;
 wire booth_b64_m37;
 wire booth_b64_m38;
 wire booth_b64_m39;
 wire booth_b64_m4;
 wire booth_b64_m40;
 wire booth_b64_m41;
 wire booth_b64_m42;
 wire booth_b64_m43;
 wire booth_b64_m44;
 wire booth_b64_m45;
 wire booth_b64_m46;
 wire booth_b64_m47;
 wire booth_b64_m48;
 wire booth_b64_m49;
 wire booth_b64_m5;
 wire booth_b64_m50;
 wire booth_b64_m51;
 wire booth_b64_m52;
 wire booth_b64_m53;
 wire booth_b64_m54;
 wire booth_b64_m55;
 wire booth_b64_m56;
 wire booth_b64_m57;
 wire booth_b64_m58;
 wire booth_b64_m59;
 wire booth_b64_m6;
 wire booth_b64_m60;
 wire booth_b64_m61;
 wire booth_b64_m62;
 wire booth_b64_m63;
 wire booth_b64_m7;
 wire booth_b64_m8;
 wire booth_b64_m9;
 wire booth_b6_m0;
 wire booth_b6_m1;
 wire booth_b6_m10;
 wire booth_b6_m11;
 wire booth_b6_m12;
 wire booth_b6_m13;
 wire booth_b6_m14;
 wire booth_b6_m15;
 wire booth_b6_m16;
 wire booth_b6_m17;
 wire booth_b6_m18;
 wire booth_b6_m19;
 wire booth_b6_m2;
 wire booth_b6_m20;
 wire booth_b6_m21;
 wire booth_b6_m22;
 wire booth_b6_m23;
 wire booth_b6_m24;
 wire booth_b6_m25;
 wire booth_b6_m26;
 wire booth_b6_m27;
 wire booth_b6_m28;
 wire booth_b6_m29;
 wire booth_b6_m3;
 wire booth_b6_m30;
 wire booth_b6_m31;
 wire booth_b6_m32;
 wire booth_b6_m33;
 wire booth_b6_m34;
 wire booth_b6_m35;
 wire booth_b6_m36;
 wire booth_b6_m37;
 wire booth_b6_m38;
 wire booth_b6_m39;
 wire booth_b6_m4;
 wire booth_b6_m40;
 wire booth_b6_m41;
 wire booth_b6_m42;
 wire booth_b6_m43;
 wire booth_b6_m44;
 wire booth_b6_m45;
 wire booth_b6_m46;
 wire booth_b6_m47;
 wire booth_b6_m48;
 wire booth_b6_m49;
 wire booth_b6_m5;
 wire booth_b6_m50;
 wire booth_b6_m51;
 wire booth_b6_m52;
 wire booth_b6_m53;
 wire booth_b6_m54;
 wire booth_b6_m55;
 wire booth_b6_m56;
 wire booth_b6_m57;
 wire booth_b6_m58;
 wire booth_b6_m59;
 wire booth_b6_m6;
 wire booth_b6_m60;
 wire booth_b6_m61;
 wire booth_b6_m62;
 wire booth_b6_m63;
 wire booth_b6_m64;
 wire booth_b6_m7;
 wire booth_b6_m8;
 wire booth_b6_m9;
 wire booth_b8_m0;
 wire booth_b8_m1;
 wire booth_b8_m10;
 wire booth_b8_m11;
 wire booth_b8_m12;
 wire booth_b8_m13;
 wire booth_b8_m14;
 wire booth_b8_m15;
 wire booth_b8_m16;
 wire booth_b8_m17;
 wire booth_b8_m18;
 wire booth_b8_m19;
 wire booth_b8_m2;
 wire booth_b8_m20;
 wire booth_b8_m21;
 wire booth_b8_m22;
 wire booth_b8_m23;
 wire booth_b8_m24;
 wire booth_b8_m25;
 wire booth_b8_m26;
 wire booth_b8_m27;
 wire booth_b8_m28;
 wire booth_b8_m29;
 wire booth_b8_m3;
 wire booth_b8_m30;
 wire booth_b8_m31;
 wire booth_b8_m32;
 wire booth_b8_m33;
 wire booth_b8_m34;
 wire booth_b8_m35;
 wire booth_b8_m36;
 wire booth_b8_m37;
 wire booth_b8_m38;
 wire booth_b8_m39;
 wire booth_b8_m4;
 wire booth_b8_m40;
 wire booth_b8_m41;
 wire booth_b8_m42;
 wire booth_b8_m43;
 wire booth_b8_m44;
 wire booth_b8_m45;
 wire booth_b8_m46;
 wire booth_b8_m47;
 wire booth_b8_m48;
 wire booth_b8_m49;
 wire booth_b8_m5;
 wire booth_b8_m50;
 wire booth_b8_m51;
 wire booth_b8_m52;
 wire booth_b8_m53;
 wire booth_b8_m54;
 wire booth_b8_m55;
 wire booth_b8_m56;
 wire booth_b8_m57;
 wire booth_b8_m58;
 wire booth_b8_m59;
 wire booth_b8_m6;
 wire booth_b8_m60;
 wire booth_b8_m61;
 wire booth_b8_m62;
 wire booth_b8_m63;
 wire booth_b8_m64;
 wire booth_b8_m7;
 wire booth_b8_m8;
 wire booth_b8_m9;
 wire \c$1 ;
 wire \c$10 ;
 wire \c$100 ;
 wire \c$1000 ;
 wire \c$1002 ;
 wire \c$1004 ;
 wire \c$1006 ;
 wire \c$1008 ;
 wire \c$1010 ;
 wire \c$1012 ;
 wire \c$1014 ;
 wire \c$1016 ;
 wire \c$1018 ;
 wire \c$102 ;
 wire \c$1020 ;
 wire \c$1022 ;
 wire \c$1024 ;
 wire \c$1026 ;
 wire \c$1028 ;
 wire \c$1030 ;
 wire \c$1032 ;
 wire \c$1034 ;
 wire \c$1036 ;
 wire \c$1038 ;
 wire \c$104 ;
 wire \c$1040 ;
 wire \c$1042 ;
 wire \c$1044 ;
 wire \c$1046 ;
 wire \c$1048 ;
 wire \c$1050 ;
 wire \c$1052 ;
 wire \c$1054 ;
 wire \c$1056 ;
 wire \c$1058 ;
 wire \c$106 ;
 wire \c$1060 ;
 wire \c$1062 ;
 wire \c$1064 ;
 wire \c$1066 ;
 wire \c$1068 ;
 wire \c$1070 ;
 wire \c$1072 ;
 wire \c$1074 ;
 wire \c$1076 ;
 wire \c$1078 ;
 wire \c$108 ;
 wire \c$1080 ;
 wire \c$1082 ;
 wire \c$1084 ;
 wire \c$1086 ;
 wire \c$1088 ;
 wire \c$1090 ;
 wire \c$1092 ;
 wire \c$1094 ;
 wire \c$1096 ;
 wire \c$1098 ;
 wire \c$110 ;
 wire \c$1100 ;
 wire \c$1102 ;
 wire \c$1104 ;
 wire \c$1106 ;
 wire \c$1108 ;
 wire \c$1110 ;
 wire \c$1112 ;
 wire \c$1114 ;
 wire \c$1116 ;
 wire \c$1118 ;
 wire \c$112 ;
 wire \c$1120 ;
 wire \c$1122 ;
 wire \c$1124 ;
 wire \c$1126 ;
 wire \c$1128 ;
 wire \c$1130 ;
 wire \c$1132 ;
 wire \c$1134 ;
 wire \c$1136 ;
 wire \c$1138 ;
 wire \c$114 ;
 wire \c$1140 ;
 wire \c$1142 ;
 wire \c$1144 ;
 wire \c$1146 ;
 wire \c$1148 ;
 wire \c$1150 ;
 wire \c$1152 ;
 wire \c$1154 ;
 wire \c$1156 ;
 wire \c$1158 ;
 wire \c$116 ;
 wire \c$1160 ;
 wire \c$1162 ;
 wire \c$1164 ;
 wire \c$1166 ;
 wire \c$1168 ;
 wire \c$1170 ;
 wire \c$1172 ;
 wire \c$1174 ;
 wire \c$1176 ;
 wire \c$1178 ;
 wire \c$118 ;
 wire \c$1180 ;
 wire \c$1182 ;
 wire \c$1184 ;
 wire \c$1186 ;
 wire \c$1188 ;
 wire \c$1190 ;
 wire \c$1192 ;
 wire \c$1194 ;
 wire \c$1196 ;
 wire \c$1198 ;
 wire \c$12 ;
 wire \c$120 ;
 wire \c$1200 ;
 wire \c$1202 ;
 wire \c$1204 ;
 wire \c$1206 ;
 wire \c$1208 ;
 wire \c$1210 ;
 wire \c$1212 ;
 wire \c$1214 ;
 wire \c$1216 ;
 wire \c$1218 ;
 wire \c$122 ;
 wire \c$1220 ;
 wire \c$1222 ;
 wire \c$1224 ;
 wire \c$1226 ;
 wire \c$1228 ;
 wire \c$1230 ;
 wire \c$1232 ;
 wire \c$1234 ;
 wire \c$1236 ;
 wire \c$1238 ;
 wire \c$124 ;
 wire \c$1240 ;
 wire \c$1242 ;
 wire \c$1244 ;
 wire \c$1246 ;
 wire \c$1248 ;
 wire \c$1250 ;
 wire \c$1252 ;
 wire \c$1254 ;
 wire \c$1256 ;
 wire \c$1258 ;
 wire \c$126 ;
 wire \c$1260 ;
 wire \c$1262 ;
 wire \c$1264 ;
 wire \c$1266 ;
 wire \c$1268 ;
 wire \c$1270 ;
 wire \c$1272 ;
 wire \c$1274 ;
 wire \c$1276 ;
 wire \c$1278 ;
 wire \c$128 ;
 wire \c$1280 ;
 wire \c$1282 ;
 wire \c$1284 ;
 wire \c$1286 ;
 wire \c$1288 ;
 wire \c$1290 ;
 wire \c$1292 ;
 wire \c$1294 ;
 wire \c$1296 ;
 wire \c$1298 ;
 wire \c$130 ;
 wire \c$1300 ;
 wire \c$1302 ;
 wire \c$1304 ;
 wire \c$1306 ;
 wire \c$1308 ;
 wire \c$1310 ;
 wire \c$1312 ;
 wire \c$1314 ;
 wire \c$1316 ;
 wire \c$1318 ;
 wire \c$132 ;
 wire \c$1320 ;
 wire \c$1322 ;
 wire \c$1324 ;
 wire \c$1326 ;
 wire \c$1328 ;
 wire \c$1330 ;
 wire \c$1332 ;
 wire \c$1334 ;
 wire \c$1336 ;
 wire \c$1338 ;
 wire \c$134 ;
 wire \c$1340 ;
 wire \c$1342 ;
 wire \c$1344 ;
 wire \c$1346 ;
 wire \c$1348 ;
 wire \c$1350 ;
 wire \c$1352 ;
 wire \c$1354 ;
 wire \c$1356 ;
 wire \c$1358 ;
 wire \c$136 ;
 wire \c$1360 ;
 wire \c$1362 ;
 wire \c$1364 ;
 wire \c$1366 ;
 wire \c$1368 ;
 wire \c$1370 ;
 wire \c$1372 ;
 wire \c$1374 ;
 wire \c$1376 ;
 wire \c$1378 ;
 wire \c$138 ;
 wire \c$1380 ;
 wire \c$1382 ;
 wire \c$1384 ;
 wire \c$1386 ;
 wire \c$1388 ;
 wire \c$1390 ;
 wire \c$1392 ;
 wire \c$1394 ;
 wire \c$1396 ;
 wire \c$1398 ;
 wire \c$14 ;
 wire \c$140 ;
 wire \c$1400 ;
 wire \c$1402 ;
 wire \c$1404 ;
 wire \c$1406 ;
 wire \c$1408 ;
 wire \c$1410 ;
 wire \c$1412 ;
 wire \c$1414 ;
 wire \c$1416 ;
 wire \c$1418 ;
 wire \c$142 ;
 wire \c$1420 ;
 wire \c$1422 ;
 wire \c$1424 ;
 wire \c$1426 ;
 wire \c$1428 ;
 wire \c$1430 ;
 wire \c$1432 ;
 wire \c$1434 ;
 wire \c$1436 ;
 wire \c$1438 ;
 wire \c$144 ;
 wire \c$1440 ;
 wire \c$1442 ;
 wire \c$1444 ;
 wire \c$1446 ;
 wire \c$1448 ;
 wire \c$1450 ;
 wire \c$1452 ;
 wire \c$1454 ;
 wire \c$1456 ;
 wire \c$1458 ;
 wire \c$146 ;
 wire \c$1460 ;
 wire \c$1462 ;
 wire \c$1464 ;
 wire \c$1466 ;
 wire \c$1468 ;
 wire \c$1470 ;
 wire \c$1472 ;
 wire \c$1474 ;
 wire \c$1476 ;
 wire \c$1478 ;
 wire \c$148 ;
 wire \c$1480 ;
 wire \c$1482 ;
 wire \c$1484 ;
 wire \c$1486 ;
 wire \c$1488 ;
 wire \c$1490 ;
 wire \c$1492 ;
 wire \c$1494 ;
 wire \c$1496 ;
 wire \c$1498 ;
 wire \c$150 ;
 wire \c$1500 ;
 wire \c$1502 ;
 wire \c$1504 ;
 wire \c$1506 ;
 wire \c$1508 ;
 wire \c$1510 ;
 wire \c$1512 ;
 wire \c$1514 ;
 wire \c$1516 ;
 wire \c$1518 ;
 wire \c$152 ;
 wire \c$1520 ;
 wire \c$1522 ;
 wire \c$1524 ;
 wire \c$1526 ;
 wire \c$1528 ;
 wire \c$1530 ;
 wire \c$1532 ;
 wire \c$1534 ;
 wire \c$1536 ;
 wire \c$1538 ;
 wire \c$154 ;
 wire \c$1540 ;
 wire \c$1542 ;
 wire \c$1544 ;
 wire \c$1546 ;
 wire \c$1548 ;
 wire \c$1550 ;
 wire \c$1552 ;
 wire \c$1554 ;
 wire \c$1556 ;
 wire \c$1558 ;
 wire \c$156 ;
 wire \c$1560 ;
 wire \c$1562 ;
 wire \c$1564 ;
 wire \c$1566 ;
 wire \c$1568 ;
 wire \c$1570 ;
 wire \c$1572 ;
 wire \c$1574 ;
 wire \c$1576 ;
 wire \c$1578 ;
 wire \c$158 ;
 wire \c$1580 ;
 wire \c$1582 ;
 wire \c$1584 ;
 wire \c$1586 ;
 wire \c$1588 ;
 wire \c$1590 ;
 wire \c$1592 ;
 wire \c$1594 ;
 wire \c$1596 ;
 wire \c$1598 ;
 wire \c$16 ;
 wire \c$160 ;
 wire \c$1600 ;
 wire \c$1602 ;
 wire \c$1604 ;
 wire \c$1606 ;
 wire \c$1608 ;
 wire \c$1610 ;
 wire \c$1612 ;
 wire \c$1614 ;
 wire \c$1616 ;
 wire \c$1618 ;
 wire \c$162 ;
 wire \c$1620 ;
 wire \c$1622 ;
 wire \c$1624 ;
 wire \c$1626 ;
 wire \c$1628 ;
 wire \c$1630 ;
 wire \c$1632 ;
 wire \c$1634 ;
 wire \c$1636 ;
 wire \c$1638 ;
 wire \c$164 ;
 wire \c$1640 ;
 wire \c$1642 ;
 wire \c$1644 ;
 wire \c$1646 ;
 wire \c$1648 ;
 wire \c$1650 ;
 wire \c$1652 ;
 wire \c$1654 ;
 wire \c$1656 ;
 wire \c$1658 ;
 wire \c$166 ;
 wire \c$1660 ;
 wire \c$1662 ;
 wire \c$1664 ;
 wire \c$1666 ;
 wire \c$1668 ;
 wire \c$1670 ;
 wire \c$1672 ;
 wire \c$1674 ;
 wire \c$1676 ;
 wire \c$1678 ;
 wire \c$168 ;
 wire \c$1680 ;
 wire \c$1682 ;
 wire \c$1684 ;
 wire \c$1686 ;
 wire \c$1688 ;
 wire \c$1690 ;
 wire \c$1692 ;
 wire \c$1694 ;
 wire \c$1696 ;
 wire \c$1698 ;
 wire \c$170 ;
 wire \c$1700 ;
 wire \c$1702 ;
 wire \c$1704 ;
 wire \c$1706 ;
 wire \c$1708 ;
 wire \c$1710 ;
 wire \c$1712 ;
 wire \c$1714 ;
 wire \c$1716 ;
 wire \c$1718 ;
 wire \c$172 ;
 wire \c$1720 ;
 wire \c$1722 ;
 wire \c$1724 ;
 wire \c$1726 ;
 wire \c$1728 ;
 wire \c$1730 ;
 wire \c$1732 ;
 wire \c$1734 ;
 wire \c$1736 ;
 wire \c$1738 ;
 wire \c$174 ;
 wire \c$1740 ;
 wire \c$1742 ;
 wire \c$1744 ;
 wire \c$1746 ;
 wire \c$1748 ;
 wire \c$1750 ;
 wire \c$1752 ;
 wire \c$1754 ;
 wire \c$1756 ;
 wire \c$1758 ;
 wire \c$176 ;
 wire \c$1760 ;
 wire \c$1762 ;
 wire \c$1764 ;
 wire \c$1766 ;
 wire \c$1768 ;
 wire \c$1770 ;
 wire \c$1772 ;
 wire \c$1774 ;
 wire \c$1776 ;
 wire \c$1778 ;
 wire \c$178 ;
 wire \c$1780 ;
 wire \c$1782 ;
 wire \c$1784 ;
 wire \c$1786 ;
 wire \c$1788 ;
 wire \c$1790 ;
 wire \c$1792 ;
 wire \c$1794 ;
 wire \c$1796 ;
 wire \c$1798 ;
 wire \c$18 ;
 wire \c$180 ;
 wire \c$1800 ;
 wire \c$1802 ;
 wire \c$1804 ;
 wire \c$1806 ;
 wire \c$1808 ;
 wire \c$1810 ;
 wire \c$1812 ;
 wire \c$1814 ;
 wire \c$1816 ;
 wire \c$1818 ;
 wire \c$182 ;
 wire \c$1820 ;
 wire \c$1822 ;
 wire \c$1824 ;
 wire \c$1826 ;
 wire \c$1828 ;
 wire \c$1830 ;
 wire \c$1832 ;
 wire \c$1834 ;
 wire \c$1836 ;
 wire \c$1838 ;
 wire \c$184 ;
 wire \c$1840 ;
 wire \c$1842 ;
 wire \c$1844 ;
 wire \c$1846 ;
 wire \c$1848 ;
 wire \c$1850 ;
 wire \c$1852 ;
 wire \c$1854 ;
 wire \c$1856 ;
 wire \c$1858 ;
 wire \c$186 ;
 wire \c$1860 ;
 wire \c$1862 ;
 wire \c$1864 ;
 wire \c$1866 ;
 wire \c$1868 ;
 wire \c$1870 ;
 wire \c$1872 ;
 wire \c$1874 ;
 wire \c$1876 ;
 wire \c$1878 ;
 wire \c$188 ;
 wire \c$1880 ;
 wire \c$1882 ;
 wire \c$1884 ;
 wire \c$1886 ;
 wire \c$1888 ;
 wire \c$1890 ;
 wire \c$1892 ;
 wire \c$1894 ;
 wire \c$1896 ;
 wire \c$1898 ;
 wire \c$190 ;
 wire \c$1900 ;
 wire \c$1902 ;
 wire \c$1904 ;
 wire \c$1906 ;
 wire \c$1908 ;
 wire \c$1910 ;
 wire \c$1912 ;
 wire \c$1914 ;
 wire \c$1916 ;
 wire \c$1918 ;
 wire \c$192 ;
 wire \c$1920 ;
 wire \c$1922 ;
 wire \c$1924 ;
 wire \c$1926 ;
 wire \c$1928 ;
 wire \c$1930 ;
 wire \c$1932 ;
 wire \c$1934 ;
 wire \c$1936 ;
 wire \c$1938 ;
 wire \c$194 ;
 wire \c$1940 ;
 wire \c$1942 ;
 wire \c$1944 ;
 wire \c$1946 ;
 wire \c$1948 ;
 wire \c$1950 ;
 wire \c$1952 ;
 wire \c$1954 ;
 wire \c$1956 ;
 wire \c$1958 ;
 wire \c$196 ;
 wire \c$1960 ;
 wire \c$1962 ;
 wire \c$1964 ;
 wire \c$1966 ;
 wire \c$1968 ;
 wire \c$1970 ;
 wire \c$1972 ;
 wire \c$1974 ;
 wire \c$1976 ;
 wire \c$1978 ;
 wire \c$198 ;
 wire \c$1980 ;
 wire \c$1982 ;
 wire \c$1984 ;
 wire \c$1986 ;
 wire \c$1988 ;
 wire \c$1990 ;
 wire \c$1992 ;
 wire \c$1994 ;
 wire \c$1996 ;
 wire \c$1998 ;
 wire \c$2 ;
 wire \c$20 ;
 wire \c$200 ;
 wire \c$2000 ;
 wire \c$2002 ;
 wire \c$2004 ;
 wire \c$2006 ;
 wire \c$2008 ;
 wire \c$2010 ;
 wire \c$2012 ;
 wire \c$2014 ;
 wire \c$2016 ;
 wire \c$2018 ;
 wire \c$202 ;
 wire \c$2020 ;
 wire \c$2022 ;
 wire \c$2024 ;
 wire \c$2026 ;
 wire \c$2028 ;
 wire \c$2030 ;
 wire \c$2032 ;
 wire \c$2034 ;
 wire \c$2036 ;
 wire \c$2038 ;
 wire \c$204 ;
 wire \c$2040 ;
 wire \c$2042 ;
 wire \c$2044 ;
 wire \c$2046 ;
 wire \c$2048 ;
 wire \c$2050 ;
 wire \c$2052 ;
 wire \c$2054 ;
 wire \c$2056 ;
 wire \c$2058 ;
 wire \c$206 ;
 wire \c$2060 ;
 wire \c$2062 ;
 wire \c$2064 ;
 wire \c$2066 ;
 wire \c$2068 ;
 wire \c$2070 ;
 wire \c$2072 ;
 wire \c$2074 ;
 wire \c$2076 ;
 wire \c$2078 ;
 wire \c$208 ;
 wire \c$2080 ;
 wire \c$2082 ;
 wire \c$2084 ;
 wire \c$2086 ;
 wire \c$2088 ;
 wire \c$2090 ;
 wire \c$2092 ;
 wire \c$2094 ;
 wire \c$2096 ;
 wire \c$2098 ;
 wire \c$210 ;
 wire \c$2100 ;
 wire \c$2102 ;
 wire \c$2104 ;
 wire \c$2106 ;
 wire \c$2108 ;
 wire \c$2110 ;
 wire \c$2112 ;
 wire \c$2114 ;
 wire \c$2116 ;
 wire \c$2118 ;
 wire \c$212 ;
 wire \c$2120 ;
 wire \c$2122 ;
 wire \c$2124 ;
 wire \c$2126 ;
 wire \c$2128 ;
 wire \c$2130 ;
 wire \c$2132 ;
 wire \c$2134 ;
 wire \c$2136 ;
 wire \c$2138 ;
 wire \c$214 ;
 wire \c$2140 ;
 wire \c$2142 ;
 wire \c$2144 ;
 wire \c$2146 ;
 wire \c$2148 ;
 wire \c$2150 ;
 wire \c$2152 ;
 wire \c$2154 ;
 wire \c$2156 ;
 wire \c$2158 ;
 wire \c$216 ;
 wire \c$2160 ;
 wire \c$2162 ;
 wire \c$2164 ;
 wire \c$2166 ;
 wire \c$2168 ;
 wire \c$2170 ;
 wire \c$2172 ;
 wire \c$2174 ;
 wire \c$2176 ;
 wire \c$2178 ;
 wire \c$218 ;
 wire \c$2180 ;
 wire \c$2182 ;
 wire \c$2184 ;
 wire \c$2186 ;
 wire \c$2188 ;
 wire \c$2190 ;
 wire \c$2192 ;
 wire \c$2194 ;
 wire \c$2196 ;
 wire \c$2198 ;
 wire \c$22 ;
 wire \c$220 ;
 wire \c$2200 ;
 wire \c$2202 ;
 wire \c$2204 ;
 wire \c$2206 ;
 wire \c$2208 ;
 wire \c$2210 ;
 wire \c$2212 ;
 wire \c$2214 ;
 wire \c$2216 ;
 wire \c$2218 ;
 wire \c$222 ;
 wire \c$2220 ;
 wire \c$2222 ;
 wire \c$2224 ;
 wire \c$2226 ;
 wire \c$2228 ;
 wire \c$2230 ;
 wire \c$2232 ;
 wire \c$2234 ;
 wire \c$2236 ;
 wire \c$2238 ;
 wire \c$224 ;
 wire \c$2240 ;
 wire \c$2242 ;
 wire \c$2244 ;
 wire \c$2246 ;
 wire \c$2248 ;
 wire \c$2250 ;
 wire \c$2252 ;
 wire \c$2254 ;
 wire \c$2256 ;
 wire \c$2258 ;
 wire \c$226 ;
 wire \c$2260 ;
 wire \c$2262 ;
 wire \c$2264 ;
 wire \c$2266 ;
 wire \c$2268 ;
 wire \c$2270 ;
 wire \c$2272 ;
 wire \c$2274 ;
 wire \c$2276 ;
 wire \c$2278 ;
 wire \c$228 ;
 wire \c$2280 ;
 wire \c$2282 ;
 wire \c$2284 ;
 wire \c$2286 ;
 wire \c$2288 ;
 wire \c$2290 ;
 wire \c$2292 ;
 wire \c$2294 ;
 wire \c$2296 ;
 wire \c$2298 ;
 wire \c$230 ;
 wire \c$2300 ;
 wire \c$2302 ;
 wire \c$2304 ;
 wire \c$2306 ;
 wire \c$2308 ;
 wire \c$2310 ;
 wire \c$2312 ;
 wire \c$2314 ;
 wire \c$2316 ;
 wire \c$2318 ;
 wire \c$232 ;
 wire \c$2320 ;
 wire \c$2322 ;
 wire \c$2324 ;
 wire \c$2326 ;
 wire \c$2328 ;
 wire \c$2330 ;
 wire \c$2332 ;
 wire \c$2334 ;
 wire \c$2336 ;
 wire \c$2338 ;
 wire \c$234 ;
 wire \c$2340 ;
 wire \c$2342 ;
 wire \c$2344 ;
 wire \c$2346 ;
 wire \c$2348 ;
 wire \c$2350 ;
 wire \c$2352 ;
 wire \c$2354 ;
 wire \c$2356 ;
 wire \c$2358 ;
 wire \c$236 ;
 wire \c$2360 ;
 wire \c$2362 ;
 wire \c$2364 ;
 wire \c$2366 ;
 wire \c$2368 ;
 wire \c$2370 ;
 wire \c$2372 ;
 wire \c$2374 ;
 wire \c$2376 ;
 wire \c$2378 ;
 wire \c$238 ;
 wire \c$2380 ;
 wire \c$2382 ;
 wire \c$2384 ;
 wire \c$2386 ;
 wire \c$2388 ;
 wire \c$2390 ;
 wire \c$2392 ;
 wire \c$2394 ;
 wire \c$2396 ;
 wire \c$2398 ;
 wire \c$24 ;
 wire \c$240 ;
 wire \c$2400 ;
 wire \c$2402 ;
 wire \c$2404 ;
 wire \c$2406 ;
 wire \c$2408 ;
 wire \c$2410 ;
 wire \c$2412 ;
 wire \c$2414 ;
 wire \c$2416 ;
 wire \c$2418 ;
 wire \c$242 ;
 wire \c$2420 ;
 wire \c$2422 ;
 wire \c$2424 ;
 wire \c$2426 ;
 wire \c$2428 ;
 wire \c$2430 ;
 wire \c$2432 ;
 wire \c$2434 ;
 wire \c$2436 ;
 wire \c$2438 ;
 wire \c$244 ;
 wire \c$2440 ;
 wire \c$2442 ;
 wire \c$2444 ;
 wire \c$2446 ;
 wire \c$2448 ;
 wire \c$2450 ;
 wire \c$2452 ;
 wire \c$2454 ;
 wire \c$2456 ;
 wire \c$2458 ;
 wire \c$246 ;
 wire \c$2460 ;
 wire \c$2462 ;
 wire \c$2464 ;
 wire \c$2466 ;
 wire \c$2468 ;
 wire \c$2470 ;
 wire \c$2472 ;
 wire \c$2474 ;
 wire \c$2476 ;
 wire \c$2478 ;
 wire \c$248 ;
 wire \c$2480 ;
 wire \c$2482 ;
 wire \c$2484 ;
 wire \c$2486 ;
 wire \c$2488 ;
 wire \c$2490 ;
 wire \c$2492 ;
 wire \c$2494 ;
 wire \c$2496 ;
 wire \c$2498 ;
 wire \c$250 ;
 wire \c$2500 ;
 wire \c$2502 ;
 wire \c$2504 ;
 wire \c$2506 ;
 wire \c$2508 ;
 wire \c$2510 ;
 wire \c$2512 ;
 wire \c$2514 ;
 wire \c$2516 ;
 wire \c$2518 ;
 wire \c$252 ;
 wire \c$2520 ;
 wire \c$2522 ;
 wire \c$2524 ;
 wire \c$2526 ;
 wire \c$2528 ;
 wire \c$2530 ;
 wire \c$2532 ;
 wire \c$2534 ;
 wire \c$2536 ;
 wire \c$2538 ;
 wire \c$254 ;
 wire \c$2540 ;
 wire \c$2542 ;
 wire \c$2544 ;
 wire \c$2546 ;
 wire \c$2548 ;
 wire \c$2550 ;
 wire \c$2552 ;
 wire \c$2554 ;
 wire \c$2556 ;
 wire \c$2558 ;
 wire \c$256 ;
 wire \c$2560 ;
 wire \c$2562 ;
 wire \c$2564 ;
 wire \c$2566 ;
 wire \c$2568 ;
 wire \c$2570 ;
 wire \c$2572 ;
 wire \c$2574 ;
 wire \c$2576 ;
 wire \c$2578 ;
 wire \c$258 ;
 wire \c$2580 ;
 wire \c$2582 ;
 wire \c$2584 ;
 wire \c$2586 ;
 wire \c$2588 ;
 wire \c$2590 ;
 wire \c$2592 ;
 wire \c$2594 ;
 wire \c$2596 ;
 wire \c$2598 ;
 wire \c$26 ;
 wire \c$260 ;
 wire \c$2600 ;
 wire \c$2602 ;
 wire \c$2604 ;
 wire \c$2606 ;
 wire \c$2608 ;
 wire \c$2610 ;
 wire \c$2612 ;
 wire \c$2614 ;
 wire \c$2616 ;
 wire \c$2618 ;
 wire \c$262 ;
 wire \c$2620 ;
 wire \c$2622 ;
 wire \c$2624 ;
 wire \c$2626 ;
 wire \c$2628 ;
 wire \c$2630 ;
 wire \c$2632 ;
 wire \c$2634 ;
 wire \c$2636 ;
 wire \c$2638 ;
 wire \c$264 ;
 wire \c$2640 ;
 wire \c$2642 ;
 wire \c$2644 ;
 wire \c$2646 ;
 wire \c$2648 ;
 wire \c$2650 ;
 wire \c$2652 ;
 wire \c$2654 ;
 wire \c$2656 ;
 wire \c$2658 ;
 wire \c$266 ;
 wire \c$2660 ;
 wire \c$2662 ;
 wire \c$2664 ;
 wire \c$2666 ;
 wire \c$2668 ;
 wire \c$2670 ;
 wire \c$2672 ;
 wire \c$2674 ;
 wire \c$2676 ;
 wire \c$2678 ;
 wire \c$268 ;
 wire \c$2680 ;
 wire \c$2682 ;
 wire \c$2684 ;
 wire \c$2686 ;
 wire \c$2688 ;
 wire \c$2690 ;
 wire \c$2692 ;
 wire \c$2694 ;
 wire \c$2696 ;
 wire \c$2698 ;
 wire \c$270 ;
 wire \c$2700 ;
 wire \c$2702 ;
 wire \c$2704 ;
 wire \c$2706 ;
 wire \c$2708 ;
 wire \c$2710 ;
 wire \c$2712 ;
 wire \c$2714 ;
 wire \c$2716 ;
 wire \c$2718 ;
 wire \c$272 ;
 wire \c$2720 ;
 wire \c$2722 ;
 wire \c$2724 ;
 wire \c$2726 ;
 wire \c$2728 ;
 wire \c$2730 ;
 wire \c$2732 ;
 wire \c$2734 ;
 wire \c$2736 ;
 wire \c$2738 ;
 wire \c$274 ;
 wire \c$2740 ;
 wire \c$2742 ;
 wire \c$2744 ;
 wire \c$2746 ;
 wire \c$2748 ;
 wire \c$2750 ;
 wire \c$2752 ;
 wire \c$2754 ;
 wire \c$2756 ;
 wire \c$2758 ;
 wire \c$276 ;
 wire \c$2760 ;
 wire \c$2762 ;
 wire \c$2764 ;
 wire \c$2766 ;
 wire \c$2768 ;
 wire \c$2770 ;
 wire \c$2772 ;
 wire \c$2774 ;
 wire \c$2776 ;
 wire \c$2778 ;
 wire \c$278 ;
 wire \c$2780 ;
 wire \c$2782 ;
 wire \c$2784 ;
 wire \c$2786 ;
 wire \c$2788 ;
 wire \c$2790 ;
 wire \c$2792 ;
 wire \c$2794 ;
 wire \c$2796 ;
 wire \c$2798 ;
 wire \c$28 ;
 wire \c$280 ;
 wire \c$2800 ;
 wire \c$2802 ;
 wire \c$2804 ;
 wire \c$2806 ;
 wire \c$2808 ;
 wire \c$2810 ;
 wire \c$2812 ;
 wire \c$2814 ;
 wire \c$2816 ;
 wire \c$2818 ;
 wire \c$282 ;
 wire \c$2820 ;
 wire \c$2822 ;
 wire \c$2824 ;
 wire \c$2826 ;
 wire \c$2828 ;
 wire \c$2830 ;
 wire \c$2832 ;
 wire \c$2834 ;
 wire \c$2836 ;
 wire \c$2838 ;
 wire \c$284 ;
 wire \c$2840 ;
 wire \c$2842 ;
 wire \c$2844 ;
 wire \c$2846 ;
 wire \c$2848 ;
 wire \c$2850 ;
 wire \c$2852 ;
 wire \c$2854 ;
 wire \c$2856 ;
 wire \c$2858 ;
 wire \c$286 ;
 wire \c$2860 ;
 wire \c$2862 ;
 wire \c$2864 ;
 wire \c$2866 ;
 wire \c$2868 ;
 wire \c$2870 ;
 wire \c$2872 ;
 wire \c$2874 ;
 wire \c$2876 ;
 wire \c$2878 ;
 wire \c$288 ;
 wire \c$2880 ;
 wire \c$2882 ;
 wire \c$2884 ;
 wire \c$2886 ;
 wire \c$2888 ;
 wire \c$2890 ;
 wire \c$2892 ;
 wire \c$2894 ;
 wire \c$2896 ;
 wire \c$2898 ;
 wire \c$290 ;
 wire \c$2900 ;
 wire \c$2902 ;
 wire \c$2904 ;
 wire \c$2906 ;
 wire \c$2908 ;
 wire \c$2910 ;
 wire \c$2912 ;
 wire \c$2914 ;
 wire \c$2916 ;
 wire \c$2918 ;
 wire \c$292 ;
 wire \c$2920 ;
 wire \c$2922 ;
 wire \c$2924 ;
 wire \c$2926 ;
 wire \c$2928 ;
 wire \c$2930 ;
 wire \c$2932 ;
 wire \c$2934 ;
 wire \c$2936 ;
 wire \c$2938 ;
 wire \c$294 ;
 wire \c$2940 ;
 wire \c$2942 ;
 wire \c$2944 ;
 wire \c$2946 ;
 wire \c$2948 ;
 wire \c$2950 ;
 wire \c$2952 ;
 wire \c$2954 ;
 wire \c$2956 ;
 wire \c$2958 ;
 wire \c$296 ;
 wire \c$2960 ;
 wire \c$2962 ;
 wire \c$2964 ;
 wire \c$2966 ;
 wire \c$2968 ;
 wire \c$2970 ;
 wire \c$2972 ;
 wire \c$2974 ;
 wire \c$2976 ;
 wire \c$2978 ;
 wire \c$298 ;
 wire \c$2980 ;
 wire \c$2982 ;
 wire \c$2984 ;
 wire \c$2986 ;
 wire \c$2988 ;
 wire \c$2990 ;
 wire \c$2992 ;
 wire \c$2994 ;
 wire \c$2996 ;
 wire \c$2998 ;
 wire \c$30 ;
 wire \c$300 ;
 wire \c$3000 ;
 wire \c$3002 ;
 wire \c$3004 ;
 wire \c$3006 ;
 wire \c$3008 ;
 wire \c$3010 ;
 wire \c$3012 ;
 wire \c$3014 ;
 wire \c$3016 ;
 wire \c$3018 ;
 wire \c$302 ;
 wire \c$3020 ;
 wire \c$3022 ;
 wire \c$3024 ;
 wire \c$3026 ;
 wire \c$3028 ;
 wire \c$3030 ;
 wire \c$3032 ;
 wire \c$3034 ;
 wire \c$3036 ;
 wire \c$3038 ;
 wire \c$304 ;
 wire \c$3040 ;
 wire \c$3042 ;
 wire \c$3044 ;
 wire \c$3046 ;
 wire \c$3048 ;
 wire \c$3050 ;
 wire \c$3052 ;
 wire \c$3054 ;
 wire \c$3056 ;
 wire \c$3058 ;
 wire \c$306 ;
 wire \c$3060 ;
 wire \c$3062 ;
 wire \c$3064 ;
 wire \c$3066 ;
 wire \c$3068 ;
 wire \c$3070 ;
 wire \c$3072 ;
 wire \c$3074 ;
 wire \c$3076 ;
 wire \c$3078 ;
 wire \c$308 ;
 wire \c$3080 ;
 wire \c$3082 ;
 wire \c$3084 ;
 wire \c$3086 ;
 wire \c$3088 ;
 wire \c$3090 ;
 wire \c$3092 ;
 wire \c$3094 ;
 wire \c$3096 ;
 wire \c$3098 ;
 wire \c$310 ;
 wire \c$3100 ;
 wire \c$3102 ;
 wire \c$3104 ;
 wire \c$3106 ;
 wire \c$3108 ;
 wire \c$3110 ;
 wire \c$3112 ;
 wire \c$3114 ;
 wire \c$3116 ;
 wire \c$3118 ;
 wire \c$312 ;
 wire \c$3120 ;
 wire \c$3122 ;
 wire \c$3124 ;
 wire \c$3126 ;
 wire \c$3128 ;
 wire \c$3130 ;
 wire \c$3132 ;
 wire \c$3134 ;
 wire \c$3136 ;
 wire \c$3138 ;
 wire \c$314 ;
 wire \c$3140 ;
 wire \c$3142 ;
 wire \c$3144 ;
 wire \c$3146 ;
 wire \c$3148 ;
 wire \c$3150 ;
 wire \c$3152 ;
 wire \c$3154 ;
 wire \c$3156 ;
 wire \c$3158 ;
 wire \c$316 ;
 wire \c$3160 ;
 wire \c$3162 ;
 wire \c$3164 ;
 wire \c$3166 ;
 wire \c$3168 ;
 wire \c$3170 ;
 wire \c$3172 ;
 wire \c$3174 ;
 wire \c$3176 ;
 wire \c$3178 ;
 wire \c$318 ;
 wire \c$3180 ;
 wire \c$3182 ;
 wire \c$3184 ;
 wire \c$3186 ;
 wire \c$3188 ;
 wire \c$3190 ;
 wire \c$3192 ;
 wire \c$3194 ;
 wire \c$3196 ;
 wire \c$3198 ;
 wire \c$32 ;
 wire \c$320 ;
 wire \c$3200 ;
 wire \c$3202 ;
 wire \c$3204 ;
 wire \c$3206 ;
 wire \c$3208 ;
 wire \c$3210 ;
 wire \c$3212 ;
 wire \c$3214 ;
 wire \c$3216 ;
 wire \c$3218 ;
 wire \c$322 ;
 wire \c$3220 ;
 wire \c$3222 ;
 wire \c$3224 ;
 wire \c$3226 ;
 wire \c$3228 ;
 wire \c$3230 ;
 wire \c$3232 ;
 wire \c$3234 ;
 wire \c$3236 ;
 wire \c$3238 ;
 wire \c$324 ;
 wire \c$3240 ;
 wire \c$3242 ;
 wire \c$3244 ;
 wire \c$3246 ;
 wire \c$3248 ;
 wire \c$3250 ;
 wire \c$3252 ;
 wire \c$3254 ;
 wire \c$3256 ;
 wire \c$3258 ;
 wire \c$326 ;
 wire \c$3260 ;
 wire \c$3262 ;
 wire \c$3264 ;
 wire \c$3266 ;
 wire \c$3268 ;
 wire \c$3270 ;
 wire \c$3272 ;
 wire \c$3274 ;
 wire \c$3276 ;
 wire \c$3278 ;
 wire \c$328 ;
 wire \c$3280 ;
 wire \c$3282 ;
 wire \c$3284 ;
 wire \c$3286 ;
 wire \c$3288 ;
 wire \c$3290 ;
 wire \c$3292 ;
 wire \c$3294 ;
 wire \c$3296 ;
 wire \c$3298 ;
 wire \c$330 ;
 wire \c$3300 ;
 wire \c$3302 ;
 wire \c$3304 ;
 wire \c$3306 ;
 wire \c$3308 ;
 wire \c$3310 ;
 wire \c$3312 ;
 wire \c$3314 ;
 wire \c$3316 ;
 wire \c$3318 ;
 wire \c$332 ;
 wire \c$3320 ;
 wire \c$3322 ;
 wire \c$3324 ;
 wire \c$3326 ;
 wire \c$3328 ;
 wire \c$3330 ;
 wire \c$3332 ;
 wire \c$3334 ;
 wire \c$3336 ;
 wire \c$3338 ;
 wire \c$334 ;
 wire \c$3340 ;
 wire \c$3342 ;
 wire \c$3344 ;
 wire \c$3346 ;
 wire \c$3348 ;
 wire \c$3350 ;
 wire \c$3352 ;
 wire \c$3354 ;
 wire \c$3356 ;
 wire \c$3358 ;
 wire \c$336 ;
 wire \c$3360 ;
 wire \c$3362 ;
 wire \c$3364 ;
 wire \c$3366 ;
 wire \c$3368 ;
 wire \c$3370 ;
 wire \c$3372 ;
 wire \c$3374 ;
 wire \c$3376 ;
 wire \c$3378 ;
 wire \c$338 ;
 wire \c$3380 ;
 wire \c$3382 ;
 wire \c$3384 ;
 wire \c$3386 ;
 wire \c$3388 ;
 wire \c$3390 ;
 wire \c$3392 ;
 wire \c$3394 ;
 wire \c$3396 ;
 wire \c$3398 ;
 wire \c$34 ;
 wire \c$340 ;
 wire \c$3400 ;
 wire \c$3402 ;
 wire \c$3404 ;
 wire \c$3406 ;
 wire \c$3408 ;
 wire \c$3410 ;
 wire \c$3412 ;
 wire \c$3414 ;
 wire \c$3416 ;
 wire \c$3418 ;
 wire \c$342 ;
 wire \c$3420 ;
 wire \c$3422 ;
 wire \c$3424 ;
 wire \c$3426 ;
 wire \c$3428 ;
 wire \c$3430 ;
 wire \c$3432 ;
 wire \c$3434 ;
 wire \c$3436 ;
 wire \c$3438 ;
 wire \c$344 ;
 wire \c$3440 ;
 wire \c$3442 ;
 wire \c$3444 ;
 wire \c$3446 ;
 wire \c$3448 ;
 wire \c$3450 ;
 wire \c$3452 ;
 wire \c$3454 ;
 wire \c$3456 ;
 wire \c$3458 ;
 wire \c$346 ;
 wire \c$3460 ;
 wire \c$3462 ;
 wire \c$3464 ;
 wire \c$3466 ;
 wire \c$3468 ;
 wire \c$3470 ;
 wire \c$3472 ;
 wire \c$3474 ;
 wire \c$3476 ;
 wire \c$3478 ;
 wire \c$348 ;
 wire \c$3480 ;
 wire \c$3482 ;
 wire \c$3484 ;
 wire \c$3486 ;
 wire \c$3488 ;
 wire \c$3490 ;
 wire \c$3492 ;
 wire \c$3494 ;
 wire \c$3496 ;
 wire \c$3498 ;
 wire \c$350 ;
 wire \c$3500 ;
 wire \c$3502 ;
 wire \c$3504 ;
 wire \c$3506 ;
 wire \c$3508 ;
 wire \c$3510 ;
 wire \c$3512 ;
 wire \c$3514 ;
 wire \c$3516 ;
 wire \c$3518 ;
 wire \c$352 ;
 wire \c$3520 ;
 wire \c$3522 ;
 wire \c$3524 ;
 wire \c$3526 ;
 wire \c$3528 ;
 wire \c$3530 ;
 wire \c$3532 ;
 wire \c$3534 ;
 wire \c$3536 ;
 wire \c$3538 ;
 wire \c$354 ;
 wire \c$3540 ;
 wire \c$3542 ;
 wire \c$3544 ;
 wire \c$3546 ;
 wire \c$3548 ;
 wire \c$3550 ;
 wire \c$3552 ;
 wire \c$3554 ;
 wire \c$3556 ;
 wire \c$3558 ;
 wire \c$356 ;
 wire \c$3560 ;
 wire \c$3562 ;
 wire \c$3564 ;
 wire \c$3566 ;
 wire \c$3568 ;
 wire \c$3570 ;
 wire \c$3572 ;
 wire \c$3574 ;
 wire \c$3576 ;
 wire \c$3578 ;
 wire \c$358 ;
 wire \c$3580 ;
 wire \c$3582 ;
 wire \c$3584 ;
 wire \c$3586 ;
 wire \c$3588 ;
 wire \c$3590 ;
 wire \c$3592 ;
 wire \c$3594 ;
 wire \c$3596 ;
 wire \c$3598 ;
 wire \c$36 ;
 wire \c$360 ;
 wire \c$3600 ;
 wire \c$3602 ;
 wire \c$3604 ;
 wire \c$3606 ;
 wire \c$3608 ;
 wire \c$3610 ;
 wire \c$3612 ;
 wire \c$3614 ;
 wire \c$3616 ;
 wire \c$3618 ;
 wire \c$362 ;
 wire \c$3620 ;
 wire \c$3622 ;
 wire \c$3624 ;
 wire \c$3626 ;
 wire \c$3628 ;
 wire \c$3630 ;
 wire \c$3632 ;
 wire \c$3634 ;
 wire \c$3636 ;
 wire \c$3638 ;
 wire \c$364 ;
 wire \c$3640 ;
 wire \c$3642 ;
 wire \c$3644 ;
 wire \c$3646 ;
 wire \c$3648 ;
 wire \c$3650 ;
 wire \c$3652 ;
 wire \c$3654 ;
 wire \c$3656 ;
 wire \c$3658 ;
 wire \c$366 ;
 wire \c$3660 ;
 wire \c$3662 ;
 wire \c$3664 ;
 wire \c$3666 ;
 wire \c$3668 ;
 wire \c$3670 ;
 wire \c$3672 ;
 wire \c$3674 ;
 wire \c$3676 ;
 wire \c$3678 ;
 wire \c$368 ;
 wire \c$3680 ;
 wire \c$3682 ;
 wire \c$3684 ;
 wire \c$3686 ;
 wire \c$3688 ;
 wire \c$3690 ;
 wire \c$3692 ;
 wire \c$3694 ;
 wire \c$3696 ;
 wire \c$3698 ;
 wire \c$370 ;
 wire \c$3700 ;
 wire \c$3702 ;
 wire \c$3704 ;
 wire \c$3706 ;
 wire \c$3708 ;
 wire \c$3710 ;
 wire \c$3712 ;
 wire \c$3714 ;
 wire \c$3716 ;
 wire \c$3718 ;
 wire \c$372 ;
 wire \c$3720 ;
 wire \c$3722 ;
 wire \c$3724 ;
 wire \c$3726 ;
 wire \c$3728 ;
 wire \c$3730 ;
 wire \c$3732 ;
 wire \c$3734 ;
 wire \c$3736 ;
 wire \c$3738 ;
 wire \c$374 ;
 wire \c$3740 ;
 wire \c$3742 ;
 wire \c$3744 ;
 wire \c$3746 ;
 wire \c$3748 ;
 wire \c$3750 ;
 wire \c$3752 ;
 wire \c$3754 ;
 wire \c$3756 ;
 wire \c$3758 ;
 wire \c$376 ;
 wire \c$3760 ;
 wire \c$3762 ;
 wire \c$3764 ;
 wire \c$3766 ;
 wire \c$3768 ;
 wire \c$3770 ;
 wire \c$3772 ;
 wire \c$3774 ;
 wire \c$3776 ;
 wire \c$3778 ;
 wire \c$378 ;
 wire \c$3780 ;
 wire \c$3782 ;
 wire \c$3784 ;
 wire \c$3786 ;
 wire \c$3788 ;
 wire \c$3790 ;
 wire \c$3792 ;
 wire \c$3794 ;
 wire \c$3796 ;
 wire \c$3798 ;
 wire \c$38 ;
 wire \c$380 ;
 wire \c$3800 ;
 wire \c$3802 ;
 wire \c$3804 ;
 wire \c$3806 ;
 wire \c$3808 ;
 wire \c$3810 ;
 wire \c$3812 ;
 wire \c$3814 ;
 wire \c$3816 ;
 wire \c$3818 ;
 wire \c$382 ;
 wire \c$3820 ;
 wire \c$3822 ;
 wire \c$3824 ;
 wire \c$3826 ;
 wire \c$3828 ;
 wire \c$3830 ;
 wire \c$3832 ;
 wire \c$3834 ;
 wire \c$3836 ;
 wire \c$3838 ;
 wire \c$384 ;
 wire \c$3840 ;
 wire \c$3842 ;
 wire \c$3844 ;
 wire \c$3846 ;
 wire \c$3848 ;
 wire \c$3850 ;
 wire \c$3852 ;
 wire \c$3854 ;
 wire \c$3856 ;
 wire \c$3858 ;
 wire \c$386 ;
 wire \c$3860 ;
 wire \c$3862 ;
 wire \c$3864 ;
 wire \c$3866 ;
 wire \c$3868 ;
 wire \c$3870 ;
 wire \c$3872 ;
 wire \c$3874 ;
 wire \c$3876 ;
 wire \c$3878 ;
 wire \c$388 ;
 wire \c$3880 ;
 wire \c$3882 ;
 wire \c$3884 ;
 wire \c$3886 ;
 wire \c$3888 ;
 wire \c$3890 ;
 wire \c$3892 ;
 wire \c$3894 ;
 wire \c$3896 ;
 wire \c$3898 ;
 wire \c$390 ;
 wire \c$3900 ;
 wire \c$3902 ;
 wire \c$3904 ;
 wire \c$3906 ;
 wire \c$3908 ;
 wire \c$3910 ;
 wire \c$3912 ;
 wire \c$3914 ;
 wire \c$3916 ;
 wire \c$3918 ;
 wire \c$392 ;
 wire \c$3920 ;
 wire \c$3922 ;
 wire \c$3924 ;
 wire \c$3926 ;
 wire \c$3928 ;
 wire \c$3930 ;
 wire \c$3932 ;
 wire \c$3934 ;
 wire \c$3936 ;
 wire \c$3938 ;
 wire \c$394 ;
 wire \c$3940 ;
 wire \c$3942 ;
 wire \c$3944 ;
 wire \c$3946 ;
 wire \c$3948 ;
 wire \c$3950 ;
 wire \c$3952 ;
 wire \c$3954 ;
 wire \c$3956 ;
 wire \c$3958 ;
 wire \c$396 ;
 wire \c$3960 ;
 wire \c$3962 ;
 wire \c$3964 ;
 wire \c$3966 ;
 wire \c$3968 ;
 wire \c$3970 ;
 wire \c$3972 ;
 wire \c$3974 ;
 wire \c$3976 ;
 wire \c$3978 ;
 wire \c$398 ;
 wire \c$3980 ;
 wire \c$3982 ;
 wire \c$3984 ;
 wire \c$3986 ;
 wire \c$3988 ;
 wire \c$3990 ;
 wire \c$3992 ;
 wire \c$3994 ;
 wire \c$3996 ;
 wire \c$3998 ;
 wire \c$4 ;
 wire \c$40 ;
 wire \c$400 ;
 wire \c$4000 ;
 wire \c$4002 ;
 wire \c$4004 ;
 wire \c$4006 ;
 wire \c$4008 ;
 wire \c$4010 ;
 wire \c$4012 ;
 wire \c$4014 ;
 wire \c$4016 ;
 wire \c$4018 ;
 wire \c$402 ;
 wire \c$4020 ;
 wire \c$4022 ;
 wire \c$4024 ;
 wire \c$4026 ;
 wire \c$4028 ;
 wire \c$4030 ;
 wire \c$4032 ;
 wire \c$4034 ;
 wire \c$4036 ;
 wire \c$4038 ;
 wire \c$404 ;
 wire \c$4040 ;
 wire \c$4042 ;
 wire \c$4044 ;
 wire \c$4046 ;
 wire \c$4048 ;
 wire \c$4050 ;
 wire \c$4052 ;
 wire \c$4054 ;
 wire \c$4056 ;
 wire \c$4058 ;
 wire \c$406 ;
 wire \c$4060 ;
 wire \c$4062 ;
 wire \c$4064 ;
 wire \c$4066 ;
 wire \c$4068 ;
 wire \c$4070 ;
 wire \c$4072 ;
 wire \c$4074 ;
 wire \c$4076 ;
 wire \c$4078 ;
 wire \c$408 ;
 wire \c$4080 ;
 wire \c$4082 ;
 wire \c$4084 ;
 wire \c$4086 ;
 wire \c$4088 ;
 wire \c$4090 ;
 wire \c$4092 ;
 wire \c$4094 ;
 wire \c$4096 ;
 wire \c$4098 ;
 wire \c$410 ;
 wire \c$4100 ;
 wire \c$4102 ;
 wire \c$4104 ;
 wire \c$4106 ;
 wire \c$4108 ;
 wire \c$4110 ;
 wire \c$4112 ;
 wire \c$4114 ;
 wire \c$4116 ;
 wire \c$4118 ;
 wire \c$412 ;
 wire \c$4120 ;
 wire \c$4122 ;
 wire \c$4124 ;
 wire \c$4126 ;
 wire \c$4128 ;
 wire \c$4130 ;
 wire \c$4132 ;
 wire \c$4134 ;
 wire \c$4136 ;
 wire \c$4138 ;
 wire \c$414 ;
 wire \c$4140 ;
 wire \c$4142 ;
 wire \c$4144 ;
 wire \c$4146 ;
 wire \c$4148 ;
 wire \c$4150 ;
 wire \c$4152 ;
 wire \c$4154 ;
 wire \c$4156 ;
 wire \c$4158 ;
 wire \c$416 ;
 wire \c$4160 ;
 wire \c$4162 ;
 wire \c$4164 ;
 wire \c$4166 ;
 wire \c$4168 ;
 wire \c$4170 ;
 wire \c$4172 ;
 wire \c$4174 ;
 wire \c$4176 ;
 wire \c$4178 ;
 wire \c$418 ;
 wire \c$4180 ;
 wire \c$4182 ;
 wire \c$4184 ;
 wire \c$4186 ;
 wire \c$4188 ;
 wire \c$4190 ;
 wire \c$4192 ;
 wire \c$4194 ;
 wire \c$4196 ;
 wire \c$4198 ;
 wire \c$42 ;
 wire \c$420 ;
 wire \c$4200 ;
 wire \c$4202 ;
 wire \c$4204 ;
 wire \c$4206 ;
 wire \c$4208 ;
 wire \c$4210 ;
 wire \c$4212 ;
 wire \c$4214 ;
 wire \c$4216 ;
 wire \c$4218 ;
 wire \c$422 ;
 wire \c$4220 ;
 wire \c$4222 ;
 wire \c$4224 ;
 wire \c$4226 ;
 wire \c$4228 ;
 wire \c$4230 ;
 wire \c$4232 ;
 wire \c$4234 ;
 wire \c$4236 ;
 wire \c$4238 ;
 wire \c$424 ;
 wire \c$4240 ;
 wire \c$4242 ;
 wire \c$4244 ;
 wire \c$4246 ;
 wire \c$4248 ;
 wire \c$4250 ;
 wire \c$4252 ;
 wire \c$4254 ;
 wire \c$4256 ;
 wire \c$4258 ;
 wire \c$426 ;
 wire \c$4260 ;
 wire \c$4262 ;
 wire \c$4264 ;
 wire \c$4266 ;
 wire \c$4268 ;
 wire \c$4270 ;
 wire \c$4272 ;
 wire \c$4274 ;
 wire \c$4276 ;
 wire \c$4278 ;
 wire \c$428 ;
 wire \c$4280 ;
 wire \c$4282 ;
 wire \c$4284 ;
 wire \c$4286 ;
 wire \c$4288 ;
 wire \c$4290 ;
 wire \c$4292 ;
 wire \c$4294 ;
 wire \c$4296 ;
 wire \c$4298 ;
 wire \c$430 ;
 wire \c$4300 ;
 wire \c$4302 ;
 wire \c$4304 ;
 wire \c$4306 ;
 wire \c$4308 ;
 wire \c$4310 ;
 wire \c$4312 ;
 wire \c$4314 ;
 wire \c$4316 ;
 wire \c$4318 ;
 wire \c$432 ;
 wire \c$4320 ;
 wire \c$4322 ;
 wire \c$4324 ;
 wire \c$4326 ;
 wire \c$4328 ;
 wire \c$4330 ;
 wire \c$4332 ;
 wire \c$4334 ;
 wire \c$4336 ;
 wire \c$4338 ;
 wire \c$434 ;
 wire \c$4340 ;
 wire \c$4342 ;
 wire \c$4344 ;
 wire \c$4346 ;
 wire \c$4348 ;
 wire \c$4350 ;
 wire \c$4352 ;
 wire \c$4354 ;
 wire \c$4356 ;
 wire \c$4358 ;
 wire \c$436 ;
 wire \c$4360 ;
 wire \c$4362 ;
 wire \c$4364 ;
 wire \c$4366 ;
 wire \c$4368 ;
 wire \c$4370 ;
 wire \c$4372 ;
 wire \c$4374 ;
 wire \c$4376 ;
 wire \c$4378 ;
 wire \c$438 ;
 wire \c$4380 ;
 wire \c$4382 ;
 wire \c$4384 ;
 wire \c$4386 ;
 wire \c$4388 ;
 wire \c$4390 ;
 wire \c$4392 ;
 wire \c$4394 ;
 wire \c$4396 ;
 wire \c$4398 ;
 wire \c$44 ;
 wire \c$440 ;
 wire \c$4400 ;
 wire \c$4402 ;
 wire \c$4404 ;
 wire \c$4406 ;
 wire \c$442 ;
 wire \c$444 ;
 wire \c$446 ;
 wire \c$448 ;
 wire \c$450 ;
 wire \c$452 ;
 wire \c$454 ;
 wire \c$456 ;
 wire \c$458 ;
 wire \c$46 ;
 wire \c$460 ;
 wire \c$462 ;
 wire \c$464 ;
 wire \c$466 ;
 wire \c$468 ;
 wire \c$470 ;
 wire \c$472 ;
 wire \c$474 ;
 wire \c$476 ;
 wire \c$478 ;
 wire \c$48 ;
 wire \c$480 ;
 wire \c$482 ;
 wire \c$484 ;
 wire \c$486 ;
 wire \c$488 ;
 wire \c$490 ;
 wire \c$492 ;
 wire \c$494 ;
 wire \c$496 ;
 wire \c$498 ;
 wire \c$50 ;
 wire \c$500 ;
 wire \c$502 ;
 wire \c$504 ;
 wire \c$506 ;
 wire \c$508 ;
 wire \c$510 ;
 wire \c$512 ;
 wire \c$514 ;
 wire \c$516 ;
 wire \c$518 ;
 wire \c$52 ;
 wire \c$520 ;
 wire \c$522 ;
 wire \c$524 ;
 wire \c$526 ;
 wire \c$528 ;
 wire \c$530 ;
 wire \c$532 ;
 wire \c$534 ;
 wire \c$536 ;
 wire \c$538 ;
 wire \c$54 ;
 wire \c$540 ;
 wire \c$542 ;
 wire \c$544 ;
 wire \c$546 ;
 wire \c$548 ;
 wire \c$550 ;
 wire \c$552 ;
 wire \c$554 ;
 wire \c$556 ;
 wire \c$558 ;
 wire \c$56 ;
 wire \c$560 ;
 wire \c$562 ;
 wire \c$564 ;
 wire \c$566 ;
 wire \c$568 ;
 wire \c$570 ;
 wire \c$572 ;
 wire \c$574 ;
 wire \c$576 ;
 wire \c$578 ;
 wire \c$58 ;
 wire \c$580 ;
 wire \c$582 ;
 wire \c$584 ;
 wire \c$586 ;
 wire \c$588 ;
 wire \c$590 ;
 wire \c$592 ;
 wire \c$594 ;
 wire \c$596 ;
 wire \c$598 ;
 wire \c$6 ;
 wire \c$60 ;
 wire \c$600 ;
 wire \c$602 ;
 wire \c$604 ;
 wire \c$606 ;
 wire \c$608 ;
 wire \c$610 ;
 wire \c$612 ;
 wire \c$614 ;
 wire \c$616 ;
 wire \c$618 ;
 wire \c$62 ;
 wire \c$620 ;
 wire \c$622 ;
 wire \c$624 ;
 wire \c$626 ;
 wire \c$628 ;
 wire \c$630 ;
 wire \c$632 ;
 wire \c$634 ;
 wire \c$636 ;
 wire \c$638 ;
 wire \c$64 ;
 wire \c$640 ;
 wire \c$642 ;
 wire \c$644 ;
 wire \c$646 ;
 wire \c$648 ;
 wire \c$650 ;
 wire \c$652 ;
 wire \c$654 ;
 wire \c$656 ;
 wire \c$658 ;
 wire \c$66 ;
 wire \c$660 ;
 wire \c$662 ;
 wire \c$664 ;
 wire \c$666 ;
 wire \c$668 ;
 wire \c$670 ;
 wire \c$672 ;
 wire \c$674 ;
 wire \c$676 ;
 wire \c$678 ;
 wire \c$68 ;
 wire \c$680 ;
 wire \c$682 ;
 wire \c$684 ;
 wire \c$686 ;
 wire \c$688 ;
 wire \c$690 ;
 wire \c$692 ;
 wire \c$694 ;
 wire \c$696 ;
 wire \c$698 ;
 wire \c$70 ;
 wire \c$700 ;
 wire \c$702 ;
 wire \c$704 ;
 wire \c$706 ;
 wire \c$708 ;
 wire \c$710 ;
 wire \c$712 ;
 wire \c$714 ;
 wire \c$716 ;
 wire \c$718 ;
 wire \c$72 ;
 wire \c$720 ;
 wire \c$722 ;
 wire \c$724 ;
 wire \c$726 ;
 wire \c$728 ;
 wire \c$730 ;
 wire \c$732 ;
 wire \c$734 ;
 wire \c$736 ;
 wire \c$738 ;
 wire \c$74 ;
 wire \c$740 ;
 wire \c$742 ;
 wire \c$744 ;
 wire \c$746 ;
 wire \c$748 ;
 wire \c$750 ;
 wire \c$752 ;
 wire \c$754 ;
 wire \c$756 ;
 wire \c$758 ;
 wire \c$76 ;
 wire \c$760 ;
 wire \c$762 ;
 wire \c$764 ;
 wire \c$766 ;
 wire \c$768 ;
 wire \c$770 ;
 wire \c$772 ;
 wire \c$774 ;
 wire \c$776 ;
 wire \c$778 ;
 wire \c$78 ;
 wire \c$780 ;
 wire \c$782 ;
 wire \c$784 ;
 wire \c$786 ;
 wire \c$788 ;
 wire \c$790 ;
 wire \c$792 ;
 wire \c$794 ;
 wire \c$796 ;
 wire \c$798 ;
 wire \c$8 ;
 wire \c$80 ;
 wire \c$800 ;
 wire \c$802 ;
 wire \c$804 ;
 wire \c$806 ;
 wire \c$808 ;
 wire \c$810 ;
 wire \c$812 ;
 wire \c$814 ;
 wire \c$816 ;
 wire \c$818 ;
 wire \c$82 ;
 wire \c$820 ;
 wire \c$822 ;
 wire \c$824 ;
 wire \c$826 ;
 wire \c$828 ;
 wire \c$830 ;
 wire \c$832 ;
 wire \c$834 ;
 wire \c$836 ;
 wire \c$838 ;
 wire \c$84 ;
 wire \c$840 ;
 wire \c$842 ;
 wire \c$844 ;
 wire \c$846 ;
 wire \c$848 ;
 wire \c$850 ;
 wire \c$852 ;
 wire \c$854 ;
 wire \c$856 ;
 wire \c$858 ;
 wire \c$86 ;
 wire \c$860 ;
 wire \c$862 ;
 wire \c$864 ;
 wire \c$866 ;
 wire \c$868 ;
 wire \c$870 ;
 wire \c$872 ;
 wire \c$874 ;
 wire \c$876 ;
 wire \c$878 ;
 wire \c$88 ;
 wire \c$880 ;
 wire \c$882 ;
 wire \c$884 ;
 wire \c$886 ;
 wire \c$888 ;
 wire \c$890 ;
 wire \c$892 ;
 wire \c$894 ;
 wire \c$896 ;
 wire \c$898 ;
 wire \c$90 ;
 wire \c$900 ;
 wire \c$902 ;
 wire \c$904 ;
 wire \c$906 ;
 wire \c$908 ;
 wire \c$910 ;
 wire \c$912 ;
 wire \c$914 ;
 wire \c$916 ;
 wire \c$918 ;
 wire \c$92 ;
 wire \c$920 ;
 wire \c$922 ;
 wire \c$924 ;
 wire \c$926 ;
 wire \c$928 ;
 wire \c$930 ;
 wire \c$932 ;
 wire \c$934 ;
 wire \c$936 ;
 wire \c$938 ;
 wire \c$94 ;
 wire \c$940 ;
 wire \c$942 ;
 wire \c$944 ;
 wire \c$946 ;
 wire \c$948 ;
 wire \c$950 ;
 wire \c$952 ;
 wire \c$954 ;
 wire \c$956 ;
 wire \c$958 ;
 wire \c$96 ;
 wire \c$960 ;
 wire \c$962 ;
 wire \c$964 ;
 wire \c$966 ;
 wire \c$968 ;
 wire \c$970 ;
 wire \c$972 ;
 wire \c$974 ;
 wire \c$976 ;
 wire \c$978 ;
 wire \c$98 ;
 wire \c$980 ;
 wire \c$982 ;
 wire \c$984 ;
 wire \c$986 ;
 wire \c$988 ;
 wire \c$990 ;
 wire \c$992 ;
 wire \c$994 ;
 wire \c$996 ;
 wire \c$998 ;
 wire \final_adder.$signal ;
 wire \final_adder.$signal$1 ;
 wire \final_adder.$signal$10 ;
 wire \final_adder.$signal$100 ;
 wire \final_adder.$signal$101 ;
 wire \final_adder.$signal$102 ;
 wire \final_adder.$signal$103 ;
 wire \final_adder.$signal$104 ;
 wire \final_adder.$signal$105 ;
 wire \final_adder.$signal$106 ;
 wire \final_adder.$signal$107 ;
 wire \final_adder.$signal$108 ;
 wire \final_adder.$signal$109 ;
 wire \final_adder.$signal$1091 ;
 wire \final_adder.$signal$1092 ;
 wire \final_adder.$signal$1093 ;
 wire \final_adder.$signal$1094 ;
 wire \final_adder.$signal$1095 ;
 wire \final_adder.$signal$1096 ;
 wire \final_adder.$signal$1097 ;
 wire \final_adder.$signal$1098 ;
 wire \final_adder.$signal$1099 ;
 wire \final_adder.$signal$110 ;
 wire \final_adder.$signal$1100 ;
 wire \final_adder.$signal$1101 ;
 wire \final_adder.$signal$1102 ;
 wire \final_adder.$signal$1103 ;
 wire \final_adder.$signal$1104 ;
 wire \final_adder.$signal$1105 ;
 wire \final_adder.$signal$1106 ;
 wire \final_adder.$signal$1107 ;
 wire \final_adder.$signal$1108 ;
 wire \final_adder.$signal$1109 ;
 wire \final_adder.$signal$111 ;
 wire \final_adder.$signal$1110 ;
 wire \final_adder.$signal$1111 ;
 wire \final_adder.$signal$1112 ;
 wire \final_adder.$signal$1113 ;
 wire \final_adder.$signal$1114 ;
 wire \final_adder.$signal$1115 ;
 wire \final_adder.$signal$1116 ;
 wire \final_adder.$signal$1117 ;
 wire \final_adder.$signal$1118 ;
 wire \final_adder.$signal$1119 ;
 wire \final_adder.$signal$112 ;
 wire \final_adder.$signal$1120 ;
 wire \final_adder.$signal$1121 ;
 wire \final_adder.$signal$1122 ;
 wire \final_adder.$signal$1123 ;
 wire \final_adder.$signal$1124 ;
 wire \final_adder.$signal$1125 ;
 wire \final_adder.$signal$1126 ;
 wire \final_adder.$signal$1127 ;
 wire \final_adder.$signal$1128 ;
 wire \final_adder.$signal$1129 ;
 wire \final_adder.$signal$113 ;
 wire \final_adder.$signal$1130 ;
 wire \final_adder.$signal$1131 ;
 wire \final_adder.$signal$1132 ;
 wire \final_adder.$signal$1133 ;
 wire \final_adder.$signal$1134 ;
 wire \final_adder.$signal$1135 ;
 wire \final_adder.$signal$1136 ;
 wire \final_adder.$signal$1137 ;
 wire \final_adder.$signal$1138 ;
 wire \final_adder.$signal$114 ;
 wire \final_adder.$signal$1146 ;
 wire \final_adder.$signal$1147 ;
 wire \final_adder.$signal$1148 ;
 wire \final_adder.$signal$1149 ;
 wire \final_adder.$signal$1150 ;
 wire \final_adder.$signal$1151 ;
 wire \final_adder.$signal$1152 ;
 wire \final_adder.$signal$1153 ;
 wire \final_adder.$signal$1154 ;
 wire \final_adder.$signal$1155 ;
 wire \final_adder.$signal$1156 ;
 wire \final_adder.$signal$1157 ;
 wire \final_adder.$signal$1158 ;
 wire \final_adder.$signal$1159 ;
 wire \final_adder.$signal$116 ;
 wire \final_adder.$signal$1160 ;
 wire \final_adder.$signal$1161 ;
 wire \final_adder.$signal$1162 ;
 wire \final_adder.$signal$1163 ;
 wire \final_adder.$signal$1164 ;
 wire \final_adder.$signal$1165 ;
 wire \final_adder.$signal$1166 ;
 wire \final_adder.$signal$1167 ;
 wire \final_adder.$signal$1168 ;
 wire \final_adder.$signal$1169 ;
 wire \final_adder.$signal$1170 ;
 wire \final_adder.$signal$1171 ;
 wire \final_adder.$signal$1172 ;
 wire \final_adder.$signal$1173 ;
 wire \final_adder.$signal$1174 ;
 wire \final_adder.$signal$1175 ;
 wire \final_adder.$signal$1176 ;
 wire \final_adder.$signal$1177 ;
 wire \final_adder.$signal$1178 ;
 wire \final_adder.$signal$1179 ;
 wire \final_adder.$signal$118 ;
 wire \final_adder.$signal$1180 ;
 wire \final_adder.$signal$1181 ;
 wire \final_adder.$signal$1182 ;
 wire \final_adder.$signal$1183 ;
 wire \final_adder.$signal$1184 ;
 wire \final_adder.$signal$1185 ;
 wire \final_adder.$signal$1186 ;
 wire \final_adder.$signal$1187 ;
 wire \final_adder.$signal$1188 ;
 wire \final_adder.$signal$1189 ;
 wire \final_adder.$signal$1190 ;
 wire \final_adder.$signal$1191 ;
 wire \final_adder.$signal$1192 ;
 wire \final_adder.$signal$1193 ;
 wire \final_adder.$signal$1194 ;
 wire \final_adder.$signal$1195 ;
 wire \final_adder.$signal$1196 ;
 wire \final_adder.$signal$1197 ;
 wire \final_adder.$signal$1198 ;
 wire \final_adder.$signal$1199 ;
 wire \final_adder.$signal$12 ;
 wire \final_adder.$signal$120 ;
 wire \final_adder.$signal$1200 ;
 wire \final_adder.$signal$1201 ;
 wire \final_adder.$signal$1202 ;
 wire \final_adder.$signal$1203 ;
 wire \final_adder.$signal$1204 ;
 wire \final_adder.$signal$1205 ;
 wire \final_adder.$signal$1206 ;
 wire \final_adder.$signal$1207 ;
 wire \final_adder.$signal$1208 ;
 wire \final_adder.$signal$1209 ;
 wire \final_adder.$signal$1210 ;
 wire \final_adder.$signal$1211 ;
 wire \final_adder.$signal$1212 ;
 wire \final_adder.$signal$1213 ;
 wire \final_adder.$signal$1214 ;
 wire \final_adder.$signal$1215 ;
 wire \final_adder.$signal$1216 ;
 wire \final_adder.$signal$1217 ;
 wire \final_adder.$signal$122 ;
 wire \final_adder.$signal$124 ;
 wire \final_adder.$signal$126 ;
 wire \final_adder.$signal$128 ;
 wire \final_adder.$signal$130 ;
 wire \final_adder.$signal$132 ;
 wire \final_adder.$signal$134 ;
 wire \final_adder.$signal$136 ;
 wire \final_adder.$signal$138 ;
 wire \final_adder.$signal$14 ;
 wire \final_adder.$signal$140 ;
 wire \final_adder.$signal$142 ;
 wire \final_adder.$signal$144 ;
 wire \final_adder.$signal$146 ;
 wire \final_adder.$signal$148 ;
 wire \final_adder.$signal$150 ;
 wire \final_adder.$signal$152 ;
 wire \final_adder.$signal$154 ;
 wire \final_adder.$signal$156 ;
 wire \final_adder.$signal$158 ;
 wire \final_adder.$signal$16 ;
 wire \final_adder.$signal$160 ;
 wire \final_adder.$signal$162 ;
 wire \final_adder.$signal$164 ;
 wire \final_adder.$signal$166 ;
 wire \final_adder.$signal$168 ;
 wire \final_adder.$signal$170 ;
 wire \final_adder.$signal$172 ;
 wire \final_adder.$signal$174 ;
 wire \final_adder.$signal$176 ;
 wire \final_adder.$signal$178 ;
 wire \final_adder.$signal$18 ;
 wire \final_adder.$signal$180 ;
 wire \final_adder.$signal$182 ;
 wire \final_adder.$signal$184 ;
 wire \final_adder.$signal$186 ;
 wire \final_adder.$signal$188 ;
 wire \final_adder.$signal$190 ;
 wire \final_adder.$signal$192 ;
 wire \final_adder.$signal$194 ;
 wire \final_adder.$signal$196 ;
 wire \final_adder.$signal$198 ;
 wire \final_adder.$signal$20 ;
 wire \final_adder.$signal$200 ;
 wire \final_adder.$signal$202 ;
 wire \final_adder.$signal$204 ;
 wire \final_adder.$signal$206 ;
 wire \final_adder.$signal$208 ;
 wire \final_adder.$signal$210 ;
 wire \final_adder.$signal$212 ;
 wire \final_adder.$signal$214 ;
 wire \final_adder.$signal$216 ;
 wire \final_adder.$signal$218 ;
 wire \final_adder.$signal$22 ;
 wire \final_adder.$signal$220 ;
 wire \final_adder.$signal$222 ;
 wire \final_adder.$signal$224 ;
 wire \final_adder.$signal$226 ;
 wire \final_adder.$signal$228 ;
 wire \final_adder.$signal$230 ;
 wire \final_adder.$signal$232 ;
 wire \final_adder.$signal$234 ;
 wire \final_adder.$signal$236 ;
 wire \final_adder.$signal$238 ;
 wire \final_adder.$signal$24 ;
 wire \final_adder.$signal$240 ;
 wire \final_adder.$signal$242 ;
 wire \final_adder.$signal$244 ;
 wire \final_adder.$signal$246 ;
 wire \final_adder.$signal$248 ;
 wire \final_adder.$signal$250 ;
 wire \final_adder.$signal$252 ;
 wire \final_adder.$signal$254 ;
 wire \final_adder.$signal$256 ;
 wire \final_adder.$signal$26 ;
 wire \final_adder.$signal$28 ;
 wire \final_adder.$signal$30 ;
 wire \final_adder.$signal$32 ;
 wire \final_adder.$signal$34 ;
 wire \final_adder.$signal$36 ;
 wire \final_adder.$signal$38 ;
 wire \final_adder.$signal$4 ;
 wire \final_adder.$signal$40 ;
 wire \final_adder.$signal$42 ;
 wire \final_adder.$signal$44 ;
 wire \final_adder.$signal$46 ;
 wire \final_adder.$signal$48 ;
 wire \final_adder.$signal$50 ;
 wire \final_adder.$signal$52 ;
 wire \final_adder.$signal$54 ;
 wire \final_adder.$signal$56 ;
 wire \final_adder.$signal$58 ;
 wire \final_adder.$signal$6 ;
 wire \final_adder.$signal$60 ;
 wire \final_adder.$signal$62 ;
 wire \final_adder.$signal$64 ;
 wire \final_adder.$signal$66 ;
 wire \final_adder.$signal$68 ;
 wire \final_adder.$signal$70 ;
 wire \final_adder.$signal$72 ;
 wire \final_adder.$signal$74 ;
 wire \final_adder.$signal$76 ;
 wire \final_adder.$signal$78 ;
 wire \final_adder.$signal$8 ;
 wire \final_adder.$signal$80 ;
 wire \final_adder.$signal$82 ;
 wire \final_adder.$signal$84 ;
 wire \final_adder.$signal$86 ;
 wire \final_adder.$signal$88 ;
 wire \final_adder.$signal$90 ;
 wire \final_adder.$signal$92 ;
 wire \final_adder.$signal$94 ;
 wire \final_adder.$signal$96 ;
 wire \final_adder.$signal$98 ;
 wire \final_adder.g_new$1001 ;
 wire \final_adder.g_new$1003 ;
 wire \final_adder.g_new$1005 ;
 wire \final_adder.g_new$1007 ;
 wire \final_adder.g_new$1009 ;
 wire \final_adder.g_new$1011 ;
 wire \final_adder.g_new$1013 ;
 wire \final_adder.g_new$1015 ;
 wire \final_adder.g_new$1017 ;
 wire \final_adder.g_new$1019 ;
 wire \final_adder.g_new$1021 ;
 wire \final_adder.g_new$1023 ;
 wire \final_adder.g_new$1025 ;
 wire \final_adder.g_new$1026 ;
 wire \final_adder.g_new$1027 ;
 wire \final_adder.g_new$1028 ;
 wire \final_adder.g_new$1029 ;
 wire \final_adder.g_new$1030 ;
 wire \final_adder.g_new$1031 ;
 wire \final_adder.g_new$1032 ;
 wire \final_adder.g_new$1033 ;
 wire \final_adder.g_new$1034 ;
 wire \final_adder.g_new$1035 ;
 wire \final_adder.g_new$1036 ;
 wire \final_adder.g_new$1037 ;
 wire \final_adder.g_new$1038 ;
 wire \final_adder.g_new$1039 ;
 wire \final_adder.g_new$1040 ;
 wire \final_adder.g_new$1041 ;
 wire \final_adder.g_new$1042 ;
 wire \final_adder.g_new$1043 ;
 wire \final_adder.g_new$1044 ;
 wire \final_adder.g_new$1045 ;
 wire \final_adder.g_new$1046 ;
 wire \final_adder.g_new$1047 ;
 wire \final_adder.g_new$1048 ;
 wire \final_adder.g_new$1049 ;
 wire \final_adder.g_new$1050 ;
 wire \final_adder.g_new$1051 ;
 wire \final_adder.g_new$1052 ;
 wire \final_adder.g_new$1053 ;
 wire \final_adder.g_new$1054 ;
 wire \final_adder.g_new$1055 ;
 wire \final_adder.g_new$1056 ;
 wire \final_adder.g_new$1057 ;
 wire \final_adder.g_new$1058 ;
 wire \final_adder.g_new$1059 ;
 wire \final_adder.g_new$1060 ;
 wire \final_adder.g_new$1061 ;
 wire \final_adder.g_new$1062 ;
 wire \final_adder.g_new$1063 ;
 wire \final_adder.g_new$1064 ;
 wire \final_adder.g_new$1065 ;
 wire \final_adder.g_new$1066 ;
 wire \final_adder.g_new$1067 ;
 wire \final_adder.g_new$1068 ;
 wire \final_adder.g_new$1069 ;
 wire \final_adder.g_new$1070 ;
 wire \final_adder.g_new$1071 ;
 wire \final_adder.g_new$1072 ;
 wire \final_adder.g_new$1073 ;
 wire \final_adder.g_new$1074 ;
 wire \final_adder.g_new$1075 ;
 wire \final_adder.g_new$1076 ;
 wire \final_adder.g_new$1077 ;
 wire \final_adder.g_new$1078 ;
 wire \final_adder.g_new$1079 ;
 wire \final_adder.g_new$1080 ;
 wire \final_adder.g_new$1081 ;
 wire \final_adder.g_new$1082 ;
 wire \final_adder.g_new$1083 ;
 wire \final_adder.g_new$1084 ;
 wire \final_adder.g_new$1085 ;
 wire \final_adder.g_new$1086 ;
 wire \final_adder.g_new$1087 ;
 wire \final_adder.g_new$1088 ;
 wire \final_adder.g_new$259 ;
 wire \final_adder.g_new$261 ;
 wire \final_adder.g_new$263 ;
 wire \final_adder.g_new$265 ;
 wire \final_adder.g_new$267 ;
 wire \final_adder.g_new$269 ;
 wire \final_adder.g_new$271 ;
 wire \final_adder.g_new$273 ;
 wire \final_adder.g_new$275 ;
 wire \final_adder.g_new$277 ;
 wire \final_adder.g_new$279 ;
 wire \final_adder.g_new$281 ;
 wire \final_adder.g_new$283 ;
 wire \final_adder.g_new$285 ;
 wire \final_adder.g_new$287 ;
 wire \final_adder.g_new$289 ;
 wire \final_adder.g_new$291 ;
 wire \final_adder.g_new$293 ;
 wire \final_adder.g_new$295 ;
 wire \final_adder.g_new$297 ;
 wire \final_adder.g_new$299 ;
 wire \final_adder.g_new$301 ;
 wire \final_adder.g_new$303 ;
 wire \final_adder.g_new$305 ;
 wire \final_adder.g_new$307 ;
 wire \final_adder.g_new$309 ;
 wire \final_adder.g_new$311 ;
 wire \final_adder.g_new$313 ;
 wire \final_adder.g_new$315 ;
 wire \final_adder.g_new$317 ;
 wire \final_adder.g_new$319 ;
 wire \final_adder.g_new$321 ;
 wire \final_adder.g_new$323 ;
 wire \final_adder.g_new$325 ;
 wire \final_adder.g_new$327 ;
 wire \final_adder.g_new$329 ;
 wire \final_adder.g_new$331 ;
 wire \final_adder.g_new$333 ;
 wire \final_adder.g_new$335 ;
 wire \final_adder.g_new$337 ;
 wire \final_adder.g_new$339 ;
 wire \final_adder.g_new$341 ;
 wire \final_adder.g_new$343 ;
 wire \final_adder.g_new$345 ;
 wire \final_adder.g_new$347 ;
 wire \final_adder.g_new$349 ;
 wire \final_adder.g_new$351 ;
 wire \final_adder.g_new$353 ;
 wire \final_adder.g_new$355 ;
 wire \final_adder.g_new$357 ;
 wire \final_adder.g_new$359 ;
 wire \final_adder.g_new$361 ;
 wire \final_adder.g_new$363 ;
 wire \final_adder.g_new$365 ;
 wire \final_adder.g_new$367 ;
 wire \final_adder.g_new$369 ;
 wire \final_adder.g_new$371 ;
 wire \final_adder.g_new$373 ;
 wire \final_adder.g_new$375 ;
 wire \final_adder.g_new$377 ;
 wire \final_adder.g_new$379 ;
 wire \final_adder.g_new$381 ;
 wire \final_adder.g_new$383 ;
 wire \final_adder.g_new$387 ;
 wire \final_adder.g_new$389 ;
 wire \final_adder.g_new$391 ;
 wire \final_adder.g_new$393 ;
 wire \final_adder.g_new$395 ;
 wire \final_adder.g_new$397 ;
 wire \final_adder.g_new$399 ;
 wire \final_adder.g_new$401 ;
 wire \final_adder.g_new$403 ;
 wire \final_adder.g_new$405 ;
 wire \final_adder.g_new$407 ;
 wire \final_adder.g_new$409 ;
 wire \final_adder.g_new$411 ;
 wire \final_adder.g_new$413 ;
 wire \final_adder.g_new$415 ;
 wire \final_adder.g_new$417 ;
 wire \final_adder.g_new$419 ;
 wire \final_adder.g_new$421 ;
 wire \final_adder.g_new$423 ;
 wire \final_adder.g_new$425 ;
 wire \final_adder.g_new$427 ;
 wire \final_adder.g_new$429 ;
 wire \final_adder.g_new$431 ;
 wire \final_adder.g_new$433 ;
 wire \final_adder.g_new$435 ;
 wire \final_adder.g_new$437 ;
 wire \final_adder.g_new$439 ;
 wire \final_adder.g_new$441 ;
 wire \final_adder.g_new$443 ;
 wire \final_adder.g_new$445 ;
 wire \final_adder.g_new$447 ;
 wire \final_adder.g_new$449 ;
 wire \final_adder.g_new$451 ;
 wire \final_adder.g_new$453 ;
 wire \final_adder.g_new$455 ;
 wire \final_adder.g_new$457 ;
 wire \final_adder.g_new$459 ;
 wire \final_adder.g_new$461 ;
 wire \final_adder.g_new$463 ;
 wire \final_adder.g_new$465 ;
 wire \final_adder.g_new$467 ;
 wire \final_adder.g_new$469 ;
 wire \final_adder.g_new$471 ;
 wire \final_adder.g_new$473 ;
 wire \final_adder.g_new$475 ;
 wire \final_adder.g_new$477 ;
 wire \final_adder.g_new$479 ;
 wire \final_adder.g_new$481 ;
 wire \final_adder.g_new$483 ;
 wire \final_adder.g_new$485 ;
 wire \final_adder.g_new$487 ;
 wire \final_adder.g_new$489 ;
 wire \final_adder.g_new$491 ;
 wire \final_adder.g_new$493 ;
 wire \final_adder.g_new$495 ;
 wire \final_adder.g_new$497 ;
 wire \final_adder.g_new$499 ;
 wire \final_adder.g_new$501 ;
 wire \final_adder.g_new$503 ;
 wire \final_adder.g_new$505 ;
 wire \final_adder.g_new$507 ;
 wire \final_adder.g_new$509 ;
 wire \final_adder.g_new$513 ;
 wire \final_adder.g_new$515 ;
 wire \final_adder.g_new$517 ;
 wire \final_adder.g_new$519 ;
 wire \final_adder.g_new$521 ;
 wire \final_adder.g_new$523 ;
 wire \final_adder.g_new$525 ;
 wire \final_adder.g_new$527 ;
 wire \final_adder.g_new$529 ;
 wire \final_adder.g_new$531 ;
 wire \final_adder.g_new$533 ;
 wire \final_adder.g_new$535 ;
 wire \final_adder.g_new$537 ;
 wire \final_adder.g_new$539 ;
 wire \final_adder.g_new$541 ;
 wire \final_adder.g_new$543 ;
 wire \final_adder.g_new$545 ;
 wire \final_adder.g_new$547 ;
 wire \final_adder.g_new$549 ;
 wire \final_adder.g_new$551 ;
 wire \final_adder.g_new$553 ;
 wire \final_adder.g_new$555 ;
 wire \final_adder.g_new$557 ;
 wire \final_adder.g_new$559 ;
 wire \final_adder.g_new$561 ;
 wire \final_adder.g_new$563 ;
 wire \final_adder.g_new$565 ;
 wire \final_adder.g_new$567 ;
 wire \final_adder.g_new$569 ;
 wire \final_adder.g_new$571 ;
 wire \final_adder.g_new$573 ;
 wire \final_adder.g_new$575 ;
 wire \final_adder.g_new$577 ;
 wire \final_adder.g_new$579 ;
 wire \final_adder.g_new$581 ;
 wire \final_adder.g_new$583 ;
 wire \final_adder.g_new$585 ;
 wire \final_adder.g_new$587 ;
 wire \final_adder.g_new$589 ;
 wire \final_adder.g_new$591 ;
 wire \final_adder.g_new$593 ;
 wire \final_adder.g_new$595 ;
 wire \final_adder.g_new$597 ;
 wire \final_adder.g_new$599 ;
 wire \final_adder.g_new$601 ;
 wire \final_adder.g_new$603 ;
 wire \final_adder.g_new$605 ;
 wire \final_adder.g_new$607 ;
 wire \final_adder.g_new$609 ;
 wire \final_adder.g_new$611 ;
 wire \final_adder.g_new$613 ;
 wire \final_adder.g_new$615 ;
 wire \final_adder.g_new$617 ;
 wire \final_adder.g_new$619 ;
 wire \final_adder.g_new$621 ;
 wire \final_adder.g_new$623 ;
 wire \final_adder.g_new$625 ;
 wire \final_adder.g_new$627 ;
 wire \final_adder.g_new$629 ;
 wire \final_adder.g_new$631 ;
 wire \final_adder.g_new$633 ;
 wire \final_adder.g_new$637 ;
 wire \final_adder.g_new$639 ;
 wire \final_adder.g_new$641 ;
 wire \final_adder.g_new$643 ;
 wire \final_adder.g_new$645 ;
 wire \final_adder.g_new$647 ;
 wire \final_adder.g_new$649 ;
 wire \final_adder.g_new$651 ;
 wire \final_adder.g_new$653 ;
 wire \final_adder.g_new$655 ;
 wire \final_adder.g_new$657 ;
 wire \final_adder.g_new$659 ;
 wire \final_adder.g_new$661 ;
 wire \final_adder.g_new$663 ;
 wire \final_adder.g_new$665 ;
 wire \final_adder.g_new$667 ;
 wire \final_adder.g_new$669 ;
 wire \final_adder.g_new$671 ;
 wire \final_adder.g_new$673 ;
 wire \final_adder.g_new$675 ;
 wire \final_adder.g_new$677 ;
 wire \final_adder.g_new$679 ;
 wire \final_adder.g_new$681 ;
 wire \final_adder.g_new$683 ;
 wire \final_adder.g_new$685 ;
 wire \final_adder.g_new$687 ;
 wire \final_adder.g_new$689 ;
 wire \final_adder.g_new$691 ;
 wire \final_adder.g_new$693 ;
 wire \final_adder.g_new$695 ;
 wire \final_adder.g_new$697 ;
 wire \final_adder.g_new$699 ;
 wire \final_adder.g_new$701 ;
 wire \final_adder.g_new$703 ;
 wire \final_adder.g_new$705 ;
 wire \final_adder.g_new$707 ;
 wire \final_adder.g_new$709 ;
 wire \final_adder.g_new$711 ;
 wire \final_adder.g_new$713 ;
 wire \final_adder.g_new$715 ;
 wire \final_adder.g_new$717 ;
 wire \final_adder.g_new$719 ;
 wire \final_adder.g_new$721 ;
 wire \final_adder.g_new$723 ;
 wire \final_adder.g_new$725 ;
 wire \final_adder.g_new$727 ;
 wire \final_adder.g_new$729 ;
 wire \final_adder.g_new$731 ;
 wire \final_adder.g_new$733 ;
 wire \final_adder.g_new$735 ;
 wire \final_adder.g_new$737 ;
 wire \final_adder.g_new$739 ;
 wire \final_adder.g_new$741 ;
 wire \final_adder.g_new$743 ;
 wire \final_adder.g_new$745 ;
 wire \final_adder.g_new$747 ;
 wire \final_adder.g_new$749 ;
 wire \final_adder.g_new$751 ;
 wire \final_adder.g_new$753 ;
 wire \final_adder.g_new$757 ;
 wire \final_adder.g_new$759 ;
 wire \final_adder.g_new$761 ;
 wire \final_adder.g_new$763 ;
 wire \final_adder.g_new$765 ;
 wire \final_adder.g_new$767 ;
 wire \final_adder.g_new$769 ;
 wire \final_adder.g_new$771 ;
 wire \final_adder.g_new$773 ;
 wire \final_adder.g_new$775 ;
 wire \final_adder.g_new$777 ;
 wire \final_adder.g_new$779 ;
 wire \final_adder.g_new$781 ;
 wire \final_adder.g_new$783 ;
 wire \final_adder.g_new$785 ;
 wire \final_adder.g_new$787 ;
 wire \final_adder.g_new$789 ;
 wire \final_adder.g_new$791 ;
 wire \final_adder.g_new$793 ;
 wire \final_adder.g_new$795 ;
 wire \final_adder.g_new$797 ;
 wire \final_adder.g_new$799 ;
 wire \final_adder.g_new$801 ;
 wire \final_adder.g_new$803 ;
 wire \final_adder.g_new$805 ;
 wire \final_adder.g_new$807 ;
 wire \final_adder.g_new$809 ;
 wire \final_adder.g_new$811 ;
 wire \final_adder.g_new$813 ;
 wire \final_adder.g_new$815 ;
 wire \final_adder.g_new$817 ;
 wire \final_adder.g_new$819 ;
 wire \final_adder.g_new$821 ;
 wire \final_adder.g_new$823 ;
 wire \final_adder.g_new$825 ;
 wire \final_adder.g_new$827 ;
 wire \final_adder.g_new$829 ;
 wire \final_adder.g_new$831 ;
 wire \final_adder.g_new$833 ;
 wire \final_adder.g_new$835 ;
 wire \final_adder.g_new$837 ;
 wire \final_adder.g_new$839 ;
 wire \final_adder.g_new$841 ;
 wire \final_adder.g_new$843 ;
 wire \final_adder.g_new$845 ;
 wire \final_adder.g_new$847 ;
 wire \final_adder.g_new$849 ;
 wire \final_adder.g_new$851 ;
 wire \final_adder.g_new$853 ;
 wire \final_adder.g_new$855 ;
 wire \final_adder.g_new$857 ;
 wire \final_adder.g_new$859 ;
 wire \final_adder.g_new$861 ;
 wire \final_adder.g_new$863 ;
 wire \final_adder.g_new$865 ;
 wire \final_adder.g_new$869 ;
 wire \final_adder.g_new$871 ;
 wire \final_adder.g_new$873 ;
 wire \final_adder.g_new$875 ;
 wire \final_adder.g_new$877 ;
 wire \final_adder.g_new$879 ;
 wire \final_adder.g_new$881 ;
 wire \final_adder.g_new$883 ;
 wire \final_adder.g_new$885 ;
 wire \final_adder.g_new$887 ;
 wire \final_adder.g_new$889 ;
 wire \final_adder.g_new$891 ;
 wire \final_adder.g_new$893 ;
 wire \final_adder.g_new$895 ;
 wire \final_adder.g_new$897 ;
 wire \final_adder.g_new$899 ;
 wire \final_adder.g_new$901 ;
 wire \final_adder.g_new$903 ;
 wire \final_adder.g_new$905 ;
 wire \final_adder.g_new$907 ;
 wire \final_adder.g_new$909 ;
 wire \final_adder.g_new$911 ;
 wire \final_adder.g_new$913 ;
 wire \final_adder.g_new$915 ;
 wire \final_adder.g_new$917 ;
 wire \final_adder.g_new$919 ;
 wire \final_adder.g_new$921 ;
 wire \final_adder.g_new$923 ;
 wire \final_adder.g_new$925 ;
 wire \final_adder.g_new$927 ;
 wire \final_adder.g_new$929 ;
 wire \final_adder.g_new$931 ;
 wire \final_adder.g_new$933 ;
 wire \final_adder.g_new$935 ;
 wire \final_adder.g_new$937 ;
 wire \final_adder.g_new$939 ;
 wire \final_adder.g_new$941 ;
 wire \final_adder.g_new$943 ;
 wire \final_adder.g_new$945 ;
 wire \final_adder.g_new$947 ;
 wire \final_adder.g_new$949 ;
 wire \final_adder.g_new$951 ;
 wire \final_adder.g_new$953 ;
 wire \final_adder.g_new$955 ;
 wire \final_adder.g_new$957 ;
 wire \final_adder.g_new$959 ;
 wire \final_adder.g_new$961 ;
 wire \final_adder.g_new$965 ;
 wire \final_adder.g_new$967 ;
 wire \final_adder.g_new$969 ;
 wire \final_adder.g_new$971 ;
 wire \final_adder.g_new$973 ;
 wire \final_adder.g_new$975 ;
 wire \final_adder.g_new$977 ;
 wire \final_adder.g_new$979 ;
 wire \final_adder.g_new$981 ;
 wire \final_adder.g_new$983 ;
 wire \final_adder.g_new$985 ;
 wire \final_adder.g_new$987 ;
 wire \final_adder.g_new$989 ;
 wire \final_adder.g_new$991 ;
 wire \final_adder.g_new$993 ;
 wire \final_adder.g_new$995 ;
 wire \final_adder.g_new$997 ;
 wire \final_adder.g_new$999 ;
 wire \final_adder.p_new$258 ;
 wire \final_adder.p_new$260 ;
 wire \final_adder.p_new$262 ;
 wire \final_adder.p_new$264 ;
 wire \final_adder.p_new$266 ;
 wire \final_adder.p_new$268 ;
 wire \final_adder.p_new$270 ;
 wire \final_adder.p_new$272 ;
 wire \final_adder.p_new$274 ;
 wire \final_adder.p_new$276 ;
 wire \final_adder.p_new$278 ;
 wire \final_adder.p_new$280 ;
 wire \final_adder.p_new$282 ;
 wire \final_adder.p_new$284 ;
 wire \final_adder.p_new$286 ;
 wire \final_adder.p_new$288 ;
 wire \final_adder.p_new$290 ;
 wire \final_adder.p_new$292 ;
 wire \final_adder.p_new$294 ;
 wire \final_adder.p_new$296 ;
 wire \final_adder.p_new$298 ;
 wire \final_adder.p_new$300 ;
 wire \final_adder.p_new$302 ;
 wire \final_adder.p_new$304 ;
 wire \final_adder.p_new$306 ;
 wire \final_adder.p_new$308 ;
 wire \final_adder.p_new$310 ;
 wire \final_adder.p_new$312 ;
 wire \final_adder.p_new$314 ;
 wire \final_adder.p_new$316 ;
 wire \final_adder.p_new$318 ;
 wire \final_adder.p_new$320 ;
 wire \final_adder.p_new$322 ;
 wire \final_adder.p_new$324 ;
 wire \final_adder.p_new$326 ;
 wire \final_adder.p_new$328 ;
 wire \final_adder.p_new$330 ;
 wire \final_adder.p_new$332 ;
 wire \final_adder.p_new$334 ;
 wire \final_adder.p_new$336 ;
 wire \final_adder.p_new$338 ;
 wire \final_adder.p_new$340 ;
 wire \final_adder.p_new$342 ;
 wire \final_adder.p_new$344 ;
 wire \final_adder.p_new$346 ;
 wire \final_adder.p_new$348 ;
 wire \final_adder.p_new$350 ;
 wire \final_adder.p_new$352 ;
 wire \final_adder.p_new$354 ;
 wire \final_adder.p_new$356 ;
 wire \final_adder.p_new$358 ;
 wire \final_adder.p_new$360 ;
 wire \final_adder.p_new$362 ;
 wire \final_adder.p_new$364 ;
 wire \final_adder.p_new$366 ;
 wire \final_adder.p_new$368 ;
 wire \final_adder.p_new$370 ;
 wire \final_adder.p_new$372 ;
 wire \final_adder.p_new$374 ;
 wire \final_adder.p_new$376 ;
 wire \final_adder.p_new$378 ;
 wire \final_adder.p_new$380 ;
 wire \final_adder.p_new$386 ;
 wire \final_adder.p_new$388 ;
 wire \final_adder.p_new$390 ;
 wire \final_adder.p_new$392 ;
 wire \final_adder.p_new$394 ;
 wire \final_adder.p_new$396 ;
 wire \final_adder.p_new$398 ;
 wire \final_adder.p_new$400 ;
 wire \final_adder.p_new$402 ;
 wire \final_adder.p_new$404 ;
 wire \final_adder.p_new$406 ;
 wire \final_adder.p_new$408 ;
 wire \final_adder.p_new$410 ;
 wire \final_adder.p_new$412 ;
 wire \final_adder.p_new$414 ;
 wire \final_adder.p_new$416 ;
 wire \final_adder.p_new$418 ;
 wire \final_adder.p_new$420 ;
 wire \final_adder.p_new$422 ;
 wire \final_adder.p_new$424 ;
 wire \final_adder.p_new$426 ;
 wire \final_adder.p_new$428 ;
 wire \final_adder.p_new$430 ;
 wire \final_adder.p_new$432 ;
 wire \final_adder.p_new$434 ;
 wire \final_adder.p_new$436 ;
 wire \final_adder.p_new$438 ;
 wire \final_adder.p_new$440 ;
 wire \final_adder.p_new$442 ;
 wire \final_adder.p_new$444 ;
 wire \final_adder.p_new$446 ;
 wire \final_adder.p_new$448 ;
 wire \final_adder.p_new$450 ;
 wire \final_adder.p_new$452 ;
 wire \final_adder.p_new$454 ;
 wire \final_adder.p_new$456 ;
 wire \final_adder.p_new$458 ;
 wire \final_adder.p_new$460 ;
 wire \final_adder.p_new$462 ;
 wire \final_adder.p_new$464 ;
 wire \final_adder.p_new$466 ;
 wire \final_adder.p_new$468 ;
 wire \final_adder.p_new$470 ;
 wire \final_adder.p_new$472 ;
 wire \final_adder.p_new$474 ;
 wire \final_adder.p_new$476 ;
 wire \final_adder.p_new$478 ;
 wire \final_adder.p_new$480 ;
 wire \final_adder.p_new$482 ;
 wire \final_adder.p_new$484 ;
 wire \final_adder.p_new$486 ;
 wire \final_adder.p_new$488 ;
 wire \final_adder.p_new$490 ;
 wire \final_adder.p_new$492 ;
 wire \final_adder.p_new$494 ;
 wire \final_adder.p_new$496 ;
 wire \final_adder.p_new$498 ;
 wire \final_adder.p_new$500 ;
 wire \final_adder.p_new$502 ;
 wire \final_adder.p_new$504 ;
 wire \final_adder.p_new$506 ;
 wire \final_adder.p_new$512 ;
 wire \final_adder.p_new$514 ;
 wire \final_adder.p_new$516 ;
 wire \final_adder.p_new$518 ;
 wire \final_adder.p_new$520 ;
 wire \final_adder.p_new$522 ;
 wire \final_adder.p_new$524 ;
 wire \final_adder.p_new$526 ;
 wire \final_adder.p_new$528 ;
 wire \final_adder.p_new$530 ;
 wire \final_adder.p_new$532 ;
 wire \final_adder.p_new$534 ;
 wire \final_adder.p_new$536 ;
 wire \final_adder.p_new$538 ;
 wire \final_adder.p_new$540 ;
 wire \final_adder.p_new$542 ;
 wire \final_adder.p_new$544 ;
 wire \final_adder.p_new$546 ;
 wire \final_adder.p_new$548 ;
 wire \final_adder.p_new$550 ;
 wire \final_adder.p_new$552 ;
 wire \final_adder.p_new$554 ;
 wire \final_adder.p_new$556 ;
 wire \final_adder.p_new$558 ;
 wire \final_adder.p_new$560 ;
 wire \final_adder.p_new$562 ;
 wire \final_adder.p_new$564 ;
 wire \final_adder.p_new$566 ;
 wire \final_adder.p_new$568 ;
 wire \final_adder.p_new$570 ;
 wire \final_adder.p_new$572 ;
 wire \final_adder.p_new$574 ;
 wire \final_adder.p_new$576 ;
 wire \final_adder.p_new$578 ;
 wire \final_adder.p_new$580 ;
 wire \final_adder.p_new$582 ;
 wire \final_adder.p_new$584 ;
 wire \final_adder.p_new$586 ;
 wire \final_adder.p_new$588 ;
 wire \final_adder.p_new$590 ;
 wire \final_adder.p_new$592 ;
 wire \final_adder.p_new$594 ;
 wire \final_adder.p_new$596 ;
 wire \final_adder.p_new$598 ;
 wire \final_adder.p_new$600 ;
 wire \final_adder.p_new$602 ;
 wire \final_adder.p_new$604 ;
 wire \final_adder.p_new$606 ;
 wire \final_adder.p_new$608 ;
 wire \final_adder.p_new$610 ;
 wire \final_adder.p_new$612 ;
 wire \final_adder.p_new$614 ;
 wire \final_adder.p_new$616 ;
 wire \final_adder.p_new$618 ;
 wire \final_adder.p_new$620 ;
 wire \final_adder.p_new$622 ;
 wire \final_adder.p_new$624 ;
 wire \final_adder.p_new$626 ;
 wire \final_adder.p_new$628 ;
 wire \final_adder.p_new$636 ;
 wire \final_adder.p_new$638 ;
 wire \final_adder.p_new$640 ;
 wire \final_adder.p_new$642 ;
 wire \final_adder.p_new$644 ;
 wire \final_adder.p_new$646 ;
 wire \final_adder.p_new$648 ;
 wire \final_adder.p_new$650 ;
 wire \final_adder.p_new$652 ;
 wire \final_adder.p_new$654 ;
 wire \final_adder.p_new$656 ;
 wire \final_adder.p_new$658 ;
 wire \final_adder.p_new$660 ;
 wire \final_adder.p_new$662 ;
 wire \final_adder.p_new$664 ;
 wire \final_adder.p_new$666 ;
 wire \final_adder.p_new$668 ;
 wire \final_adder.p_new$670 ;
 wire \final_adder.p_new$672 ;
 wire \final_adder.p_new$674 ;
 wire \final_adder.p_new$676 ;
 wire \final_adder.p_new$678 ;
 wire \final_adder.p_new$680 ;
 wire \final_adder.p_new$682 ;
 wire \final_adder.p_new$684 ;
 wire \final_adder.p_new$686 ;
 wire \final_adder.p_new$688 ;
 wire \final_adder.p_new$690 ;
 wire \final_adder.p_new$692 ;
 wire \final_adder.p_new$694 ;
 wire \final_adder.p_new$696 ;
 wire \final_adder.p_new$698 ;
 wire \final_adder.p_new$700 ;
 wire \final_adder.p_new$702 ;
 wire \final_adder.p_new$704 ;
 wire \final_adder.p_new$706 ;
 wire \final_adder.p_new$708 ;
 wire \final_adder.p_new$710 ;
 wire \final_adder.p_new$712 ;
 wire \final_adder.p_new$714 ;
 wire \final_adder.p_new$716 ;
 wire \final_adder.p_new$718 ;
 wire \final_adder.p_new$720 ;
 wire \final_adder.p_new$722 ;
 wire \final_adder.p_new$724 ;
 wire \final_adder.p_new$726 ;
 wire \final_adder.p_new$728 ;
 wire \final_adder.p_new$730 ;
 wire \final_adder.p_new$732 ;
 wire \final_adder.p_new$734 ;
 wire \final_adder.p_new$736 ;
 wire \final_adder.p_new$738 ;
 wire \final_adder.p_new$740 ;
 wire \final_adder.p_new$742 ;
 wire \final_adder.p_new$744 ;
 wire \final_adder.p_new$756 ;
 wire \final_adder.p_new$758 ;
 wire \final_adder.p_new$760 ;
 wire \final_adder.p_new$762 ;
 wire \final_adder.p_new$764 ;
 wire \final_adder.p_new$766 ;
 wire \final_adder.p_new$768 ;
 wire \final_adder.p_new$770 ;
 wire \final_adder.p_new$772 ;
 wire \final_adder.p_new$774 ;
 wire \final_adder.p_new$776 ;
 wire \final_adder.p_new$778 ;
 wire \final_adder.p_new$780 ;
 wire \final_adder.p_new$782 ;
 wire \final_adder.p_new$784 ;
 wire \final_adder.p_new$786 ;
 wire \final_adder.p_new$788 ;
 wire \final_adder.p_new$790 ;
 wire \final_adder.p_new$792 ;
 wire \final_adder.p_new$794 ;
 wire \final_adder.p_new$796 ;
 wire \final_adder.p_new$798 ;
 wire \final_adder.p_new$800 ;
 wire \final_adder.p_new$802 ;
 wire \final_adder.p_new$804 ;
 wire \final_adder.p_new$806 ;
 wire \final_adder.p_new$808 ;
 wire \final_adder.p_new$810 ;
 wire \final_adder.p_new$812 ;
 wire \final_adder.p_new$814 ;
 wire \final_adder.p_new$816 ;
 wire \final_adder.p_new$818 ;
 wire \final_adder.p_new$820 ;
 wire \final_adder.p_new$822 ;
 wire \final_adder.p_new$824 ;
 wire \final_adder.p_new$826 ;
 wire \final_adder.p_new$828 ;
 wire \final_adder.p_new$830 ;
 wire \final_adder.p_new$832 ;
 wire \final_adder.p_new$834 ;
 wire \final_adder.p_new$836 ;
 wire \final_adder.p_new$838 ;
 wire \final_adder.p_new$840 ;
 wire \final_adder.p_new$842 ;
 wire \final_adder.p_new$844 ;
 wire \final_adder.p_new$846 ;
 wire \final_adder.p_new$848 ;
 wire \final_adder.p_new$868 ;
 wire \final_adder.p_new$870 ;
 wire \final_adder.p_new$872 ;
 wire \final_adder.p_new$874 ;
 wire \final_adder.p_new$876 ;
 wire \final_adder.p_new$878 ;
 wire \final_adder.p_new$880 ;
 wire \final_adder.p_new$882 ;
 wire \final_adder.p_new$884 ;
 wire \final_adder.p_new$886 ;
 wire \final_adder.p_new$888 ;
 wire \final_adder.p_new$890 ;
 wire \final_adder.p_new$892 ;
 wire \final_adder.p_new$894 ;
 wire \final_adder.p_new$896 ;
 wire \final_adder.p_new$898 ;
 wire \final_adder.p_new$900 ;
 wire \final_adder.p_new$902 ;
 wire \final_adder.p_new$904 ;
 wire \final_adder.p_new$906 ;
 wire \final_adder.p_new$908 ;
 wire \final_adder.p_new$910 ;
 wire \final_adder.p_new$912 ;
 wire \final_adder.p_new$914 ;
 wire \final_adder.p_new$916 ;
 wire \final_adder.p_new$918 ;
 wire \final_adder.p_new$920 ;
 wire \final_adder.p_new$922 ;
 wire \final_adder.p_new$924 ;
 wire \final_adder.p_new$926 ;
 wire \final_adder.p_new$928 ;
 wire \notblock$4475[0] ;
 wire \notblock$4475[1] ;
 wire \notblock$4475[2] ;
 wire \notblock$4545[0] ;
 wire \notblock$4545[1] ;
 wire \notblock$4545[2] ;
 wire \notblock$4615[0] ;
 wire \notblock$4615[1] ;
 wire \notblock$4615[2] ;
 wire \notblock$4685[0] ;
 wire \notblock$4685[1] ;
 wire \notblock$4685[2] ;
 wire \notblock$4755[0] ;
 wire \notblock$4755[1] ;
 wire \notblock$4755[2] ;
 wire \notblock$4825[0] ;
 wire \notblock$4825[1] ;
 wire \notblock$4825[2] ;
 wire \notblock$4895[0] ;
 wire \notblock$4895[1] ;
 wire \notblock$4895[2] ;
 wire \notblock$4965[0] ;
 wire \notblock$4965[1] ;
 wire \notblock$4965[2] ;
 wire \notblock$5035[0] ;
 wire \notblock$5035[1] ;
 wire \notblock$5035[2] ;
 wire \notblock$5105[0] ;
 wire \notblock$5105[1] ;
 wire \notblock$5105[2] ;
 wire \notblock$5175[0] ;
 wire \notblock$5175[1] ;
 wire \notblock$5175[2] ;
 wire \notblock$5245[0] ;
 wire \notblock$5245[1] ;
 wire \notblock$5245[2] ;
 wire \notblock$5315[0] ;
 wire \notblock$5315[1] ;
 wire \notblock$5315[2] ;
 wire \notblock$5385[0] ;
 wire \notblock$5385[1] ;
 wire \notblock$5385[2] ;
 wire \notblock$5455[0] ;
 wire \notblock$5455[1] ;
 wire \notblock$5455[2] ;
 wire \notblock$5525[0] ;
 wire \notblock$5525[1] ;
 wire \notblock$5525[2] ;
 wire \notblock$5595[0] ;
 wire \notblock$5595[1] ;
 wire \notblock$5595[2] ;
 wire \notblock$5665[0] ;
 wire \notblock$5665[1] ;
 wire \notblock$5665[2] ;
 wire \notblock$5735[0] ;
 wire \notblock$5735[1] ;
 wire \notblock$5735[2] ;
 wire \notblock$5805[0] ;
 wire \notblock$5805[1] ;
 wire \notblock$5805[2] ;
 wire \notblock$5875[0] ;
 wire \notblock$5875[1] ;
 wire \notblock$5875[2] ;
 wire \notblock$5945[0] ;
 wire \notblock$5945[1] ;
 wire \notblock$5945[2] ;
 wire \notblock$6015[0] ;
 wire \notblock$6015[1] ;
 wire \notblock$6015[2] ;
 wire \notblock$6085[0] ;
 wire \notblock$6085[1] ;
 wire \notblock$6085[2] ;
 wire \notblock$6155[0] ;
 wire \notblock$6155[1] ;
 wire \notblock$6155[2] ;
 wire \notblock$6225[0] ;
 wire \notblock$6225[1] ;
 wire \notblock$6225[2] ;
 wire \notblock$6295[0] ;
 wire \notblock$6295[1] ;
 wire \notblock$6295[2] ;
 wire \notblock$6365[0] ;
 wire \notblock$6365[1] ;
 wire \notblock$6365[2] ;
 wire \notblock$6435[0] ;
 wire \notblock$6435[1] ;
 wire \notblock$6435[2] ;
 wire \notblock$6505[0] ;
 wire \notblock$6505[1] ;
 wire \notblock$6505[2] ;
 wire \notblock$6575[0] ;
 wire \notblock$6575[1] ;
 wire \notblock$6575[2] ;
 wire \notblock$6645[0] ;
 wire \notblock$6645[1] ;
 wire \notblock$6645[2] ;
 wire \notblock[0] ;
 wire \notblock[1] ;
 wire \notblock[2] ;
 wire notsign;
 wire \notsign$4544 ;
 wire \notsign$4614 ;
 wire \notsign$4684 ;
 wire \notsign$4754 ;
 wire \notsign$4824 ;
 wire \notsign$4894 ;
 wire \notsign$4964 ;
 wire \notsign$5034 ;
 wire \notsign$5104 ;
 wire \notsign$5174 ;
 wire \notsign$5244 ;
 wire \notsign$5314 ;
 wire \notsign$5384 ;
 wire \notsign$5454 ;
 wire \notsign$5524 ;
 wire \notsign$5594 ;
 wire \notsign$5664 ;
 wire \notsign$5734 ;
 wire \notsign$5804 ;
 wire \notsign$5874 ;
 wire \notsign$5944 ;
 wire \notsign$6014 ;
 wire \notsign$6084 ;
 wire \notsign$6154 ;
 wire \notsign$6224 ;
 wire \notsign$6294 ;
 wire \notsign$6364 ;
 wire \notsign$6434 ;
 wire \notsign$6504 ;
 wire \notsign$6574 ;
 wire \notsign$6644 ;
 wire pp_row0_0;
 wire pp_row0_1;
 wire pp_row0_2;
 wire pp_row100_1;
 wire pp_row100_10;
 wire pp_row100_11;
 wire pp_row100_12;
 wire pp_row100_13;
 wire pp_row100_14;
 wire pp_row100_15;
 wire pp_row100_16;
 wire pp_row100_2;
 wire pp_row100_3;
 wire pp_row100_4;
 wire pp_row100_5;
 wire pp_row100_6;
 wire pp_row100_7;
 wire pp_row100_8;
 wire pp_row100_9;
 wire pp_row101_0;
 wire pp_row101_1;
 wire pp_row101_10;
 wire pp_row101_11;
 wire pp_row101_12;
 wire pp_row101_13;
 wire pp_row101_14;
 wire pp_row101_15;
 wire pp_row101_2;
 wire pp_row101_3;
 wire pp_row101_4;
 wire pp_row101_5;
 wire pp_row101_6;
 wire pp_row101_7;
 wire pp_row101_8;
 wire pp_row101_9;
 wire pp_row102_1;
 wire pp_row102_10;
 wire pp_row102_11;
 wire pp_row102_12;
 wire pp_row102_13;
 wire pp_row102_14;
 wire pp_row102_15;
 wire pp_row102_2;
 wire pp_row102_3;
 wire pp_row102_4;
 wire pp_row102_5;
 wire pp_row102_6;
 wire pp_row102_7;
 wire pp_row102_8;
 wire pp_row102_9;
 wire pp_row103_0;
 wire pp_row103_1;
 wire pp_row103_10;
 wire pp_row103_11;
 wire pp_row103_12;
 wire pp_row103_13;
 wire pp_row103_14;
 wire pp_row103_2;
 wire pp_row103_3;
 wire pp_row103_4;
 wire pp_row103_5;
 wire pp_row103_6;
 wire pp_row103_7;
 wire pp_row103_8;
 wire pp_row103_9;
 wire pp_row104_1;
 wire pp_row104_10;
 wire pp_row104_11;
 wire pp_row104_12;
 wire pp_row104_13;
 wire pp_row104_14;
 wire pp_row104_2;
 wire pp_row104_3;
 wire pp_row104_4;
 wire pp_row104_5;
 wire pp_row104_6;
 wire pp_row104_7;
 wire pp_row104_8;
 wire pp_row104_9;
 wire pp_row105_0;
 wire pp_row105_1;
 wire pp_row105_10;
 wire pp_row105_11;
 wire pp_row105_12;
 wire pp_row105_13;
 wire pp_row105_2;
 wire pp_row105_3;
 wire pp_row105_4;
 wire pp_row105_5;
 wire pp_row105_6;
 wire pp_row105_7;
 wire pp_row105_8;
 wire pp_row105_9;
 wire pp_row106_1;
 wire pp_row106_10;
 wire pp_row106_11;
 wire pp_row106_12;
 wire pp_row106_13;
 wire pp_row106_2;
 wire pp_row106_3;
 wire pp_row106_4;
 wire pp_row106_5;
 wire pp_row106_6;
 wire pp_row106_7;
 wire pp_row106_8;
 wire pp_row106_9;
 wire pp_row107_0;
 wire pp_row107_1;
 wire pp_row107_10;
 wire pp_row107_11;
 wire pp_row107_12;
 wire pp_row107_2;
 wire pp_row107_3;
 wire pp_row107_4;
 wire pp_row107_5;
 wire pp_row107_6;
 wire pp_row107_7;
 wire pp_row107_8;
 wire pp_row107_9;
 wire pp_row108_1;
 wire pp_row108_10;
 wire pp_row108_11;
 wire pp_row108_12;
 wire pp_row108_2;
 wire pp_row108_3;
 wire pp_row108_4;
 wire pp_row108_5;
 wire pp_row108_6;
 wire pp_row108_7;
 wire pp_row108_8;
 wire pp_row108_9;
 wire pp_row109_0;
 wire pp_row109_1;
 wire pp_row109_10;
 wire pp_row109_11;
 wire pp_row109_2;
 wire pp_row109_3;
 wire pp_row109_4;
 wire pp_row109_5;
 wire pp_row109_6;
 wire pp_row109_7;
 wire pp_row109_8;
 wire pp_row109_9;
 wire pp_row10_0;
 wire pp_row10_1;
 wire pp_row10_2;
 wire pp_row10_3;
 wire pp_row10_4;
 wire pp_row10_5;
 wire pp_row10_6;
 wire pp_row10_7;
 wire pp_row110_1;
 wire pp_row110_10;
 wire pp_row110_11;
 wire pp_row110_2;
 wire pp_row110_3;
 wire pp_row110_4;
 wire pp_row110_5;
 wire pp_row110_6;
 wire pp_row110_7;
 wire pp_row110_8;
 wire pp_row110_9;
 wire pp_row111_0;
 wire pp_row111_1;
 wire pp_row111_10;
 wire pp_row111_2;
 wire pp_row111_3;
 wire pp_row111_4;
 wire pp_row111_5;
 wire pp_row111_6;
 wire pp_row111_7;
 wire pp_row111_8;
 wire pp_row111_9;
 wire pp_row112_1;
 wire pp_row112_10;
 wire pp_row112_2;
 wire pp_row112_3;
 wire pp_row112_4;
 wire pp_row112_5;
 wire pp_row112_6;
 wire pp_row112_7;
 wire pp_row112_8;
 wire pp_row112_9;
 wire pp_row113_0;
 wire pp_row113_1;
 wire pp_row113_2;
 wire pp_row113_3;
 wire pp_row113_4;
 wire pp_row113_5;
 wire pp_row113_6;
 wire pp_row113_7;
 wire pp_row113_8;
 wire pp_row113_9;
 wire pp_row114_1;
 wire pp_row114_2;
 wire pp_row114_3;
 wire pp_row114_4;
 wire pp_row114_5;
 wire pp_row114_6;
 wire pp_row114_7;
 wire pp_row114_8;
 wire pp_row114_9;
 wire pp_row115_0;
 wire pp_row115_1;
 wire pp_row115_2;
 wire pp_row115_3;
 wire pp_row115_4;
 wire pp_row115_5;
 wire pp_row115_6;
 wire pp_row115_7;
 wire pp_row115_8;
 wire pp_row116_1;
 wire pp_row116_2;
 wire pp_row116_3;
 wire pp_row116_4;
 wire pp_row116_5;
 wire pp_row116_6;
 wire pp_row116_7;
 wire pp_row116_8;
 wire pp_row117_0;
 wire pp_row117_1;
 wire pp_row117_2;
 wire pp_row117_3;
 wire pp_row117_4;
 wire pp_row117_5;
 wire pp_row117_6;
 wire pp_row117_7;
 wire pp_row118_1;
 wire pp_row118_2;
 wire pp_row118_3;
 wire pp_row118_4;
 wire pp_row118_5;
 wire pp_row118_6;
 wire pp_row118_7;
 wire pp_row119_0;
 wire pp_row119_1;
 wire pp_row119_2;
 wire pp_row119_3;
 wire pp_row119_4;
 wire pp_row119_5;
 wire pp_row119_6;
 wire pp_row11_0;
 wire pp_row11_1;
 wire pp_row11_2;
 wire pp_row11_3;
 wire pp_row11_4;
 wire pp_row11_5;
 wire pp_row11_6;
 wire pp_row120_1;
 wire pp_row120_2;
 wire pp_row120_3;
 wire pp_row120_4;
 wire pp_row120_5;
 wire pp_row120_6;
 wire pp_row121_0;
 wire pp_row121_1;
 wire pp_row121_2;
 wire pp_row121_3;
 wire pp_row121_4;
 wire pp_row121_5;
 wire pp_row122_1;
 wire pp_row122_2;
 wire pp_row122_3;
 wire pp_row122_4;
 wire pp_row122_5;
 wire pp_row123_0;
 wire pp_row123_1;
 wire pp_row123_2;
 wire pp_row123_3;
 wire pp_row123_4;
 wire pp_row124_1;
 wire pp_row124_2;
 wire pp_row124_3;
 wire pp_row124_4;
 wire pp_row125_0;
 wire pp_row125_1;
 wire pp_row125_2;
 wire pp_row125_3;
 wire pp_row126_1;
 wire pp_row126_2;
 wire pp_row126_3;
 wire pp_row127_0;
 wire pp_row127_1;
 wire pp_row127_2;
 wire pp_row12_0;
 wire pp_row12_1;
 wire pp_row12_2;
 wire pp_row12_3;
 wire pp_row12_4;
 wire pp_row12_5;
 wire pp_row12_6;
 wire pp_row12_7;
 wire pp_row12_8;
 wire pp_row13_0;
 wire pp_row13_1;
 wire pp_row13_2;
 wire pp_row13_3;
 wire pp_row13_4;
 wire pp_row13_5;
 wire pp_row13_6;
 wire pp_row13_7;
 wire pp_row14_0;
 wire pp_row14_1;
 wire pp_row14_2;
 wire pp_row14_3;
 wire pp_row14_4;
 wire pp_row14_5;
 wire pp_row14_6;
 wire pp_row14_7;
 wire pp_row14_8;
 wire pp_row14_9;
 wire pp_row15_0;
 wire pp_row15_1;
 wire pp_row15_2;
 wire pp_row15_3;
 wire pp_row15_4;
 wire pp_row15_5;
 wire pp_row15_6;
 wire pp_row15_7;
 wire pp_row15_8;
 wire pp_row16_0;
 wire pp_row16_1;
 wire pp_row16_10;
 wire pp_row16_2;
 wire pp_row16_3;
 wire pp_row16_4;
 wire pp_row16_5;
 wire pp_row16_6;
 wire pp_row16_7;
 wire pp_row16_8;
 wire pp_row16_9;
 wire pp_row17_0;
 wire pp_row17_1;
 wire pp_row17_2;
 wire pp_row17_3;
 wire pp_row17_4;
 wire pp_row17_5;
 wire pp_row17_6;
 wire pp_row17_7;
 wire pp_row17_8;
 wire pp_row17_9;
 wire pp_row18_0;
 wire pp_row18_1;
 wire pp_row18_10;
 wire pp_row18_11;
 wire pp_row18_2;
 wire pp_row18_3;
 wire pp_row18_4;
 wire pp_row18_5;
 wire pp_row18_6;
 wire pp_row18_7;
 wire pp_row18_8;
 wire pp_row18_9;
 wire pp_row19_0;
 wire pp_row19_1;
 wire pp_row19_10;
 wire pp_row19_2;
 wire pp_row19_3;
 wire pp_row19_4;
 wire pp_row19_5;
 wire pp_row19_6;
 wire pp_row19_7;
 wire pp_row19_8;
 wire pp_row19_9;
 wire pp_row1_0;
 wire pp_row1_1;
 wire pp_row20_0;
 wire pp_row20_1;
 wire pp_row20_10;
 wire pp_row20_11;
 wire pp_row20_12;
 wire pp_row20_2;
 wire pp_row20_3;
 wire pp_row20_4;
 wire pp_row20_5;
 wire pp_row20_6;
 wire pp_row20_7;
 wire pp_row20_8;
 wire pp_row20_9;
 wire pp_row21_0;
 wire pp_row21_1;
 wire pp_row21_10;
 wire pp_row21_11;
 wire pp_row21_2;
 wire pp_row21_3;
 wire pp_row21_4;
 wire pp_row21_5;
 wire pp_row21_6;
 wire pp_row21_7;
 wire pp_row21_8;
 wire pp_row21_9;
 wire pp_row22_0;
 wire pp_row22_1;
 wire pp_row22_10;
 wire pp_row22_11;
 wire pp_row22_12;
 wire pp_row22_13;
 wire pp_row22_2;
 wire pp_row22_3;
 wire pp_row22_4;
 wire pp_row22_5;
 wire pp_row22_6;
 wire pp_row22_7;
 wire pp_row22_8;
 wire pp_row22_9;
 wire pp_row23_0;
 wire pp_row23_1;
 wire pp_row23_10;
 wire pp_row23_11;
 wire pp_row23_12;
 wire pp_row23_2;
 wire pp_row23_3;
 wire pp_row23_4;
 wire pp_row23_5;
 wire pp_row23_6;
 wire pp_row23_7;
 wire pp_row23_8;
 wire pp_row23_9;
 wire pp_row24_0;
 wire pp_row24_1;
 wire pp_row24_10;
 wire pp_row24_11;
 wire pp_row24_12;
 wire pp_row24_13;
 wire pp_row24_14;
 wire pp_row24_2;
 wire pp_row24_3;
 wire pp_row24_4;
 wire pp_row24_5;
 wire pp_row24_6;
 wire pp_row24_7;
 wire pp_row24_8;
 wire pp_row24_9;
 wire pp_row25_0;
 wire pp_row25_1;
 wire pp_row25_10;
 wire pp_row25_11;
 wire pp_row25_12;
 wire pp_row25_13;
 wire pp_row25_2;
 wire pp_row25_3;
 wire pp_row25_4;
 wire pp_row25_5;
 wire pp_row25_6;
 wire pp_row25_7;
 wire pp_row25_8;
 wire pp_row25_9;
 wire pp_row26_0;
 wire pp_row26_1;
 wire pp_row26_10;
 wire pp_row26_11;
 wire pp_row26_12;
 wire pp_row26_13;
 wire pp_row26_14;
 wire pp_row26_15;
 wire pp_row26_2;
 wire pp_row26_3;
 wire pp_row26_4;
 wire pp_row26_5;
 wire pp_row26_6;
 wire pp_row26_7;
 wire pp_row26_8;
 wire pp_row26_9;
 wire pp_row27_0;
 wire pp_row27_1;
 wire pp_row27_10;
 wire pp_row27_11;
 wire pp_row27_12;
 wire pp_row27_13;
 wire pp_row27_14;
 wire pp_row27_2;
 wire pp_row27_3;
 wire pp_row27_4;
 wire pp_row27_5;
 wire pp_row27_6;
 wire pp_row27_7;
 wire pp_row27_8;
 wire pp_row27_9;
 wire pp_row28_0;
 wire pp_row28_1;
 wire pp_row28_10;
 wire pp_row28_11;
 wire pp_row28_12;
 wire pp_row28_13;
 wire pp_row28_14;
 wire pp_row28_15;
 wire pp_row28_16;
 wire pp_row28_2;
 wire pp_row28_3;
 wire pp_row28_4;
 wire pp_row28_5;
 wire pp_row28_6;
 wire pp_row28_7;
 wire pp_row28_8;
 wire pp_row28_9;
 wire pp_row29_0;
 wire pp_row29_1;
 wire pp_row29_10;
 wire pp_row29_11;
 wire pp_row29_12;
 wire pp_row29_13;
 wire pp_row29_14;
 wire pp_row29_15;
 wire pp_row29_2;
 wire pp_row29_3;
 wire pp_row29_4;
 wire pp_row29_5;
 wire pp_row29_6;
 wire pp_row29_7;
 wire pp_row29_8;
 wire pp_row29_9;
 wire pp_row2_0;
 wire pp_row2_1;
 wire pp_row2_2;
 wire pp_row2_3;
 wire pp_row30_0;
 wire pp_row30_1;
 wire pp_row30_10;
 wire pp_row30_11;
 wire pp_row30_12;
 wire pp_row30_13;
 wire pp_row30_14;
 wire pp_row30_15;
 wire pp_row30_16;
 wire pp_row30_17;
 wire pp_row30_2;
 wire pp_row30_3;
 wire pp_row30_4;
 wire pp_row30_5;
 wire pp_row30_6;
 wire pp_row30_7;
 wire pp_row30_8;
 wire pp_row30_9;
 wire pp_row31_0;
 wire pp_row31_1;
 wire pp_row31_10;
 wire pp_row31_11;
 wire pp_row31_12;
 wire pp_row31_13;
 wire pp_row31_14;
 wire pp_row31_15;
 wire pp_row31_16;
 wire pp_row31_2;
 wire pp_row31_3;
 wire pp_row31_4;
 wire pp_row31_5;
 wire pp_row31_6;
 wire pp_row31_7;
 wire pp_row31_8;
 wire pp_row31_9;
 wire pp_row32_0;
 wire pp_row32_1;
 wire pp_row32_10;
 wire pp_row32_11;
 wire pp_row32_12;
 wire pp_row32_13;
 wire pp_row32_14;
 wire pp_row32_15;
 wire pp_row32_16;
 wire pp_row32_17;
 wire pp_row32_18;
 wire pp_row32_2;
 wire pp_row32_3;
 wire pp_row32_4;
 wire pp_row32_5;
 wire pp_row32_6;
 wire pp_row32_7;
 wire pp_row32_8;
 wire pp_row32_9;
 wire pp_row33_0;
 wire pp_row33_1;
 wire pp_row33_10;
 wire pp_row33_11;
 wire pp_row33_12;
 wire pp_row33_13;
 wire pp_row33_14;
 wire pp_row33_15;
 wire pp_row33_16;
 wire pp_row33_17;
 wire pp_row33_2;
 wire pp_row33_3;
 wire pp_row33_4;
 wire pp_row33_5;
 wire pp_row33_6;
 wire pp_row33_7;
 wire pp_row33_8;
 wire pp_row33_9;
 wire pp_row34_0;
 wire pp_row34_1;
 wire pp_row34_10;
 wire pp_row34_11;
 wire pp_row34_12;
 wire pp_row34_13;
 wire pp_row34_14;
 wire pp_row34_15;
 wire pp_row34_16;
 wire pp_row34_17;
 wire pp_row34_18;
 wire pp_row34_19;
 wire pp_row34_2;
 wire pp_row34_3;
 wire pp_row34_4;
 wire pp_row34_5;
 wire pp_row34_6;
 wire pp_row34_7;
 wire pp_row34_8;
 wire pp_row34_9;
 wire pp_row35_0;
 wire pp_row35_1;
 wire pp_row35_10;
 wire pp_row35_11;
 wire pp_row35_12;
 wire pp_row35_13;
 wire pp_row35_14;
 wire pp_row35_15;
 wire pp_row35_16;
 wire pp_row35_17;
 wire pp_row35_18;
 wire pp_row35_2;
 wire pp_row35_3;
 wire pp_row35_4;
 wire pp_row35_5;
 wire pp_row35_6;
 wire pp_row35_7;
 wire pp_row35_8;
 wire pp_row35_9;
 wire pp_row36_0;
 wire pp_row36_1;
 wire pp_row36_10;
 wire pp_row36_11;
 wire pp_row36_12;
 wire pp_row36_13;
 wire pp_row36_14;
 wire pp_row36_15;
 wire pp_row36_16;
 wire pp_row36_17;
 wire pp_row36_18;
 wire pp_row36_19;
 wire pp_row36_2;
 wire pp_row36_20;
 wire pp_row36_3;
 wire pp_row36_4;
 wire pp_row36_5;
 wire pp_row36_6;
 wire pp_row36_7;
 wire pp_row36_8;
 wire pp_row36_9;
 wire pp_row37_0;
 wire pp_row37_1;
 wire pp_row37_10;
 wire pp_row37_11;
 wire pp_row37_12;
 wire pp_row37_13;
 wire pp_row37_14;
 wire pp_row37_15;
 wire pp_row37_16;
 wire pp_row37_17;
 wire pp_row37_18;
 wire pp_row37_19;
 wire pp_row37_2;
 wire pp_row37_3;
 wire pp_row37_4;
 wire pp_row37_5;
 wire pp_row37_6;
 wire pp_row37_7;
 wire pp_row37_8;
 wire pp_row37_9;
 wire pp_row38_0;
 wire pp_row38_1;
 wire pp_row38_10;
 wire pp_row38_11;
 wire pp_row38_12;
 wire pp_row38_13;
 wire pp_row38_14;
 wire pp_row38_15;
 wire pp_row38_16;
 wire pp_row38_17;
 wire pp_row38_18;
 wire pp_row38_19;
 wire pp_row38_2;
 wire pp_row38_20;
 wire pp_row38_21;
 wire pp_row38_3;
 wire pp_row38_4;
 wire pp_row38_5;
 wire pp_row38_6;
 wire pp_row38_7;
 wire pp_row38_8;
 wire pp_row38_9;
 wire pp_row39_0;
 wire pp_row39_1;
 wire pp_row39_10;
 wire pp_row39_11;
 wire pp_row39_12;
 wire pp_row39_13;
 wire pp_row39_14;
 wire pp_row39_15;
 wire pp_row39_16;
 wire pp_row39_17;
 wire pp_row39_18;
 wire pp_row39_19;
 wire pp_row39_2;
 wire pp_row39_20;
 wire pp_row39_3;
 wire pp_row39_4;
 wire pp_row39_5;
 wire pp_row39_6;
 wire pp_row39_7;
 wire pp_row39_8;
 wire pp_row39_9;
 wire pp_row3_0;
 wire pp_row3_1;
 wire pp_row3_2;
 wire pp_row40_0;
 wire pp_row40_1;
 wire pp_row40_10;
 wire pp_row40_11;
 wire pp_row40_12;
 wire pp_row40_13;
 wire pp_row40_14;
 wire pp_row40_15;
 wire pp_row40_16;
 wire pp_row40_17;
 wire pp_row40_18;
 wire pp_row40_19;
 wire pp_row40_2;
 wire pp_row40_20;
 wire pp_row40_21;
 wire pp_row40_22;
 wire pp_row40_3;
 wire pp_row40_4;
 wire pp_row40_5;
 wire pp_row40_6;
 wire pp_row40_7;
 wire pp_row40_8;
 wire pp_row40_9;
 wire pp_row41_0;
 wire pp_row41_1;
 wire pp_row41_10;
 wire pp_row41_11;
 wire pp_row41_12;
 wire pp_row41_13;
 wire pp_row41_14;
 wire pp_row41_15;
 wire pp_row41_16;
 wire pp_row41_17;
 wire pp_row41_18;
 wire pp_row41_19;
 wire pp_row41_2;
 wire pp_row41_20;
 wire pp_row41_21;
 wire pp_row41_3;
 wire pp_row41_4;
 wire pp_row41_5;
 wire pp_row41_6;
 wire pp_row41_7;
 wire pp_row41_8;
 wire pp_row41_9;
 wire pp_row42_0;
 wire pp_row42_1;
 wire pp_row42_10;
 wire pp_row42_11;
 wire pp_row42_12;
 wire pp_row42_13;
 wire pp_row42_14;
 wire pp_row42_15;
 wire pp_row42_16;
 wire pp_row42_17;
 wire pp_row42_18;
 wire pp_row42_19;
 wire pp_row42_2;
 wire pp_row42_20;
 wire pp_row42_21;
 wire pp_row42_22;
 wire pp_row42_23;
 wire pp_row42_3;
 wire pp_row42_4;
 wire pp_row42_5;
 wire pp_row42_6;
 wire pp_row42_7;
 wire pp_row42_8;
 wire pp_row42_9;
 wire pp_row43_0;
 wire pp_row43_1;
 wire pp_row43_10;
 wire pp_row43_11;
 wire pp_row43_12;
 wire pp_row43_13;
 wire pp_row43_14;
 wire pp_row43_15;
 wire pp_row43_16;
 wire pp_row43_17;
 wire pp_row43_18;
 wire pp_row43_19;
 wire pp_row43_2;
 wire pp_row43_20;
 wire pp_row43_21;
 wire pp_row43_22;
 wire pp_row43_3;
 wire pp_row43_4;
 wire pp_row43_5;
 wire pp_row43_6;
 wire pp_row43_7;
 wire pp_row43_8;
 wire pp_row43_9;
 wire pp_row44_0;
 wire pp_row44_1;
 wire pp_row44_10;
 wire pp_row44_11;
 wire pp_row44_12;
 wire pp_row44_13;
 wire pp_row44_14;
 wire pp_row44_15;
 wire pp_row44_16;
 wire pp_row44_17;
 wire pp_row44_18;
 wire pp_row44_19;
 wire pp_row44_2;
 wire pp_row44_20;
 wire pp_row44_21;
 wire pp_row44_22;
 wire pp_row44_23;
 wire pp_row44_24;
 wire pp_row44_3;
 wire pp_row44_4;
 wire pp_row44_5;
 wire pp_row44_6;
 wire pp_row44_7;
 wire pp_row44_8;
 wire pp_row44_9;
 wire pp_row45_0;
 wire pp_row45_1;
 wire pp_row45_10;
 wire pp_row45_11;
 wire pp_row45_12;
 wire pp_row45_13;
 wire pp_row45_14;
 wire pp_row45_15;
 wire pp_row45_16;
 wire pp_row45_17;
 wire pp_row45_18;
 wire pp_row45_19;
 wire pp_row45_2;
 wire pp_row45_20;
 wire pp_row45_21;
 wire pp_row45_22;
 wire pp_row45_23;
 wire pp_row45_3;
 wire pp_row45_4;
 wire pp_row45_5;
 wire pp_row45_6;
 wire pp_row45_7;
 wire pp_row45_8;
 wire pp_row45_9;
 wire pp_row46_0;
 wire pp_row46_1;
 wire pp_row46_10;
 wire pp_row46_11;
 wire pp_row46_12;
 wire pp_row46_13;
 wire pp_row46_14;
 wire pp_row46_15;
 wire pp_row46_16;
 wire pp_row46_17;
 wire pp_row46_18;
 wire pp_row46_19;
 wire pp_row46_2;
 wire pp_row46_20;
 wire pp_row46_21;
 wire pp_row46_22;
 wire pp_row46_23;
 wire pp_row46_24;
 wire pp_row46_25;
 wire pp_row46_3;
 wire pp_row46_4;
 wire pp_row46_5;
 wire pp_row46_6;
 wire pp_row46_7;
 wire pp_row46_8;
 wire pp_row46_9;
 wire pp_row47_0;
 wire pp_row47_1;
 wire pp_row47_10;
 wire pp_row47_11;
 wire pp_row47_12;
 wire pp_row47_13;
 wire pp_row47_14;
 wire pp_row47_15;
 wire pp_row47_16;
 wire pp_row47_17;
 wire pp_row47_18;
 wire pp_row47_19;
 wire pp_row47_2;
 wire pp_row47_20;
 wire pp_row47_21;
 wire pp_row47_22;
 wire pp_row47_23;
 wire pp_row47_24;
 wire pp_row47_3;
 wire pp_row47_4;
 wire pp_row47_5;
 wire pp_row47_6;
 wire pp_row47_7;
 wire pp_row47_8;
 wire pp_row47_9;
 wire pp_row48_0;
 wire pp_row48_1;
 wire pp_row48_10;
 wire pp_row48_11;
 wire pp_row48_12;
 wire pp_row48_13;
 wire pp_row48_14;
 wire pp_row48_15;
 wire pp_row48_16;
 wire pp_row48_17;
 wire pp_row48_18;
 wire pp_row48_19;
 wire pp_row48_2;
 wire pp_row48_20;
 wire pp_row48_21;
 wire pp_row48_22;
 wire pp_row48_23;
 wire pp_row48_24;
 wire pp_row48_25;
 wire pp_row48_26;
 wire pp_row48_3;
 wire pp_row48_4;
 wire pp_row48_5;
 wire pp_row48_6;
 wire pp_row48_7;
 wire pp_row48_8;
 wire pp_row48_9;
 wire pp_row49_0;
 wire pp_row49_1;
 wire pp_row49_10;
 wire pp_row49_11;
 wire pp_row49_12;
 wire pp_row49_13;
 wire pp_row49_14;
 wire pp_row49_15;
 wire pp_row49_16;
 wire pp_row49_17;
 wire pp_row49_18;
 wire pp_row49_19;
 wire pp_row49_2;
 wire pp_row49_20;
 wire pp_row49_21;
 wire pp_row49_22;
 wire pp_row49_23;
 wire pp_row49_24;
 wire pp_row49_25;
 wire pp_row49_3;
 wire pp_row49_4;
 wire pp_row49_5;
 wire pp_row49_6;
 wire pp_row49_7;
 wire pp_row49_8;
 wire pp_row49_9;
 wire pp_row4_0;
 wire pp_row4_1;
 wire pp_row4_2;
 wire pp_row4_3;
 wire pp_row4_4;
 wire pp_row50_0;
 wire pp_row50_1;
 wire pp_row50_10;
 wire pp_row50_11;
 wire pp_row50_12;
 wire pp_row50_13;
 wire pp_row50_14;
 wire pp_row50_15;
 wire pp_row50_16;
 wire pp_row50_17;
 wire pp_row50_18;
 wire pp_row50_19;
 wire pp_row50_2;
 wire pp_row50_20;
 wire pp_row50_21;
 wire pp_row50_22;
 wire pp_row50_23;
 wire pp_row50_24;
 wire pp_row50_25;
 wire pp_row50_26;
 wire pp_row50_27;
 wire pp_row50_3;
 wire pp_row50_4;
 wire pp_row50_5;
 wire pp_row50_6;
 wire pp_row50_7;
 wire pp_row50_8;
 wire pp_row50_9;
 wire pp_row51_0;
 wire pp_row51_1;
 wire pp_row51_10;
 wire pp_row51_11;
 wire pp_row51_12;
 wire pp_row51_13;
 wire pp_row51_14;
 wire pp_row51_15;
 wire pp_row51_16;
 wire pp_row51_17;
 wire pp_row51_18;
 wire pp_row51_19;
 wire pp_row51_2;
 wire pp_row51_20;
 wire pp_row51_21;
 wire pp_row51_22;
 wire pp_row51_23;
 wire pp_row51_24;
 wire pp_row51_25;
 wire pp_row51_26;
 wire pp_row51_3;
 wire pp_row51_4;
 wire pp_row51_5;
 wire pp_row51_6;
 wire pp_row51_7;
 wire pp_row51_8;
 wire pp_row51_9;
 wire pp_row52_0;
 wire pp_row52_1;
 wire pp_row52_10;
 wire pp_row52_11;
 wire pp_row52_12;
 wire pp_row52_13;
 wire pp_row52_14;
 wire pp_row52_15;
 wire pp_row52_16;
 wire pp_row52_17;
 wire pp_row52_18;
 wire pp_row52_19;
 wire pp_row52_2;
 wire pp_row52_20;
 wire pp_row52_21;
 wire pp_row52_22;
 wire pp_row52_23;
 wire pp_row52_24;
 wire pp_row52_25;
 wire pp_row52_26;
 wire pp_row52_27;
 wire pp_row52_28;
 wire pp_row52_3;
 wire pp_row52_4;
 wire pp_row52_5;
 wire pp_row52_6;
 wire pp_row52_7;
 wire pp_row52_8;
 wire pp_row52_9;
 wire pp_row53_0;
 wire pp_row53_1;
 wire pp_row53_10;
 wire pp_row53_11;
 wire pp_row53_12;
 wire pp_row53_13;
 wire pp_row53_14;
 wire pp_row53_15;
 wire pp_row53_16;
 wire pp_row53_17;
 wire pp_row53_18;
 wire pp_row53_19;
 wire pp_row53_2;
 wire pp_row53_20;
 wire pp_row53_21;
 wire pp_row53_22;
 wire pp_row53_23;
 wire pp_row53_24;
 wire pp_row53_25;
 wire pp_row53_26;
 wire pp_row53_27;
 wire pp_row53_3;
 wire pp_row53_4;
 wire pp_row53_5;
 wire pp_row53_6;
 wire pp_row53_7;
 wire pp_row53_8;
 wire pp_row53_9;
 wire pp_row54_0;
 wire pp_row54_1;
 wire pp_row54_10;
 wire pp_row54_11;
 wire pp_row54_12;
 wire pp_row54_13;
 wire pp_row54_14;
 wire pp_row54_15;
 wire pp_row54_16;
 wire pp_row54_17;
 wire pp_row54_18;
 wire pp_row54_19;
 wire pp_row54_2;
 wire pp_row54_20;
 wire pp_row54_21;
 wire pp_row54_22;
 wire pp_row54_23;
 wire pp_row54_24;
 wire pp_row54_25;
 wire pp_row54_26;
 wire pp_row54_27;
 wire pp_row54_28;
 wire pp_row54_29;
 wire pp_row54_3;
 wire pp_row54_4;
 wire pp_row54_5;
 wire pp_row54_6;
 wire pp_row54_7;
 wire pp_row54_8;
 wire pp_row54_9;
 wire pp_row55_0;
 wire pp_row55_1;
 wire pp_row55_10;
 wire pp_row55_11;
 wire pp_row55_12;
 wire pp_row55_13;
 wire pp_row55_14;
 wire pp_row55_15;
 wire pp_row55_16;
 wire pp_row55_17;
 wire pp_row55_18;
 wire pp_row55_19;
 wire pp_row55_2;
 wire pp_row55_20;
 wire pp_row55_21;
 wire pp_row55_22;
 wire pp_row55_23;
 wire pp_row55_24;
 wire pp_row55_25;
 wire pp_row55_26;
 wire pp_row55_27;
 wire pp_row55_28;
 wire pp_row55_3;
 wire pp_row55_4;
 wire pp_row55_5;
 wire pp_row55_6;
 wire pp_row55_7;
 wire pp_row55_8;
 wire pp_row55_9;
 wire pp_row56_0;
 wire pp_row56_1;
 wire pp_row56_10;
 wire pp_row56_11;
 wire pp_row56_12;
 wire pp_row56_13;
 wire pp_row56_14;
 wire pp_row56_15;
 wire pp_row56_16;
 wire pp_row56_17;
 wire pp_row56_18;
 wire pp_row56_19;
 wire pp_row56_2;
 wire pp_row56_20;
 wire pp_row56_21;
 wire pp_row56_22;
 wire pp_row56_23;
 wire pp_row56_24;
 wire pp_row56_25;
 wire pp_row56_26;
 wire pp_row56_27;
 wire pp_row56_28;
 wire pp_row56_29;
 wire pp_row56_3;
 wire pp_row56_30;
 wire pp_row56_4;
 wire pp_row56_5;
 wire pp_row56_6;
 wire pp_row56_7;
 wire pp_row56_8;
 wire pp_row56_9;
 wire pp_row57_0;
 wire pp_row57_1;
 wire pp_row57_10;
 wire pp_row57_11;
 wire pp_row57_12;
 wire pp_row57_13;
 wire pp_row57_14;
 wire pp_row57_15;
 wire pp_row57_16;
 wire pp_row57_17;
 wire pp_row57_18;
 wire pp_row57_19;
 wire pp_row57_2;
 wire pp_row57_20;
 wire pp_row57_21;
 wire pp_row57_22;
 wire pp_row57_23;
 wire pp_row57_24;
 wire pp_row57_25;
 wire pp_row57_26;
 wire pp_row57_27;
 wire pp_row57_28;
 wire pp_row57_29;
 wire pp_row57_3;
 wire pp_row57_4;
 wire pp_row57_5;
 wire pp_row57_6;
 wire pp_row57_7;
 wire pp_row57_8;
 wire pp_row57_9;
 wire pp_row58_0;
 wire pp_row58_1;
 wire pp_row58_10;
 wire pp_row58_11;
 wire pp_row58_12;
 wire pp_row58_13;
 wire pp_row58_14;
 wire pp_row58_15;
 wire pp_row58_16;
 wire pp_row58_17;
 wire pp_row58_18;
 wire pp_row58_19;
 wire pp_row58_2;
 wire pp_row58_20;
 wire pp_row58_21;
 wire pp_row58_22;
 wire pp_row58_23;
 wire pp_row58_24;
 wire pp_row58_25;
 wire pp_row58_26;
 wire pp_row58_27;
 wire pp_row58_28;
 wire pp_row58_29;
 wire pp_row58_3;
 wire pp_row58_30;
 wire pp_row58_31;
 wire pp_row58_4;
 wire pp_row58_5;
 wire pp_row58_6;
 wire pp_row58_7;
 wire pp_row58_8;
 wire pp_row58_9;
 wire pp_row59_0;
 wire pp_row59_1;
 wire pp_row59_10;
 wire pp_row59_11;
 wire pp_row59_12;
 wire pp_row59_13;
 wire pp_row59_14;
 wire pp_row59_15;
 wire pp_row59_16;
 wire pp_row59_17;
 wire pp_row59_18;
 wire pp_row59_19;
 wire pp_row59_2;
 wire pp_row59_20;
 wire pp_row59_21;
 wire pp_row59_22;
 wire pp_row59_23;
 wire pp_row59_24;
 wire pp_row59_25;
 wire pp_row59_26;
 wire pp_row59_27;
 wire pp_row59_28;
 wire pp_row59_29;
 wire pp_row59_3;
 wire pp_row59_30;
 wire pp_row59_4;
 wire pp_row59_5;
 wire pp_row59_6;
 wire pp_row59_7;
 wire pp_row59_8;
 wire pp_row59_9;
 wire pp_row5_0;
 wire pp_row5_1;
 wire pp_row5_2;
 wire pp_row5_3;
 wire pp_row60_0;
 wire pp_row60_1;
 wire pp_row60_10;
 wire pp_row60_11;
 wire pp_row60_12;
 wire pp_row60_13;
 wire pp_row60_14;
 wire pp_row60_15;
 wire pp_row60_16;
 wire pp_row60_17;
 wire pp_row60_18;
 wire pp_row60_19;
 wire pp_row60_2;
 wire pp_row60_20;
 wire pp_row60_21;
 wire pp_row60_22;
 wire pp_row60_23;
 wire pp_row60_24;
 wire pp_row60_25;
 wire pp_row60_26;
 wire pp_row60_27;
 wire pp_row60_28;
 wire pp_row60_29;
 wire pp_row60_3;
 wire pp_row60_30;
 wire pp_row60_31;
 wire pp_row60_32;
 wire pp_row60_4;
 wire pp_row60_5;
 wire pp_row60_6;
 wire pp_row60_7;
 wire pp_row60_8;
 wire pp_row60_9;
 wire pp_row61_0;
 wire pp_row61_1;
 wire pp_row61_10;
 wire pp_row61_11;
 wire pp_row61_12;
 wire pp_row61_13;
 wire pp_row61_14;
 wire pp_row61_15;
 wire pp_row61_16;
 wire pp_row61_17;
 wire pp_row61_18;
 wire pp_row61_19;
 wire pp_row61_2;
 wire pp_row61_20;
 wire pp_row61_21;
 wire pp_row61_22;
 wire pp_row61_23;
 wire pp_row61_24;
 wire pp_row61_25;
 wire pp_row61_26;
 wire pp_row61_27;
 wire pp_row61_28;
 wire pp_row61_29;
 wire pp_row61_3;
 wire pp_row61_30;
 wire pp_row61_31;
 wire pp_row61_4;
 wire pp_row61_5;
 wire pp_row61_6;
 wire pp_row61_7;
 wire pp_row61_8;
 wire pp_row61_9;
 wire pp_row62_0;
 wire pp_row62_1;
 wire pp_row62_10;
 wire pp_row62_11;
 wire pp_row62_12;
 wire pp_row62_13;
 wire pp_row62_14;
 wire pp_row62_15;
 wire pp_row62_16;
 wire pp_row62_17;
 wire pp_row62_18;
 wire pp_row62_19;
 wire pp_row62_2;
 wire pp_row62_20;
 wire pp_row62_21;
 wire pp_row62_22;
 wire pp_row62_23;
 wire pp_row62_24;
 wire pp_row62_25;
 wire pp_row62_26;
 wire pp_row62_27;
 wire pp_row62_28;
 wire pp_row62_29;
 wire pp_row62_3;
 wire pp_row62_30;
 wire pp_row62_31;
 wire pp_row62_32;
 wire pp_row62_33;
 wire pp_row62_4;
 wire pp_row62_5;
 wire pp_row62_6;
 wire pp_row62_7;
 wire pp_row62_8;
 wire pp_row62_9;
 wire pp_row63_0;
 wire pp_row63_1;
 wire pp_row63_10;
 wire pp_row63_11;
 wire pp_row63_12;
 wire pp_row63_13;
 wire pp_row63_14;
 wire pp_row63_15;
 wire pp_row63_16;
 wire pp_row63_17;
 wire pp_row63_18;
 wire pp_row63_19;
 wire pp_row63_2;
 wire pp_row63_20;
 wire pp_row63_21;
 wire pp_row63_22;
 wire pp_row63_23;
 wire pp_row63_24;
 wire pp_row63_25;
 wire pp_row63_26;
 wire pp_row63_27;
 wire pp_row63_28;
 wire pp_row63_29;
 wire pp_row63_3;
 wire pp_row63_30;
 wire pp_row63_31;
 wire pp_row63_32;
 wire pp_row63_4;
 wire pp_row63_5;
 wire pp_row63_6;
 wire pp_row63_7;
 wire pp_row63_8;
 wire pp_row63_9;
 wire pp_row64_0;
 wire pp_row64_1;
 wire pp_row64_10;
 wire pp_row64_11;
 wire pp_row64_12;
 wire pp_row64_13;
 wire pp_row64_14;
 wire pp_row64_15;
 wire pp_row64_16;
 wire pp_row64_17;
 wire pp_row64_18;
 wire pp_row64_19;
 wire pp_row64_2;
 wire pp_row64_20;
 wire pp_row64_21;
 wire pp_row64_22;
 wire pp_row64_23;
 wire pp_row64_24;
 wire pp_row64_25;
 wire pp_row64_26;
 wire pp_row64_27;
 wire pp_row64_28;
 wire pp_row64_29;
 wire pp_row64_3;
 wire pp_row64_30;
 wire pp_row64_31;
 wire pp_row64_32;
 wire pp_row64_33;
 wire pp_row64_4;
 wire pp_row64_5;
 wire pp_row64_6;
 wire pp_row64_7;
 wire pp_row64_8;
 wire pp_row64_9;
 wire pp_row65_1;
 wire pp_row65_10;
 wire pp_row65_11;
 wire pp_row65_12;
 wire pp_row65_13;
 wire pp_row65_14;
 wire pp_row65_15;
 wire pp_row65_16;
 wire pp_row65_17;
 wire pp_row65_18;
 wire pp_row65_19;
 wire pp_row65_2;
 wire pp_row65_20;
 wire pp_row65_21;
 wire pp_row65_22;
 wire pp_row65_23;
 wire pp_row65_24;
 wire pp_row65_25;
 wire pp_row65_26;
 wire pp_row65_27;
 wire pp_row65_28;
 wire pp_row65_29;
 wire pp_row65_3;
 wire pp_row65_30;
 wire pp_row65_31;
 wire pp_row65_32;
 wire pp_row65_33;
 wire pp_row65_4;
 wire pp_row65_5;
 wire pp_row65_6;
 wire pp_row65_7;
 wire pp_row65_8;
 wire pp_row65_9;
 wire pp_row66_1;
 wire pp_row66_10;
 wire pp_row66_11;
 wire pp_row66_12;
 wire pp_row66_13;
 wire pp_row66_14;
 wire pp_row66_15;
 wire pp_row66_16;
 wire pp_row66_17;
 wire pp_row66_18;
 wire pp_row66_19;
 wire pp_row66_2;
 wire pp_row66_20;
 wire pp_row66_21;
 wire pp_row66_22;
 wire pp_row66_23;
 wire pp_row66_24;
 wire pp_row66_25;
 wire pp_row66_26;
 wire pp_row66_27;
 wire pp_row66_28;
 wire pp_row66_29;
 wire pp_row66_3;
 wire pp_row66_30;
 wire pp_row66_31;
 wire pp_row66_32;
 wire pp_row66_33;
 wire pp_row66_4;
 wire pp_row66_5;
 wire pp_row66_6;
 wire pp_row66_7;
 wire pp_row66_8;
 wire pp_row66_9;
 wire pp_row67_0;
 wire pp_row67_1;
 wire pp_row67_10;
 wire pp_row67_11;
 wire pp_row67_12;
 wire pp_row67_13;
 wire pp_row67_14;
 wire pp_row67_15;
 wire pp_row67_16;
 wire pp_row67_17;
 wire pp_row67_18;
 wire pp_row67_19;
 wire pp_row67_2;
 wire pp_row67_20;
 wire pp_row67_21;
 wire pp_row67_22;
 wire pp_row67_23;
 wire pp_row67_24;
 wire pp_row67_25;
 wire pp_row67_26;
 wire pp_row67_27;
 wire pp_row67_28;
 wire pp_row67_29;
 wire pp_row67_3;
 wire pp_row67_30;
 wire pp_row67_31;
 wire pp_row67_32;
 wire pp_row67_33;
 wire pp_row67_4;
 wire pp_row67_5;
 wire pp_row67_6;
 wire pp_row67_7;
 wire pp_row67_8;
 wire pp_row67_9;
 wire pp_row68_1;
 wire pp_row68_10;
 wire pp_row68_11;
 wire pp_row68_12;
 wire pp_row68_13;
 wire pp_row68_14;
 wire pp_row68_15;
 wire pp_row68_16;
 wire pp_row68_17;
 wire pp_row68_18;
 wire pp_row68_19;
 wire pp_row68_2;
 wire pp_row68_20;
 wire pp_row68_21;
 wire pp_row68_22;
 wire pp_row68_23;
 wire pp_row68_24;
 wire pp_row68_25;
 wire pp_row68_26;
 wire pp_row68_27;
 wire pp_row68_28;
 wire pp_row68_29;
 wire pp_row68_3;
 wire pp_row68_30;
 wire pp_row68_31;
 wire pp_row68_32;
 wire pp_row68_4;
 wire pp_row68_5;
 wire pp_row68_6;
 wire pp_row68_7;
 wire pp_row68_8;
 wire pp_row68_9;
 wire pp_row69_0;
 wire pp_row69_1;
 wire pp_row69_10;
 wire pp_row69_11;
 wire pp_row69_12;
 wire pp_row69_13;
 wire pp_row69_14;
 wire pp_row69_15;
 wire pp_row69_16;
 wire pp_row69_17;
 wire pp_row69_18;
 wire pp_row69_19;
 wire pp_row69_2;
 wire pp_row69_20;
 wire pp_row69_21;
 wire pp_row69_22;
 wire pp_row69_23;
 wire pp_row69_24;
 wire pp_row69_25;
 wire pp_row69_26;
 wire pp_row69_27;
 wire pp_row69_28;
 wire pp_row69_29;
 wire pp_row69_3;
 wire pp_row69_30;
 wire pp_row69_31;
 wire pp_row69_4;
 wire pp_row69_5;
 wire pp_row69_6;
 wire pp_row69_7;
 wire pp_row69_8;
 wire pp_row69_9;
 wire pp_row6_0;
 wire pp_row6_1;
 wire pp_row6_2;
 wire pp_row6_3;
 wire pp_row6_4;
 wire pp_row6_5;
 wire pp_row70_1;
 wire pp_row70_10;
 wire pp_row70_11;
 wire pp_row70_12;
 wire pp_row70_13;
 wire pp_row70_14;
 wire pp_row70_15;
 wire pp_row70_16;
 wire pp_row70_17;
 wire pp_row70_18;
 wire pp_row70_19;
 wire pp_row70_2;
 wire pp_row70_20;
 wire pp_row70_21;
 wire pp_row70_22;
 wire pp_row70_23;
 wire pp_row70_24;
 wire pp_row70_25;
 wire pp_row70_26;
 wire pp_row70_27;
 wire pp_row70_28;
 wire pp_row70_29;
 wire pp_row70_3;
 wire pp_row70_30;
 wire pp_row70_31;
 wire pp_row70_4;
 wire pp_row70_5;
 wire pp_row70_6;
 wire pp_row70_7;
 wire pp_row70_8;
 wire pp_row70_9;
 wire pp_row71_0;
 wire pp_row71_1;
 wire pp_row71_10;
 wire pp_row71_11;
 wire pp_row71_12;
 wire pp_row71_13;
 wire pp_row71_14;
 wire pp_row71_15;
 wire pp_row71_16;
 wire pp_row71_17;
 wire pp_row71_18;
 wire pp_row71_19;
 wire pp_row71_2;
 wire pp_row71_20;
 wire pp_row71_21;
 wire pp_row71_22;
 wire pp_row71_23;
 wire pp_row71_24;
 wire pp_row71_25;
 wire pp_row71_26;
 wire pp_row71_27;
 wire pp_row71_28;
 wire pp_row71_29;
 wire pp_row71_3;
 wire pp_row71_30;
 wire pp_row71_4;
 wire pp_row71_5;
 wire pp_row71_6;
 wire pp_row71_7;
 wire pp_row71_8;
 wire pp_row71_9;
 wire pp_row72_1;
 wire pp_row72_10;
 wire pp_row72_11;
 wire pp_row72_12;
 wire pp_row72_13;
 wire pp_row72_14;
 wire pp_row72_15;
 wire pp_row72_16;
 wire pp_row72_17;
 wire pp_row72_18;
 wire pp_row72_19;
 wire pp_row72_2;
 wire pp_row72_20;
 wire pp_row72_21;
 wire pp_row72_22;
 wire pp_row72_23;
 wire pp_row72_24;
 wire pp_row72_25;
 wire pp_row72_26;
 wire pp_row72_27;
 wire pp_row72_28;
 wire pp_row72_29;
 wire pp_row72_3;
 wire pp_row72_30;
 wire pp_row72_4;
 wire pp_row72_5;
 wire pp_row72_6;
 wire pp_row72_7;
 wire pp_row72_8;
 wire pp_row72_9;
 wire pp_row73_0;
 wire pp_row73_1;
 wire pp_row73_10;
 wire pp_row73_11;
 wire pp_row73_12;
 wire pp_row73_13;
 wire pp_row73_14;
 wire pp_row73_15;
 wire pp_row73_16;
 wire pp_row73_17;
 wire pp_row73_18;
 wire pp_row73_19;
 wire pp_row73_2;
 wire pp_row73_20;
 wire pp_row73_21;
 wire pp_row73_22;
 wire pp_row73_23;
 wire pp_row73_24;
 wire pp_row73_25;
 wire pp_row73_26;
 wire pp_row73_27;
 wire pp_row73_28;
 wire pp_row73_29;
 wire pp_row73_3;
 wire pp_row73_4;
 wire pp_row73_5;
 wire pp_row73_6;
 wire pp_row73_7;
 wire pp_row73_8;
 wire pp_row73_9;
 wire pp_row74_1;
 wire pp_row74_10;
 wire pp_row74_11;
 wire pp_row74_12;
 wire pp_row74_13;
 wire pp_row74_14;
 wire pp_row74_15;
 wire pp_row74_16;
 wire pp_row74_17;
 wire pp_row74_18;
 wire pp_row74_19;
 wire pp_row74_2;
 wire pp_row74_20;
 wire pp_row74_21;
 wire pp_row74_22;
 wire pp_row74_23;
 wire pp_row74_24;
 wire pp_row74_25;
 wire pp_row74_26;
 wire pp_row74_27;
 wire pp_row74_28;
 wire pp_row74_29;
 wire pp_row74_3;
 wire pp_row74_4;
 wire pp_row74_5;
 wire pp_row74_6;
 wire pp_row74_7;
 wire pp_row74_8;
 wire pp_row74_9;
 wire pp_row75_0;
 wire pp_row75_1;
 wire pp_row75_10;
 wire pp_row75_11;
 wire pp_row75_12;
 wire pp_row75_13;
 wire pp_row75_14;
 wire pp_row75_15;
 wire pp_row75_16;
 wire pp_row75_17;
 wire pp_row75_18;
 wire pp_row75_19;
 wire pp_row75_2;
 wire pp_row75_20;
 wire pp_row75_21;
 wire pp_row75_22;
 wire pp_row75_23;
 wire pp_row75_24;
 wire pp_row75_25;
 wire pp_row75_26;
 wire pp_row75_27;
 wire pp_row75_28;
 wire pp_row75_3;
 wire pp_row75_4;
 wire pp_row75_5;
 wire pp_row75_6;
 wire pp_row75_7;
 wire pp_row75_8;
 wire pp_row75_9;
 wire pp_row76_1;
 wire pp_row76_10;
 wire pp_row76_11;
 wire pp_row76_12;
 wire pp_row76_13;
 wire pp_row76_14;
 wire pp_row76_15;
 wire pp_row76_16;
 wire pp_row76_17;
 wire pp_row76_18;
 wire pp_row76_19;
 wire pp_row76_2;
 wire pp_row76_20;
 wire pp_row76_21;
 wire pp_row76_22;
 wire pp_row76_23;
 wire pp_row76_24;
 wire pp_row76_25;
 wire pp_row76_26;
 wire pp_row76_27;
 wire pp_row76_28;
 wire pp_row76_3;
 wire pp_row76_4;
 wire pp_row76_5;
 wire pp_row76_6;
 wire pp_row76_7;
 wire pp_row76_8;
 wire pp_row76_9;
 wire pp_row77_0;
 wire pp_row77_1;
 wire pp_row77_10;
 wire pp_row77_11;
 wire pp_row77_12;
 wire pp_row77_13;
 wire pp_row77_14;
 wire pp_row77_15;
 wire pp_row77_16;
 wire pp_row77_17;
 wire pp_row77_18;
 wire pp_row77_19;
 wire pp_row77_2;
 wire pp_row77_20;
 wire pp_row77_21;
 wire pp_row77_22;
 wire pp_row77_23;
 wire pp_row77_24;
 wire pp_row77_25;
 wire pp_row77_26;
 wire pp_row77_27;
 wire pp_row77_3;
 wire pp_row77_4;
 wire pp_row77_5;
 wire pp_row77_6;
 wire pp_row77_7;
 wire pp_row77_8;
 wire pp_row77_9;
 wire pp_row78_1;
 wire pp_row78_10;
 wire pp_row78_11;
 wire pp_row78_12;
 wire pp_row78_13;
 wire pp_row78_14;
 wire pp_row78_15;
 wire pp_row78_16;
 wire pp_row78_17;
 wire pp_row78_18;
 wire pp_row78_19;
 wire pp_row78_2;
 wire pp_row78_20;
 wire pp_row78_21;
 wire pp_row78_22;
 wire pp_row78_23;
 wire pp_row78_24;
 wire pp_row78_25;
 wire pp_row78_26;
 wire pp_row78_27;
 wire pp_row78_3;
 wire pp_row78_4;
 wire pp_row78_5;
 wire pp_row78_6;
 wire pp_row78_7;
 wire pp_row78_8;
 wire pp_row78_9;
 wire pp_row79_0;
 wire pp_row79_1;
 wire pp_row79_10;
 wire pp_row79_11;
 wire pp_row79_12;
 wire pp_row79_13;
 wire pp_row79_14;
 wire pp_row79_15;
 wire pp_row79_16;
 wire pp_row79_17;
 wire pp_row79_18;
 wire pp_row79_19;
 wire pp_row79_2;
 wire pp_row79_20;
 wire pp_row79_21;
 wire pp_row79_22;
 wire pp_row79_23;
 wire pp_row79_24;
 wire pp_row79_25;
 wire pp_row79_26;
 wire pp_row79_3;
 wire pp_row79_4;
 wire pp_row79_5;
 wire pp_row79_6;
 wire pp_row79_7;
 wire pp_row79_8;
 wire pp_row79_9;
 wire pp_row7_0;
 wire pp_row7_1;
 wire pp_row7_2;
 wire pp_row7_3;
 wire pp_row7_4;
 wire pp_row80_1;
 wire pp_row80_10;
 wire pp_row80_11;
 wire pp_row80_12;
 wire pp_row80_13;
 wire pp_row80_14;
 wire pp_row80_15;
 wire pp_row80_16;
 wire pp_row80_17;
 wire pp_row80_18;
 wire pp_row80_19;
 wire pp_row80_2;
 wire pp_row80_20;
 wire pp_row80_21;
 wire pp_row80_22;
 wire pp_row80_23;
 wire pp_row80_24;
 wire pp_row80_25;
 wire pp_row80_26;
 wire pp_row80_3;
 wire pp_row80_4;
 wire pp_row80_5;
 wire pp_row80_6;
 wire pp_row80_7;
 wire pp_row80_8;
 wire pp_row80_9;
 wire pp_row81_0;
 wire pp_row81_1;
 wire pp_row81_10;
 wire pp_row81_11;
 wire pp_row81_12;
 wire pp_row81_13;
 wire pp_row81_14;
 wire pp_row81_15;
 wire pp_row81_16;
 wire pp_row81_17;
 wire pp_row81_18;
 wire pp_row81_19;
 wire pp_row81_2;
 wire pp_row81_20;
 wire pp_row81_21;
 wire pp_row81_22;
 wire pp_row81_23;
 wire pp_row81_24;
 wire pp_row81_25;
 wire pp_row81_3;
 wire pp_row81_4;
 wire pp_row81_5;
 wire pp_row81_6;
 wire pp_row81_7;
 wire pp_row81_8;
 wire pp_row81_9;
 wire pp_row82_1;
 wire pp_row82_10;
 wire pp_row82_11;
 wire pp_row82_12;
 wire pp_row82_13;
 wire pp_row82_14;
 wire pp_row82_15;
 wire pp_row82_16;
 wire pp_row82_17;
 wire pp_row82_18;
 wire pp_row82_19;
 wire pp_row82_2;
 wire pp_row82_20;
 wire pp_row82_21;
 wire pp_row82_22;
 wire pp_row82_23;
 wire pp_row82_24;
 wire pp_row82_25;
 wire pp_row82_3;
 wire pp_row82_4;
 wire pp_row82_5;
 wire pp_row82_6;
 wire pp_row82_7;
 wire pp_row82_8;
 wire pp_row82_9;
 wire pp_row83_0;
 wire pp_row83_1;
 wire pp_row83_10;
 wire pp_row83_11;
 wire pp_row83_12;
 wire pp_row83_13;
 wire pp_row83_14;
 wire pp_row83_15;
 wire pp_row83_16;
 wire pp_row83_17;
 wire pp_row83_18;
 wire pp_row83_19;
 wire pp_row83_2;
 wire pp_row83_20;
 wire pp_row83_21;
 wire pp_row83_22;
 wire pp_row83_23;
 wire pp_row83_24;
 wire pp_row83_3;
 wire pp_row83_4;
 wire pp_row83_5;
 wire pp_row83_6;
 wire pp_row83_7;
 wire pp_row83_8;
 wire pp_row83_9;
 wire pp_row84_1;
 wire pp_row84_10;
 wire pp_row84_11;
 wire pp_row84_12;
 wire pp_row84_13;
 wire pp_row84_14;
 wire pp_row84_15;
 wire pp_row84_16;
 wire pp_row84_17;
 wire pp_row84_18;
 wire pp_row84_19;
 wire pp_row84_2;
 wire pp_row84_20;
 wire pp_row84_21;
 wire pp_row84_22;
 wire pp_row84_23;
 wire pp_row84_24;
 wire pp_row84_3;
 wire pp_row84_4;
 wire pp_row84_5;
 wire pp_row84_6;
 wire pp_row84_7;
 wire pp_row84_8;
 wire pp_row84_9;
 wire pp_row85_0;
 wire pp_row85_1;
 wire pp_row85_10;
 wire pp_row85_11;
 wire pp_row85_12;
 wire pp_row85_13;
 wire pp_row85_14;
 wire pp_row85_15;
 wire pp_row85_16;
 wire pp_row85_17;
 wire pp_row85_18;
 wire pp_row85_19;
 wire pp_row85_2;
 wire pp_row85_20;
 wire pp_row85_21;
 wire pp_row85_22;
 wire pp_row85_23;
 wire pp_row85_3;
 wire pp_row85_4;
 wire pp_row85_5;
 wire pp_row85_6;
 wire pp_row85_7;
 wire pp_row85_8;
 wire pp_row85_9;
 wire pp_row86_1;
 wire pp_row86_10;
 wire pp_row86_11;
 wire pp_row86_12;
 wire pp_row86_13;
 wire pp_row86_14;
 wire pp_row86_15;
 wire pp_row86_16;
 wire pp_row86_17;
 wire pp_row86_18;
 wire pp_row86_19;
 wire pp_row86_2;
 wire pp_row86_20;
 wire pp_row86_21;
 wire pp_row86_22;
 wire pp_row86_23;
 wire pp_row86_3;
 wire pp_row86_4;
 wire pp_row86_5;
 wire pp_row86_6;
 wire pp_row86_7;
 wire pp_row86_8;
 wire pp_row86_9;
 wire pp_row87_0;
 wire pp_row87_1;
 wire pp_row87_10;
 wire pp_row87_11;
 wire pp_row87_12;
 wire pp_row87_13;
 wire pp_row87_14;
 wire pp_row87_15;
 wire pp_row87_16;
 wire pp_row87_17;
 wire pp_row87_18;
 wire pp_row87_19;
 wire pp_row87_2;
 wire pp_row87_20;
 wire pp_row87_21;
 wire pp_row87_22;
 wire pp_row87_3;
 wire pp_row87_4;
 wire pp_row87_5;
 wire pp_row87_6;
 wire pp_row87_7;
 wire pp_row87_8;
 wire pp_row87_9;
 wire pp_row88_1;
 wire pp_row88_10;
 wire pp_row88_11;
 wire pp_row88_12;
 wire pp_row88_13;
 wire pp_row88_14;
 wire pp_row88_15;
 wire pp_row88_16;
 wire pp_row88_17;
 wire pp_row88_18;
 wire pp_row88_19;
 wire pp_row88_2;
 wire pp_row88_20;
 wire pp_row88_21;
 wire pp_row88_22;
 wire pp_row88_3;
 wire pp_row88_4;
 wire pp_row88_5;
 wire pp_row88_6;
 wire pp_row88_7;
 wire pp_row88_8;
 wire pp_row88_9;
 wire pp_row89_0;
 wire pp_row89_1;
 wire pp_row89_10;
 wire pp_row89_11;
 wire pp_row89_12;
 wire pp_row89_13;
 wire pp_row89_14;
 wire pp_row89_15;
 wire pp_row89_16;
 wire pp_row89_17;
 wire pp_row89_18;
 wire pp_row89_19;
 wire pp_row89_2;
 wire pp_row89_20;
 wire pp_row89_21;
 wire pp_row89_3;
 wire pp_row89_4;
 wire pp_row89_5;
 wire pp_row89_6;
 wire pp_row89_7;
 wire pp_row89_8;
 wire pp_row89_9;
 wire pp_row8_0;
 wire pp_row8_1;
 wire pp_row8_2;
 wire pp_row8_3;
 wire pp_row8_4;
 wire pp_row8_5;
 wire pp_row8_6;
 wire pp_row90_1;
 wire pp_row90_10;
 wire pp_row90_11;
 wire pp_row90_12;
 wire pp_row90_13;
 wire pp_row90_14;
 wire pp_row90_15;
 wire pp_row90_16;
 wire pp_row90_17;
 wire pp_row90_18;
 wire pp_row90_19;
 wire pp_row90_2;
 wire pp_row90_20;
 wire pp_row90_21;
 wire pp_row90_3;
 wire pp_row90_4;
 wire pp_row90_5;
 wire pp_row90_6;
 wire pp_row90_7;
 wire pp_row90_8;
 wire pp_row90_9;
 wire pp_row91_0;
 wire pp_row91_1;
 wire pp_row91_10;
 wire pp_row91_11;
 wire pp_row91_12;
 wire pp_row91_13;
 wire pp_row91_14;
 wire pp_row91_15;
 wire pp_row91_16;
 wire pp_row91_17;
 wire pp_row91_18;
 wire pp_row91_19;
 wire pp_row91_2;
 wire pp_row91_20;
 wire pp_row91_3;
 wire pp_row91_4;
 wire pp_row91_5;
 wire pp_row91_6;
 wire pp_row91_7;
 wire pp_row91_8;
 wire pp_row91_9;
 wire pp_row92_1;
 wire pp_row92_10;
 wire pp_row92_11;
 wire pp_row92_12;
 wire pp_row92_13;
 wire pp_row92_14;
 wire pp_row92_15;
 wire pp_row92_16;
 wire pp_row92_17;
 wire pp_row92_18;
 wire pp_row92_19;
 wire pp_row92_2;
 wire pp_row92_20;
 wire pp_row92_3;
 wire pp_row92_4;
 wire pp_row92_5;
 wire pp_row92_6;
 wire pp_row92_7;
 wire pp_row92_8;
 wire pp_row92_9;
 wire pp_row93_0;
 wire pp_row93_1;
 wire pp_row93_10;
 wire pp_row93_11;
 wire pp_row93_12;
 wire pp_row93_13;
 wire pp_row93_14;
 wire pp_row93_15;
 wire pp_row93_16;
 wire pp_row93_17;
 wire pp_row93_18;
 wire pp_row93_19;
 wire pp_row93_2;
 wire pp_row93_3;
 wire pp_row93_4;
 wire pp_row93_5;
 wire pp_row93_6;
 wire pp_row93_7;
 wire pp_row93_8;
 wire pp_row93_9;
 wire pp_row94_1;
 wire pp_row94_10;
 wire pp_row94_11;
 wire pp_row94_12;
 wire pp_row94_13;
 wire pp_row94_14;
 wire pp_row94_15;
 wire pp_row94_16;
 wire pp_row94_17;
 wire pp_row94_18;
 wire pp_row94_19;
 wire pp_row94_2;
 wire pp_row94_3;
 wire pp_row94_4;
 wire pp_row94_5;
 wire pp_row94_6;
 wire pp_row94_7;
 wire pp_row94_8;
 wire pp_row94_9;
 wire pp_row95_0;
 wire pp_row95_1;
 wire pp_row95_10;
 wire pp_row95_11;
 wire pp_row95_12;
 wire pp_row95_13;
 wire pp_row95_14;
 wire pp_row95_15;
 wire pp_row95_16;
 wire pp_row95_17;
 wire pp_row95_18;
 wire pp_row95_2;
 wire pp_row95_3;
 wire pp_row95_4;
 wire pp_row95_5;
 wire pp_row95_6;
 wire pp_row95_7;
 wire pp_row95_8;
 wire pp_row95_9;
 wire pp_row96_1;
 wire pp_row96_10;
 wire pp_row96_11;
 wire pp_row96_12;
 wire pp_row96_13;
 wire pp_row96_14;
 wire pp_row96_15;
 wire pp_row96_16;
 wire pp_row96_17;
 wire pp_row96_18;
 wire pp_row96_2;
 wire pp_row96_3;
 wire pp_row96_4;
 wire pp_row96_5;
 wire pp_row96_6;
 wire pp_row96_7;
 wire pp_row96_8;
 wire pp_row96_9;
 wire pp_row97_0;
 wire pp_row97_1;
 wire pp_row97_10;
 wire pp_row97_11;
 wire pp_row97_12;
 wire pp_row97_13;
 wire pp_row97_14;
 wire pp_row97_15;
 wire pp_row97_16;
 wire pp_row97_17;
 wire pp_row97_2;
 wire pp_row97_3;
 wire pp_row97_4;
 wire pp_row97_5;
 wire pp_row97_6;
 wire pp_row97_7;
 wire pp_row97_8;
 wire pp_row97_9;
 wire pp_row98_1;
 wire pp_row98_10;
 wire pp_row98_11;
 wire pp_row98_12;
 wire pp_row98_13;
 wire pp_row98_14;
 wire pp_row98_15;
 wire pp_row98_16;
 wire pp_row98_17;
 wire pp_row98_2;
 wire pp_row98_3;
 wire pp_row98_4;
 wire pp_row98_5;
 wire pp_row98_6;
 wire pp_row98_7;
 wire pp_row98_8;
 wire pp_row98_9;
 wire pp_row99_0;
 wire pp_row99_1;
 wire pp_row99_10;
 wire pp_row99_11;
 wire pp_row99_12;
 wire pp_row99_13;
 wire pp_row99_14;
 wire pp_row99_15;
 wire pp_row99_16;
 wire pp_row99_2;
 wire pp_row99_3;
 wire pp_row99_4;
 wire pp_row99_5;
 wire pp_row99_6;
 wire pp_row99_7;
 wire pp_row99_8;
 wire pp_row99_9;
 wire pp_row9_0;
 wire pp_row9_1;
 wire pp_row9_2;
 wire pp_row9_3;
 wire pp_row9_4;
 wire pp_row9_5;
 wire s;
 wire \s$1001 ;
 wire \s$1003 ;
 wire \s$1005 ;
 wire \s$1007 ;
 wire \s$1009 ;
 wire \s$101 ;
 wire \s$1011 ;
 wire \s$1013 ;
 wire \s$1015 ;
 wire \s$1017 ;
 wire \s$1019 ;
 wire \s$1021 ;
 wire \s$1023 ;
 wire \s$1025 ;
 wire \s$1027 ;
 wire \s$1029 ;
 wire \s$103 ;
 wire \s$1031 ;
 wire \s$1033 ;
 wire \s$1035 ;
 wire \s$1037 ;
 wire \s$1039 ;
 wire \s$1041 ;
 wire \s$1043 ;
 wire \s$1045 ;
 wire \s$1047 ;
 wire \s$1049 ;
 wire \s$105 ;
 wire \s$1051 ;
 wire \s$1053 ;
 wire \s$1055 ;
 wire \s$1057 ;
 wire \s$1059 ;
 wire \s$1061 ;
 wire \s$1063 ;
 wire \s$1065 ;
 wire \s$1067 ;
 wire \s$1069 ;
 wire \s$107 ;
 wire \s$1071 ;
 wire \s$1073 ;
 wire \s$1075 ;
 wire \s$1077 ;
 wire \s$1079 ;
 wire \s$1081 ;
 wire \s$1083 ;
 wire \s$1085 ;
 wire \s$1087 ;
 wire \s$1089 ;
 wire \s$109 ;
 wire \s$1091 ;
 wire \s$1093 ;
 wire \s$1095 ;
 wire \s$1097 ;
 wire \s$1099 ;
 wire \s$11 ;
 wire \s$1101 ;
 wire \s$1103 ;
 wire \s$1105 ;
 wire \s$1107 ;
 wire \s$1109 ;
 wire \s$111 ;
 wire \s$1111 ;
 wire \s$1113 ;
 wire \s$1115 ;
 wire \s$1117 ;
 wire \s$1119 ;
 wire \s$1121 ;
 wire \s$1123 ;
 wire \s$1125 ;
 wire \s$1127 ;
 wire \s$1129 ;
 wire \s$113 ;
 wire \s$1131 ;
 wire \s$1133 ;
 wire \s$1135 ;
 wire \s$1137 ;
 wire \s$1139 ;
 wire \s$1141 ;
 wire \s$1143 ;
 wire \s$1145 ;
 wire \s$1147 ;
 wire \s$1149 ;
 wire \s$115 ;
 wire \s$1151 ;
 wire \s$1153 ;
 wire \s$1155 ;
 wire \s$1157 ;
 wire \s$1159 ;
 wire \s$1161 ;
 wire \s$1163 ;
 wire \s$1165 ;
 wire \s$1167 ;
 wire \s$1169 ;
 wire \s$117 ;
 wire \s$1171 ;
 wire \s$1173 ;
 wire \s$1175 ;
 wire \s$1177 ;
 wire \s$1179 ;
 wire \s$1181 ;
 wire \s$1183 ;
 wire \s$1185 ;
 wire \s$1187 ;
 wire \s$1189 ;
 wire \s$119 ;
 wire \s$1191 ;
 wire \s$1193 ;
 wire \s$1195 ;
 wire \s$1197 ;
 wire \s$1199 ;
 wire \s$1201 ;
 wire \s$1203 ;
 wire \s$1205 ;
 wire \s$1207 ;
 wire \s$1209 ;
 wire \s$121 ;
 wire \s$1211 ;
 wire \s$1213 ;
 wire \s$1215 ;
 wire \s$1217 ;
 wire \s$1219 ;
 wire \s$1221 ;
 wire \s$1223 ;
 wire \s$1225 ;
 wire \s$1227 ;
 wire \s$1229 ;
 wire \s$123 ;
 wire \s$1231 ;
 wire \s$1233 ;
 wire \s$1235 ;
 wire \s$1237 ;
 wire \s$1239 ;
 wire \s$1241 ;
 wire \s$1243 ;
 wire \s$1245 ;
 wire \s$1247 ;
 wire \s$1249 ;
 wire \s$125 ;
 wire \s$1251 ;
 wire \s$1253 ;
 wire \s$1255 ;
 wire \s$1257 ;
 wire \s$1259 ;
 wire \s$1261 ;
 wire \s$1263 ;
 wire \s$1265 ;
 wire \s$1267 ;
 wire \s$1269 ;
 wire \s$127 ;
 wire \s$1271 ;
 wire \s$1273 ;
 wire \s$1275 ;
 wire \s$1277 ;
 wire \s$1279 ;
 wire \s$1281 ;
 wire \s$1283 ;
 wire \s$1285 ;
 wire \s$1287 ;
 wire \s$1289 ;
 wire \s$129 ;
 wire \s$1291 ;
 wire \s$1293 ;
 wire \s$1295 ;
 wire \s$1297 ;
 wire \s$1299 ;
 wire \s$13 ;
 wire \s$1301 ;
 wire \s$1303 ;
 wire \s$1305 ;
 wire \s$1307 ;
 wire \s$1309 ;
 wire \s$131 ;
 wire \s$1311 ;
 wire \s$1313 ;
 wire \s$1315 ;
 wire \s$1317 ;
 wire \s$1319 ;
 wire \s$1321 ;
 wire \s$1323 ;
 wire \s$1325 ;
 wire \s$1327 ;
 wire \s$1329 ;
 wire \s$133 ;
 wire \s$1331 ;
 wire \s$1333 ;
 wire \s$1335 ;
 wire \s$1337 ;
 wire \s$1339 ;
 wire \s$1341 ;
 wire \s$1343 ;
 wire \s$1345 ;
 wire \s$1347 ;
 wire \s$1349 ;
 wire \s$135 ;
 wire \s$1351 ;
 wire \s$1353 ;
 wire \s$1355 ;
 wire \s$1357 ;
 wire \s$1359 ;
 wire \s$1361 ;
 wire \s$1363 ;
 wire \s$1365 ;
 wire \s$1367 ;
 wire \s$1369 ;
 wire \s$137 ;
 wire \s$1371 ;
 wire \s$1373 ;
 wire \s$1375 ;
 wire \s$1377 ;
 wire \s$1379 ;
 wire \s$1381 ;
 wire \s$1383 ;
 wire \s$1385 ;
 wire \s$1387 ;
 wire \s$1389 ;
 wire \s$139 ;
 wire \s$1391 ;
 wire \s$1393 ;
 wire \s$1395 ;
 wire \s$1397 ;
 wire \s$1399 ;
 wire \s$1401 ;
 wire \s$1403 ;
 wire \s$1405 ;
 wire \s$1407 ;
 wire \s$1409 ;
 wire \s$141 ;
 wire \s$1411 ;
 wire \s$1413 ;
 wire \s$1415 ;
 wire \s$1417 ;
 wire \s$1419 ;
 wire \s$1421 ;
 wire \s$1423 ;
 wire \s$1425 ;
 wire \s$1427 ;
 wire \s$1429 ;
 wire \s$143 ;
 wire \s$1431 ;
 wire \s$1433 ;
 wire \s$1435 ;
 wire \s$1437 ;
 wire \s$1439 ;
 wire \s$1441 ;
 wire \s$1443 ;
 wire \s$1445 ;
 wire \s$1447 ;
 wire \s$1449 ;
 wire \s$145 ;
 wire \s$1451 ;
 wire \s$1453 ;
 wire \s$1455 ;
 wire \s$1457 ;
 wire \s$1459 ;
 wire \s$1461 ;
 wire \s$1463 ;
 wire \s$1465 ;
 wire \s$1467 ;
 wire \s$1469 ;
 wire \s$147 ;
 wire \s$1471 ;
 wire \s$1473 ;
 wire \s$1475 ;
 wire \s$1477 ;
 wire \s$1479 ;
 wire \s$1481 ;
 wire \s$1483 ;
 wire \s$1485 ;
 wire \s$1487 ;
 wire \s$1489 ;
 wire \s$149 ;
 wire \s$1491 ;
 wire \s$1493 ;
 wire \s$1495 ;
 wire \s$1497 ;
 wire \s$1499 ;
 wire \s$15 ;
 wire \s$1501 ;
 wire \s$1503 ;
 wire \s$1505 ;
 wire \s$1507 ;
 wire \s$1509 ;
 wire \s$151 ;
 wire \s$1511 ;
 wire \s$1513 ;
 wire \s$1515 ;
 wire \s$1517 ;
 wire \s$1519 ;
 wire \s$1521 ;
 wire \s$1523 ;
 wire \s$1525 ;
 wire \s$1527 ;
 wire \s$1529 ;
 wire \s$153 ;
 wire \s$1531 ;
 wire \s$1533 ;
 wire \s$1535 ;
 wire \s$1537 ;
 wire \s$1539 ;
 wire \s$1541 ;
 wire \s$1543 ;
 wire \s$1545 ;
 wire \s$1547 ;
 wire \s$1549 ;
 wire \s$155 ;
 wire \s$1551 ;
 wire \s$1553 ;
 wire \s$1555 ;
 wire \s$1557 ;
 wire \s$1559 ;
 wire \s$1561 ;
 wire \s$1563 ;
 wire \s$1565 ;
 wire \s$1567 ;
 wire \s$1569 ;
 wire \s$157 ;
 wire \s$1571 ;
 wire \s$1573 ;
 wire \s$1575 ;
 wire \s$1577 ;
 wire \s$1579 ;
 wire \s$1581 ;
 wire \s$1583 ;
 wire \s$1585 ;
 wire \s$1587 ;
 wire \s$1589 ;
 wire \s$159 ;
 wire \s$1591 ;
 wire \s$1593 ;
 wire \s$1595 ;
 wire \s$1597 ;
 wire \s$1599 ;
 wire \s$1601 ;
 wire \s$1603 ;
 wire \s$1605 ;
 wire \s$1607 ;
 wire \s$1609 ;
 wire \s$161 ;
 wire \s$1611 ;
 wire \s$1613 ;
 wire \s$1615 ;
 wire \s$1617 ;
 wire \s$1619 ;
 wire \s$1621 ;
 wire \s$1623 ;
 wire \s$1625 ;
 wire \s$1627 ;
 wire \s$1629 ;
 wire \s$163 ;
 wire \s$1631 ;
 wire \s$1633 ;
 wire \s$1635 ;
 wire \s$1637 ;
 wire \s$1639 ;
 wire \s$1641 ;
 wire \s$1643 ;
 wire \s$1645 ;
 wire \s$1647 ;
 wire \s$1649 ;
 wire \s$165 ;
 wire \s$1651 ;
 wire \s$1653 ;
 wire \s$1655 ;
 wire \s$1657 ;
 wire \s$1659 ;
 wire \s$1661 ;
 wire \s$1663 ;
 wire \s$1665 ;
 wire \s$1667 ;
 wire \s$1669 ;
 wire \s$167 ;
 wire \s$1671 ;
 wire \s$1673 ;
 wire \s$1675 ;
 wire \s$1677 ;
 wire \s$1679 ;
 wire \s$1681 ;
 wire \s$1683 ;
 wire \s$1685 ;
 wire \s$1687 ;
 wire \s$1689 ;
 wire \s$169 ;
 wire \s$1691 ;
 wire \s$1693 ;
 wire \s$1695 ;
 wire \s$1697 ;
 wire \s$1699 ;
 wire \s$17 ;
 wire \s$1701 ;
 wire \s$1703 ;
 wire \s$1705 ;
 wire \s$1707 ;
 wire \s$1709 ;
 wire \s$171 ;
 wire \s$1711 ;
 wire \s$1713 ;
 wire \s$1715 ;
 wire \s$1717 ;
 wire \s$1719 ;
 wire \s$1721 ;
 wire \s$1723 ;
 wire \s$1725 ;
 wire \s$1727 ;
 wire \s$1729 ;
 wire \s$173 ;
 wire \s$1731 ;
 wire \s$1733 ;
 wire \s$1735 ;
 wire \s$1737 ;
 wire \s$1739 ;
 wire \s$1741 ;
 wire \s$1743 ;
 wire \s$1745 ;
 wire \s$1747 ;
 wire \s$1749 ;
 wire \s$175 ;
 wire \s$1751 ;
 wire \s$1753 ;
 wire \s$1755 ;
 wire \s$1757 ;
 wire \s$1759 ;
 wire \s$1761 ;
 wire \s$1763 ;
 wire \s$1765 ;
 wire \s$1767 ;
 wire \s$1769 ;
 wire \s$177 ;
 wire \s$1771 ;
 wire \s$1773 ;
 wire \s$1775 ;
 wire \s$1777 ;
 wire \s$1779 ;
 wire \s$1781 ;
 wire \s$1783 ;
 wire \s$1785 ;
 wire \s$1787 ;
 wire \s$1789 ;
 wire \s$179 ;
 wire \s$1791 ;
 wire \s$1793 ;
 wire \s$1795 ;
 wire \s$1797 ;
 wire \s$1799 ;
 wire \s$1801 ;
 wire \s$1803 ;
 wire \s$1805 ;
 wire \s$1807 ;
 wire \s$1809 ;
 wire \s$181 ;
 wire \s$1811 ;
 wire \s$1813 ;
 wire \s$1815 ;
 wire \s$1817 ;
 wire \s$1819 ;
 wire \s$1821 ;
 wire \s$1823 ;
 wire \s$1825 ;
 wire \s$1827 ;
 wire \s$1829 ;
 wire \s$183 ;
 wire \s$1831 ;
 wire \s$1833 ;
 wire \s$1835 ;
 wire \s$1837 ;
 wire \s$1839 ;
 wire \s$1841 ;
 wire \s$1843 ;
 wire \s$1845 ;
 wire \s$1847 ;
 wire \s$1849 ;
 wire \s$185 ;
 wire \s$1851 ;
 wire \s$1853 ;
 wire \s$1855 ;
 wire \s$1857 ;
 wire \s$1859 ;
 wire \s$1861 ;
 wire \s$1863 ;
 wire \s$1865 ;
 wire \s$1867 ;
 wire \s$1869 ;
 wire \s$187 ;
 wire \s$1871 ;
 wire \s$1873 ;
 wire \s$1875 ;
 wire \s$1877 ;
 wire \s$1879 ;
 wire \s$1881 ;
 wire \s$1883 ;
 wire \s$1885 ;
 wire \s$1887 ;
 wire \s$1889 ;
 wire \s$189 ;
 wire \s$1891 ;
 wire \s$1893 ;
 wire \s$1895 ;
 wire \s$1897 ;
 wire \s$1899 ;
 wire \s$19 ;
 wire \s$1901 ;
 wire \s$1903 ;
 wire \s$1905 ;
 wire \s$1907 ;
 wire \s$1909 ;
 wire \s$191 ;
 wire \s$1911 ;
 wire \s$1913 ;
 wire \s$1915 ;
 wire \s$1917 ;
 wire \s$1919 ;
 wire \s$1921 ;
 wire \s$1923 ;
 wire \s$1925 ;
 wire \s$1927 ;
 wire \s$1929 ;
 wire \s$193 ;
 wire \s$1931 ;
 wire \s$1933 ;
 wire \s$1935 ;
 wire \s$1937 ;
 wire \s$1939 ;
 wire \s$1941 ;
 wire \s$1943 ;
 wire \s$1945 ;
 wire \s$1947 ;
 wire \s$1949 ;
 wire \s$195 ;
 wire \s$1951 ;
 wire \s$1953 ;
 wire \s$1955 ;
 wire \s$1957 ;
 wire \s$1959 ;
 wire \s$1961 ;
 wire \s$1963 ;
 wire \s$1965 ;
 wire \s$1967 ;
 wire \s$1969 ;
 wire \s$197 ;
 wire \s$1971 ;
 wire \s$1973 ;
 wire \s$1975 ;
 wire \s$1977 ;
 wire \s$1979 ;
 wire \s$1981 ;
 wire \s$1983 ;
 wire \s$1985 ;
 wire \s$1987 ;
 wire \s$1989 ;
 wire \s$199 ;
 wire \s$1991 ;
 wire \s$1993 ;
 wire \s$1995 ;
 wire \s$1997 ;
 wire \s$1999 ;
 wire \s$2001 ;
 wire \s$2003 ;
 wire \s$2005 ;
 wire \s$2007 ;
 wire \s$2009 ;
 wire \s$201 ;
 wire \s$2011 ;
 wire \s$2013 ;
 wire \s$2015 ;
 wire \s$2017 ;
 wire \s$2019 ;
 wire \s$2021 ;
 wire \s$2023 ;
 wire \s$2025 ;
 wire \s$2027 ;
 wire \s$2029 ;
 wire \s$203 ;
 wire \s$2031 ;
 wire \s$2033 ;
 wire \s$2035 ;
 wire \s$2037 ;
 wire \s$2039 ;
 wire \s$2041 ;
 wire \s$2043 ;
 wire \s$2045 ;
 wire \s$2047 ;
 wire \s$2049 ;
 wire \s$205 ;
 wire \s$2051 ;
 wire \s$2053 ;
 wire \s$2055 ;
 wire \s$2057 ;
 wire \s$2059 ;
 wire \s$2061 ;
 wire \s$2063 ;
 wire \s$2065 ;
 wire \s$2067 ;
 wire \s$2069 ;
 wire \s$207 ;
 wire \s$2071 ;
 wire \s$2073 ;
 wire \s$2075 ;
 wire \s$2077 ;
 wire \s$2079 ;
 wire \s$2081 ;
 wire \s$2083 ;
 wire \s$2085 ;
 wire \s$2087 ;
 wire \s$2089 ;
 wire \s$209 ;
 wire \s$2091 ;
 wire \s$2093 ;
 wire \s$2095 ;
 wire \s$2097 ;
 wire \s$2099 ;
 wire \s$21 ;
 wire \s$2101 ;
 wire \s$2103 ;
 wire \s$2105 ;
 wire \s$2107 ;
 wire \s$2109 ;
 wire \s$211 ;
 wire \s$2111 ;
 wire \s$2113 ;
 wire \s$2115 ;
 wire \s$2117 ;
 wire \s$2119 ;
 wire \s$2121 ;
 wire \s$2123 ;
 wire \s$2125 ;
 wire \s$2127 ;
 wire \s$2129 ;
 wire \s$213 ;
 wire \s$2131 ;
 wire \s$2133 ;
 wire \s$2135 ;
 wire \s$2137 ;
 wire \s$2139 ;
 wire \s$2141 ;
 wire \s$2143 ;
 wire \s$2145 ;
 wire \s$2147 ;
 wire \s$2149 ;
 wire \s$215 ;
 wire \s$2151 ;
 wire \s$2153 ;
 wire \s$2155 ;
 wire \s$2157 ;
 wire \s$2159 ;
 wire \s$2161 ;
 wire \s$2163 ;
 wire \s$2165 ;
 wire \s$2167 ;
 wire \s$2169 ;
 wire \s$217 ;
 wire \s$2171 ;
 wire \s$2173 ;
 wire \s$2175 ;
 wire \s$2177 ;
 wire \s$2179 ;
 wire \s$2181 ;
 wire \s$2183 ;
 wire \s$2185 ;
 wire \s$2187 ;
 wire \s$2189 ;
 wire \s$219 ;
 wire \s$2191 ;
 wire \s$2193 ;
 wire \s$2195 ;
 wire \s$2197 ;
 wire \s$2199 ;
 wire \s$2201 ;
 wire \s$2203 ;
 wire \s$2205 ;
 wire \s$2207 ;
 wire \s$2209 ;
 wire \s$221 ;
 wire \s$2211 ;
 wire \s$2213 ;
 wire \s$2215 ;
 wire \s$2217 ;
 wire \s$2219 ;
 wire \s$2221 ;
 wire \s$2223 ;
 wire \s$2225 ;
 wire \s$2227 ;
 wire \s$2229 ;
 wire \s$223 ;
 wire \s$2231 ;
 wire \s$2233 ;
 wire \s$2235 ;
 wire \s$2237 ;
 wire \s$2239 ;
 wire \s$2241 ;
 wire \s$2243 ;
 wire \s$2245 ;
 wire \s$2247 ;
 wire \s$2249 ;
 wire \s$225 ;
 wire \s$2251 ;
 wire \s$2253 ;
 wire \s$2255 ;
 wire \s$2257 ;
 wire \s$2259 ;
 wire \s$2261 ;
 wire \s$2263 ;
 wire \s$2265 ;
 wire \s$2267 ;
 wire \s$2269 ;
 wire \s$227 ;
 wire \s$2271 ;
 wire \s$2273 ;
 wire \s$2275 ;
 wire \s$2277 ;
 wire \s$2279 ;
 wire \s$2281 ;
 wire \s$2283 ;
 wire \s$2285 ;
 wire \s$2287 ;
 wire \s$2289 ;
 wire \s$229 ;
 wire \s$2291 ;
 wire \s$2293 ;
 wire \s$2295 ;
 wire \s$2297 ;
 wire \s$2299 ;
 wire \s$23 ;
 wire \s$2301 ;
 wire \s$2303 ;
 wire \s$2305 ;
 wire \s$2307 ;
 wire \s$2309 ;
 wire \s$231 ;
 wire \s$2311 ;
 wire \s$2313 ;
 wire \s$2315 ;
 wire \s$2317 ;
 wire \s$2319 ;
 wire \s$2321 ;
 wire \s$2323 ;
 wire \s$2325 ;
 wire \s$2327 ;
 wire \s$2329 ;
 wire \s$233 ;
 wire \s$2331 ;
 wire \s$2333 ;
 wire \s$2335 ;
 wire \s$2337 ;
 wire \s$2339 ;
 wire \s$2341 ;
 wire \s$2343 ;
 wire \s$2345 ;
 wire \s$2347 ;
 wire \s$2349 ;
 wire \s$235 ;
 wire \s$2351 ;
 wire \s$2353 ;
 wire \s$2355 ;
 wire \s$2357 ;
 wire \s$2359 ;
 wire \s$2361 ;
 wire \s$2363 ;
 wire \s$2365 ;
 wire \s$2367 ;
 wire \s$2369 ;
 wire \s$237 ;
 wire \s$2371 ;
 wire \s$2373 ;
 wire \s$2375 ;
 wire \s$2377 ;
 wire \s$2379 ;
 wire \s$2381 ;
 wire \s$2383 ;
 wire \s$2385 ;
 wire \s$2387 ;
 wire \s$2389 ;
 wire \s$239 ;
 wire \s$2391 ;
 wire \s$2393 ;
 wire \s$2395 ;
 wire \s$2397 ;
 wire \s$2399 ;
 wire \s$2401 ;
 wire \s$2403 ;
 wire \s$2405 ;
 wire \s$2407 ;
 wire \s$2409 ;
 wire \s$241 ;
 wire \s$2411 ;
 wire \s$2413 ;
 wire \s$2415 ;
 wire \s$2417 ;
 wire \s$2419 ;
 wire \s$2421 ;
 wire \s$2423 ;
 wire \s$2425 ;
 wire \s$2427 ;
 wire \s$2429 ;
 wire \s$243 ;
 wire \s$2431 ;
 wire \s$2433 ;
 wire \s$2435 ;
 wire \s$2437 ;
 wire \s$2439 ;
 wire \s$2441 ;
 wire \s$2443 ;
 wire \s$2445 ;
 wire \s$2447 ;
 wire \s$2449 ;
 wire \s$245 ;
 wire \s$2451 ;
 wire \s$2453 ;
 wire \s$2455 ;
 wire \s$2457 ;
 wire \s$2459 ;
 wire \s$2461 ;
 wire \s$2463 ;
 wire \s$2465 ;
 wire \s$2467 ;
 wire \s$2469 ;
 wire \s$247 ;
 wire \s$2471 ;
 wire \s$2473 ;
 wire \s$2475 ;
 wire \s$2477 ;
 wire \s$2479 ;
 wire \s$2481 ;
 wire \s$2483 ;
 wire \s$2485 ;
 wire \s$2487 ;
 wire \s$2489 ;
 wire \s$249 ;
 wire \s$2491 ;
 wire \s$2493 ;
 wire \s$2495 ;
 wire \s$2497 ;
 wire \s$2499 ;
 wire \s$25 ;
 wire \s$2501 ;
 wire \s$2503 ;
 wire \s$2505 ;
 wire \s$2507 ;
 wire \s$2509 ;
 wire \s$251 ;
 wire \s$2511 ;
 wire \s$2513 ;
 wire \s$2515 ;
 wire \s$2517 ;
 wire \s$2519 ;
 wire \s$2521 ;
 wire \s$2523 ;
 wire \s$2525 ;
 wire \s$2527 ;
 wire \s$2529 ;
 wire \s$253 ;
 wire \s$2531 ;
 wire \s$2533 ;
 wire \s$2535 ;
 wire \s$2537 ;
 wire \s$2539 ;
 wire \s$2541 ;
 wire \s$2543 ;
 wire \s$2545 ;
 wire \s$2547 ;
 wire \s$2549 ;
 wire \s$255 ;
 wire \s$2551 ;
 wire \s$2553 ;
 wire \s$2555 ;
 wire \s$2557 ;
 wire \s$2559 ;
 wire \s$2561 ;
 wire \s$2563 ;
 wire \s$2565 ;
 wire \s$2567 ;
 wire \s$2569 ;
 wire \s$257 ;
 wire \s$2571 ;
 wire \s$2573 ;
 wire \s$2575 ;
 wire \s$2577 ;
 wire \s$2579 ;
 wire \s$2581 ;
 wire \s$2583 ;
 wire \s$2585 ;
 wire \s$2587 ;
 wire \s$2589 ;
 wire \s$259 ;
 wire \s$2591 ;
 wire \s$2593 ;
 wire \s$2595 ;
 wire \s$2597 ;
 wire \s$2599 ;
 wire \s$2601 ;
 wire \s$2603 ;
 wire \s$2605 ;
 wire \s$2607 ;
 wire \s$2609 ;
 wire \s$261 ;
 wire \s$2611 ;
 wire \s$2613 ;
 wire \s$2615 ;
 wire \s$2617 ;
 wire \s$2619 ;
 wire \s$2621 ;
 wire \s$2623 ;
 wire \s$2625 ;
 wire \s$2627 ;
 wire \s$2629 ;
 wire \s$263 ;
 wire \s$2631 ;
 wire \s$2633 ;
 wire \s$2635 ;
 wire \s$2637 ;
 wire \s$2639 ;
 wire \s$2641 ;
 wire \s$2643 ;
 wire \s$2645 ;
 wire \s$2647 ;
 wire \s$2649 ;
 wire \s$265 ;
 wire \s$2651 ;
 wire \s$2653 ;
 wire \s$2655 ;
 wire \s$2657 ;
 wire \s$2659 ;
 wire \s$2661 ;
 wire \s$2663 ;
 wire \s$2665 ;
 wire \s$2667 ;
 wire \s$2669 ;
 wire \s$267 ;
 wire \s$2671 ;
 wire \s$2673 ;
 wire \s$2675 ;
 wire \s$2677 ;
 wire \s$2679 ;
 wire \s$2681 ;
 wire \s$2683 ;
 wire \s$2685 ;
 wire \s$2687 ;
 wire \s$2689 ;
 wire \s$269 ;
 wire \s$2691 ;
 wire \s$2693 ;
 wire \s$2695 ;
 wire \s$2697 ;
 wire \s$2699 ;
 wire \s$27 ;
 wire \s$2701 ;
 wire \s$2703 ;
 wire \s$2705 ;
 wire \s$2707 ;
 wire \s$2709 ;
 wire \s$271 ;
 wire \s$2711 ;
 wire \s$2713 ;
 wire \s$2715 ;
 wire \s$2717 ;
 wire \s$2719 ;
 wire \s$2721 ;
 wire \s$2723 ;
 wire \s$2725 ;
 wire \s$2727 ;
 wire \s$2729 ;
 wire \s$273 ;
 wire \s$2731 ;
 wire \s$2733 ;
 wire \s$2735 ;
 wire \s$2737 ;
 wire \s$2739 ;
 wire \s$2741 ;
 wire \s$2743 ;
 wire \s$2745 ;
 wire \s$2747 ;
 wire \s$2749 ;
 wire \s$275 ;
 wire \s$2751 ;
 wire \s$2753 ;
 wire \s$2755 ;
 wire \s$2757 ;
 wire \s$2759 ;
 wire \s$2761 ;
 wire \s$2763 ;
 wire \s$2765 ;
 wire \s$2767 ;
 wire \s$2769 ;
 wire \s$277 ;
 wire \s$2771 ;
 wire \s$2773 ;
 wire \s$2775 ;
 wire \s$2777 ;
 wire \s$2779 ;
 wire \s$2781 ;
 wire \s$2783 ;
 wire \s$2785 ;
 wire \s$2787 ;
 wire \s$2789 ;
 wire \s$279 ;
 wire \s$2791 ;
 wire \s$2793 ;
 wire \s$2795 ;
 wire \s$2797 ;
 wire \s$2799 ;
 wire \s$2801 ;
 wire \s$2803 ;
 wire \s$2805 ;
 wire \s$2807 ;
 wire \s$2809 ;
 wire \s$281 ;
 wire \s$2811 ;
 wire \s$2813 ;
 wire \s$2815 ;
 wire \s$2817 ;
 wire \s$2819 ;
 wire \s$2821 ;
 wire \s$2823 ;
 wire \s$2825 ;
 wire \s$2827 ;
 wire \s$2829 ;
 wire \s$283 ;
 wire \s$2831 ;
 wire \s$2833 ;
 wire \s$2835 ;
 wire \s$2837 ;
 wire \s$2839 ;
 wire \s$2841 ;
 wire \s$2843 ;
 wire \s$2845 ;
 wire \s$2847 ;
 wire \s$2849 ;
 wire \s$285 ;
 wire \s$2851 ;
 wire \s$2853 ;
 wire \s$2855 ;
 wire \s$2857 ;
 wire \s$2859 ;
 wire \s$2861 ;
 wire \s$2863 ;
 wire \s$2865 ;
 wire \s$2867 ;
 wire \s$2869 ;
 wire \s$287 ;
 wire \s$2871 ;
 wire \s$2873 ;
 wire \s$2875 ;
 wire \s$2877 ;
 wire \s$2879 ;
 wire \s$2881 ;
 wire \s$2883 ;
 wire \s$2885 ;
 wire \s$2887 ;
 wire \s$2889 ;
 wire \s$289 ;
 wire \s$2891 ;
 wire \s$2893 ;
 wire \s$2895 ;
 wire \s$2897 ;
 wire \s$2899 ;
 wire \s$29 ;
 wire \s$2901 ;
 wire \s$2903 ;
 wire \s$2905 ;
 wire \s$2907 ;
 wire \s$2909 ;
 wire \s$291 ;
 wire \s$2911 ;
 wire \s$2913 ;
 wire \s$2915 ;
 wire \s$2917 ;
 wire \s$2919 ;
 wire \s$2921 ;
 wire \s$2923 ;
 wire \s$2925 ;
 wire \s$2927 ;
 wire \s$2929 ;
 wire \s$293 ;
 wire \s$2931 ;
 wire \s$2933 ;
 wire \s$2935 ;
 wire \s$2937 ;
 wire \s$2939 ;
 wire \s$2941 ;
 wire \s$2943 ;
 wire \s$2945 ;
 wire \s$2947 ;
 wire \s$2949 ;
 wire \s$295 ;
 wire \s$2951 ;
 wire \s$2953 ;
 wire \s$2955 ;
 wire \s$2957 ;
 wire \s$2959 ;
 wire \s$2961 ;
 wire \s$2963 ;
 wire \s$2965 ;
 wire \s$2967 ;
 wire \s$2969 ;
 wire \s$297 ;
 wire \s$2971 ;
 wire \s$2973 ;
 wire \s$2975 ;
 wire \s$2977 ;
 wire \s$2979 ;
 wire \s$2981 ;
 wire \s$2983 ;
 wire \s$2985 ;
 wire \s$2987 ;
 wire \s$2989 ;
 wire \s$299 ;
 wire \s$2991 ;
 wire \s$2993 ;
 wire \s$2995 ;
 wire \s$2997 ;
 wire \s$2999 ;
 wire \s$3 ;
 wire \s$3001 ;
 wire \s$3003 ;
 wire \s$3005 ;
 wire \s$3007 ;
 wire \s$3009 ;
 wire \s$301 ;
 wire \s$3011 ;
 wire \s$3013 ;
 wire \s$3015 ;
 wire \s$3017 ;
 wire \s$3019 ;
 wire \s$3021 ;
 wire \s$3023 ;
 wire \s$3025 ;
 wire \s$3027 ;
 wire \s$3029 ;
 wire \s$303 ;
 wire \s$3031 ;
 wire \s$3033 ;
 wire \s$3035 ;
 wire \s$3037 ;
 wire \s$3039 ;
 wire \s$3041 ;
 wire \s$3043 ;
 wire \s$3045 ;
 wire \s$3047 ;
 wire \s$3049 ;
 wire \s$305 ;
 wire \s$3051 ;
 wire \s$3053 ;
 wire \s$3055 ;
 wire \s$3057 ;
 wire \s$3059 ;
 wire \s$3061 ;
 wire \s$3063 ;
 wire \s$3065 ;
 wire \s$3067 ;
 wire \s$3069 ;
 wire \s$307 ;
 wire \s$3071 ;
 wire \s$3073 ;
 wire \s$3075 ;
 wire \s$3077 ;
 wire \s$3079 ;
 wire \s$3081 ;
 wire \s$3083 ;
 wire \s$3085 ;
 wire \s$3087 ;
 wire \s$3089 ;
 wire \s$309 ;
 wire \s$3091 ;
 wire \s$3093 ;
 wire \s$3095 ;
 wire \s$3097 ;
 wire \s$3099 ;
 wire \s$31 ;
 wire \s$3101 ;
 wire \s$3103 ;
 wire \s$3105 ;
 wire \s$3107 ;
 wire \s$3109 ;
 wire \s$311 ;
 wire \s$3111 ;
 wire \s$3113 ;
 wire \s$3115 ;
 wire \s$3117 ;
 wire \s$3119 ;
 wire \s$3121 ;
 wire \s$3123 ;
 wire \s$3125 ;
 wire \s$3127 ;
 wire \s$3129 ;
 wire \s$313 ;
 wire \s$3131 ;
 wire \s$3133 ;
 wire \s$3135 ;
 wire \s$3137 ;
 wire \s$3139 ;
 wire \s$3141 ;
 wire \s$3143 ;
 wire \s$3145 ;
 wire \s$3147 ;
 wire \s$3149 ;
 wire \s$315 ;
 wire \s$3151 ;
 wire \s$3153 ;
 wire \s$3155 ;
 wire \s$3157 ;
 wire \s$3159 ;
 wire \s$3161 ;
 wire \s$3163 ;
 wire \s$3165 ;
 wire \s$3167 ;
 wire \s$3169 ;
 wire \s$317 ;
 wire \s$3171 ;
 wire \s$3173 ;
 wire \s$3175 ;
 wire \s$3177 ;
 wire \s$3179 ;
 wire \s$3181 ;
 wire \s$3183 ;
 wire \s$3185 ;
 wire \s$3187 ;
 wire \s$3189 ;
 wire \s$319 ;
 wire \s$3191 ;
 wire \s$3193 ;
 wire \s$3195 ;
 wire \s$3197 ;
 wire \s$3199 ;
 wire \s$3201 ;
 wire \s$3203 ;
 wire \s$3205 ;
 wire \s$3207 ;
 wire \s$3209 ;
 wire \s$321 ;
 wire \s$3211 ;
 wire \s$3213 ;
 wire \s$3215 ;
 wire \s$3217 ;
 wire \s$3219 ;
 wire \s$3221 ;
 wire \s$3223 ;
 wire \s$3225 ;
 wire \s$3227 ;
 wire \s$3229 ;
 wire \s$323 ;
 wire \s$3231 ;
 wire \s$3233 ;
 wire \s$3235 ;
 wire \s$3237 ;
 wire \s$3239 ;
 wire \s$3241 ;
 wire \s$3243 ;
 wire \s$3245 ;
 wire \s$3247 ;
 wire \s$3249 ;
 wire \s$325 ;
 wire \s$3251 ;
 wire \s$3253 ;
 wire \s$3255 ;
 wire \s$3257 ;
 wire \s$3259 ;
 wire \s$3261 ;
 wire \s$3263 ;
 wire \s$3265 ;
 wire \s$3267 ;
 wire \s$3269 ;
 wire \s$327 ;
 wire \s$3271 ;
 wire \s$3273 ;
 wire \s$3275 ;
 wire \s$3277 ;
 wire \s$3279 ;
 wire \s$3281 ;
 wire \s$3283 ;
 wire \s$3285 ;
 wire \s$3287 ;
 wire \s$3289 ;
 wire \s$329 ;
 wire \s$3291 ;
 wire \s$3293 ;
 wire \s$3295 ;
 wire \s$3297 ;
 wire \s$3299 ;
 wire \s$33 ;
 wire \s$3301 ;
 wire \s$3303 ;
 wire \s$3305 ;
 wire \s$3307 ;
 wire \s$3309 ;
 wire \s$331 ;
 wire \s$3311 ;
 wire \s$3313 ;
 wire \s$3315 ;
 wire \s$3317 ;
 wire \s$3319 ;
 wire \s$3321 ;
 wire \s$3323 ;
 wire \s$3325 ;
 wire \s$3327 ;
 wire \s$3329 ;
 wire \s$333 ;
 wire \s$3331 ;
 wire \s$3333 ;
 wire \s$3335 ;
 wire \s$3337 ;
 wire \s$3339 ;
 wire \s$3341 ;
 wire \s$3343 ;
 wire \s$3345 ;
 wire \s$3347 ;
 wire \s$3349 ;
 wire \s$335 ;
 wire \s$3351 ;
 wire \s$3353 ;
 wire \s$3355 ;
 wire \s$3357 ;
 wire \s$3359 ;
 wire \s$3361 ;
 wire \s$3363 ;
 wire \s$3365 ;
 wire \s$3367 ;
 wire \s$3369 ;
 wire \s$337 ;
 wire \s$3371 ;
 wire \s$3373 ;
 wire \s$3375 ;
 wire \s$3377 ;
 wire \s$3379 ;
 wire \s$3381 ;
 wire \s$3383 ;
 wire \s$3385 ;
 wire \s$3387 ;
 wire \s$3389 ;
 wire \s$339 ;
 wire \s$3391 ;
 wire \s$3393 ;
 wire \s$3395 ;
 wire \s$3397 ;
 wire \s$3399 ;
 wire \s$3401 ;
 wire \s$3403 ;
 wire \s$3405 ;
 wire \s$3407 ;
 wire \s$3409 ;
 wire \s$341 ;
 wire \s$3411 ;
 wire \s$3413 ;
 wire \s$3415 ;
 wire \s$3417 ;
 wire \s$3419 ;
 wire \s$3421 ;
 wire \s$3423 ;
 wire \s$3425 ;
 wire \s$3427 ;
 wire \s$3429 ;
 wire \s$343 ;
 wire \s$3431 ;
 wire \s$3433 ;
 wire \s$3435 ;
 wire \s$3437 ;
 wire \s$3439 ;
 wire \s$3441 ;
 wire \s$3443 ;
 wire \s$3445 ;
 wire \s$3447 ;
 wire \s$3449 ;
 wire \s$345 ;
 wire \s$3451 ;
 wire \s$3453 ;
 wire \s$3455 ;
 wire \s$3457 ;
 wire \s$3459 ;
 wire \s$3461 ;
 wire \s$3463 ;
 wire \s$3465 ;
 wire \s$3467 ;
 wire \s$3469 ;
 wire \s$347 ;
 wire \s$3471 ;
 wire \s$3473 ;
 wire \s$3475 ;
 wire \s$3477 ;
 wire \s$3479 ;
 wire \s$3481 ;
 wire \s$3483 ;
 wire \s$3485 ;
 wire \s$3487 ;
 wire \s$3489 ;
 wire \s$349 ;
 wire \s$3491 ;
 wire \s$3493 ;
 wire \s$3495 ;
 wire \s$3497 ;
 wire \s$3499 ;
 wire \s$35 ;
 wire \s$3501 ;
 wire \s$3503 ;
 wire \s$3505 ;
 wire \s$3507 ;
 wire \s$3509 ;
 wire \s$351 ;
 wire \s$3511 ;
 wire \s$3513 ;
 wire \s$3515 ;
 wire \s$3517 ;
 wire \s$3519 ;
 wire \s$3521 ;
 wire \s$3523 ;
 wire \s$3525 ;
 wire \s$3527 ;
 wire \s$3529 ;
 wire \s$353 ;
 wire \s$3531 ;
 wire \s$3533 ;
 wire \s$3535 ;
 wire \s$3537 ;
 wire \s$3539 ;
 wire \s$3541 ;
 wire \s$3543 ;
 wire \s$3545 ;
 wire \s$3547 ;
 wire \s$3549 ;
 wire \s$355 ;
 wire \s$3551 ;
 wire \s$3553 ;
 wire \s$3555 ;
 wire \s$3557 ;
 wire \s$3559 ;
 wire \s$3561 ;
 wire \s$3563 ;
 wire \s$3565 ;
 wire \s$3567 ;
 wire \s$3569 ;
 wire \s$357 ;
 wire \s$3571 ;
 wire \s$3573 ;
 wire \s$3575 ;
 wire \s$3577 ;
 wire \s$3579 ;
 wire \s$3581 ;
 wire \s$3583 ;
 wire \s$3585 ;
 wire \s$3587 ;
 wire \s$3589 ;
 wire \s$359 ;
 wire \s$3591 ;
 wire \s$3593 ;
 wire \s$3595 ;
 wire \s$3597 ;
 wire \s$3599 ;
 wire \s$3601 ;
 wire \s$3603 ;
 wire \s$3605 ;
 wire \s$3607 ;
 wire \s$3609 ;
 wire \s$361 ;
 wire \s$3611 ;
 wire \s$3613 ;
 wire \s$3615 ;
 wire \s$3617 ;
 wire \s$3619 ;
 wire \s$3621 ;
 wire \s$3623 ;
 wire \s$3625 ;
 wire \s$3627 ;
 wire \s$3629 ;
 wire \s$363 ;
 wire \s$3631 ;
 wire \s$3633 ;
 wire \s$3635 ;
 wire \s$3637 ;
 wire \s$3639 ;
 wire \s$3641 ;
 wire \s$3643 ;
 wire \s$3645 ;
 wire \s$3647 ;
 wire \s$3649 ;
 wire \s$365 ;
 wire \s$3651 ;
 wire \s$3653 ;
 wire \s$3655 ;
 wire \s$3657 ;
 wire \s$3659 ;
 wire \s$3661 ;
 wire \s$3663 ;
 wire \s$3665 ;
 wire \s$3667 ;
 wire \s$3669 ;
 wire \s$367 ;
 wire \s$3671 ;
 wire \s$3673 ;
 wire \s$3675 ;
 wire \s$3677 ;
 wire \s$3679 ;
 wire \s$3681 ;
 wire \s$3683 ;
 wire \s$3685 ;
 wire \s$3687 ;
 wire \s$3689 ;
 wire \s$369 ;
 wire \s$3691 ;
 wire \s$3693 ;
 wire \s$3695 ;
 wire \s$3697 ;
 wire \s$3699 ;
 wire \s$37 ;
 wire \s$3701 ;
 wire \s$3703 ;
 wire \s$3705 ;
 wire \s$3707 ;
 wire \s$3709 ;
 wire \s$371 ;
 wire \s$3711 ;
 wire \s$3713 ;
 wire \s$3715 ;
 wire \s$3717 ;
 wire \s$3719 ;
 wire \s$3721 ;
 wire \s$3723 ;
 wire \s$3725 ;
 wire \s$3727 ;
 wire \s$3729 ;
 wire \s$373 ;
 wire \s$3731 ;
 wire \s$3733 ;
 wire \s$3735 ;
 wire \s$3737 ;
 wire \s$3739 ;
 wire \s$3741 ;
 wire \s$3743 ;
 wire \s$3745 ;
 wire \s$3747 ;
 wire \s$3749 ;
 wire \s$375 ;
 wire \s$3751 ;
 wire \s$3753 ;
 wire \s$3755 ;
 wire \s$3757 ;
 wire \s$3759 ;
 wire \s$3761 ;
 wire \s$3763 ;
 wire \s$3765 ;
 wire \s$3767 ;
 wire \s$3769 ;
 wire \s$377 ;
 wire \s$3771 ;
 wire \s$3773 ;
 wire \s$3775 ;
 wire \s$3777 ;
 wire \s$3779 ;
 wire \s$3781 ;
 wire \s$3783 ;
 wire \s$3785 ;
 wire \s$3787 ;
 wire \s$3789 ;
 wire \s$379 ;
 wire \s$3791 ;
 wire \s$3793 ;
 wire \s$3795 ;
 wire \s$3797 ;
 wire \s$3799 ;
 wire \s$3801 ;
 wire \s$3803 ;
 wire \s$3805 ;
 wire \s$3807 ;
 wire \s$3809 ;
 wire \s$381 ;
 wire \s$3811 ;
 wire \s$3813 ;
 wire \s$3815 ;
 wire \s$3817 ;
 wire \s$3819 ;
 wire \s$3821 ;
 wire \s$3823 ;
 wire \s$3825 ;
 wire \s$3827 ;
 wire \s$3829 ;
 wire \s$383 ;
 wire \s$3831 ;
 wire \s$3833 ;
 wire \s$3835 ;
 wire \s$3837 ;
 wire \s$3839 ;
 wire \s$3841 ;
 wire \s$3843 ;
 wire \s$3845 ;
 wire \s$3847 ;
 wire \s$3849 ;
 wire \s$385 ;
 wire \s$3851 ;
 wire \s$3853 ;
 wire \s$3855 ;
 wire \s$3857 ;
 wire \s$3859 ;
 wire \s$3861 ;
 wire \s$3863 ;
 wire \s$3865 ;
 wire \s$3867 ;
 wire \s$3869 ;
 wire \s$387 ;
 wire \s$3871 ;
 wire \s$3873 ;
 wire \s$3875 ;
 wire \s$3877 ;
 wire \s$3879 ;
 wire \s$3881 ;
 wire \s$3883 ;
 wire \s$3885 ;
 wire \s$3887 ;
 wire \s$3889 ;
 wire \s$389 ;
 wire \s$3891 ;
 wire \s$3893 ;
 wire \s$3895 ;
 wire \s$3897 ;
 wire \s$3899 ;
 wire \s$39 ;
 wire \s$3901 ;
 wire \s$3903 ;
 wire \s$3905 ;
 wire \s$3907 ;
 wire \s$3909 ;
 wire \s$391 ;
 wire \s$3911 ;
 wire \s$3913 ;
 wire \s$3915 ;
 wire \s$3917 ;
 wire \s$3919 ;
 wire \s$3921 ;
 wire \s$3923 ;
 wire \s$3925 ;
 wire \s$3927 ;
 wire \s$3929 ;
 wire \s$393 ;
 wire \s$3931 ;
 wire \s$3933 ;
 wire \s$3935 ;
 wire \s$3937 ;
 wire \s$3939 ;
 wire \s$3941 ;
 wire \s$3943 ;
 wire \s$3945 ;
 wire \s$3947 ;
 wire \s$3949 ;
 wire \s$395 ;
 wire \s$3951 ;
 wire \s$3953 ;
 wire \s$3955 ;
 wire \s$3957 ;
 wire \s$3959 ;
 wire \s$3961 ;
 wire \s$3963 ;
 wire \s$3965 ;
 wire \s$3967 ;
 wire \s$3969 ;
 wire \s$397 ;
 wire \s$3971 ;
 wire \s$3973 ;
 wire \s$3975 ;
 wire \s$3977 ;
 wire \s$3979 ;
 wire \s$3981 ;
 wire \s$3983 ;
 wire \s$3985 ;
 wire \s$3987 ;
 wire \s$3989 ;
 wire \s$399 ;
 wire \s$3991 ;
 wire \s$3993 ;
 wire \s$3995 ;
 wire \s$3997 ;
 wire \s$3999 ;
 wire \s$4001 ;
 wire \s$4003 ;
 wire \s$4005 ;
 wire \s$4007 ;
 wire \s$4009 ;
 wire \s$401 ;
 wire \s$4011 ;
 wire \s$4013 ;
 wire \s$4015 ;
 wire \s$4017 ;
 wire \s$4019 ;
 wire \s$4021 ;
 wire \s$4023 ;
 wire \s$4025 ;
 wire \s$4027 ;
 wire \s$4029 ;
 wire \s$403 ;
 wire \s$4031 ;
 wire \s$4033 ;
 wire \s$4035 ;
 wire \s$4037 ;
 wire \s$4039 ;
 wire \s$4041 ;
 wire \s$4043 ;
 wire \s$4045 ;
 wire \s$4047 ;
 wire \s$4049 ;
 wire \s$405 ;
 wire \s$4051 ;
 wire \s$4053 ;
 wire \s$4055 ;
 wire \s$4057 ;
 wire \s$4059 ;
 wire \s$4061 ;
 wire \s$4063 ;
 wire \s$4065 ;
 wire \s$4067 ;
 wire \s$4069 ;
 wire \s$407 ;
 wire \s$4071 ;
 wire \s$4073 ;
 wire \s$4075 ;
 wire \s$4077 ;
 wire \s$4079 ;
 wire \s$4081 ;
 wire \s$4083 ;
 wire \s$4085 ;
 wire \s$4087 ;
 wire \s$4089 ;
 wire \s$409 ;
 wire \s$4091 ;
 wire \s$4093 ;
 wire \s$4095 ;
 wire \s$4097 ;
 wire \s$4099 ;
 wire \s$41 ;
 wire \s$4101 ;
 wire \s$4103 ;
 wire \s$4105 ;
 wire \s$4107 ;
 wire \s$4109 ;
 wire \s$411 ;
 wire \s$4111 ;
 wire \s$4113 ;
 wire \s$4115 ;
 wire \s$4117 ;
 wire \s$4119 ;
 wire \s$4121 ;
 wire \s$4123 ;
 wire \s$4125 ;
 wire \s$4127 ;
 wire \s$4129 ;
 wire \s$413 ;
 wire \s$4131 ;
 wire \s$4133 ;
 wire \s$4135 ;
 wire \s$4137 ;
 wire \s$4139 ;
 wire \s$4141 ;
 wire \s$4143 ;
 wire \s$4145 ;
 wire \s$4147 ;
 wire \s$4149 ;
 wire \s$415 ;
 wire \s$4151 ;
 wire \s$4153 ;
 wire \s$4155 ;
 wire \s$4157 ;
 wire \s$4159 ;
 wire \s$4161 ;
 wire \s$4163 ;
 wire \s$4165 ;
 wire \s$4167 ;
 wire \s$4169 ;
 wire \s$417 ;
 wire \s$4171 ;
 wire \s$4173 ;
 wire \s$4175 ;
 wire \s$4177 ;
 wire \s$4179 ;
 wire \s$4181 ;
 wire \s$4183 ;
 wire \s$4185 ;
 wire \s$4187 ;
 wire \s$4189 ;
 wire \s$419 ;
 wire \s$4191 ;
 wire \s$4193 ;
 wire \s$4195 ;
 wire \s$4197 ;
 wire \s$4199 ;
 wire \s$4201 ;
 wire \s$4203 ;
 wire \s$4205 ;
 wire \s$4207 ;
 wire \s$4209 ;
 wire \s$421 ;
 wire \s$4211 ;
 wire \s$4213 ;
 wire \s$4215 ;
 wire \s$4217 ;
 wire \s$4219 ;
 wire \s$4221 ;
 wire \s$4223 ;
 wire \s$4225 ;
 wire \s$4227 ;
 wire \s$4229 ;
 wire \s$423 ;
 wire \s$4231 ;
 wire \s$4233 ;
 wire \s$4235 ;
 wire \s$4237 ;
 wire \s$4239 ;
 wire \s$4241 ;
 wire \s$4243 ;
 wire \s$4245 ;
 wire \s$4247 ;
 wire \s$4249 ;
 wire \s$425 ;
 wire \s$4251 ;
 wire \s$4253 ;
 wire \s$4255 ;
 wire \s$4257 ;
 wire \s$4259 ;
 wire \s$4261 ;
 wire \s$4263 ;
 wire \s$4265 ;
 wire \s$4267 ;
 wire \s$4269 ;
 wire \s$427 ;
 wire \s$4271 ;
 wire \s$4273 ;
 wire \s$4275 ;
 wire \s$4277 ;
 wire \s$4279 ;
 wire \s$4281 ;
 wire \s$4283 ;
 wire \s$4285 ;
 wire \s$4287 ;
 wire \s$4289 ;
 wire \s$429 ;
 wire \s$4291 ;
 wire \s$4293 ;
 wire \s$4295 ;
 wire \s$4297 ;
 wire \s$4299 ;
 wire \s$43 ;
 wire \s$4301 ;
 wire \s$4303 ;
 wire \s$4305 ;
 wire \s$4307 ;
 wire \s$4309 ;
 wire \s$431 ;
 wire \s$4311 ;
 wire \s$4313 ;
 wire \s$4315 ;
 wire \s$4317 ;
 wire \s$4319 ;
 wire \s$4321 ;
 wire \s$4323 ;
 wire \s$4325 ;
 wire \s$4327 ;
 wire \s$4329 ;
 wire \s$433 ;
 wire \s$4331 ;
 wire \s$4333 ;
 wire \s$4335 ;
 wire \s$4337 ;
 wire \s$4339 ;
 wire \s$4341 ;
 wire \s$4343 ;
 wire \s$4345 ;
 wire \s$4347 ;
 wire \s$4349 ;
 wire \s$435 ;
 wire \s$4351 ;
 wire \s$4353 ;
 wire \s$4355 ;
 wire \s$4357 ;
 wire \s$4359 ;
 wire \s$4361 ;
 wire \s$4363 ;
 wire \s$4365 ;
 wire \s$4367 ;
 wire \s$4369 ;
 wire \s$437 ;
 wire \s$4371 ;
 wire \s$4373 ;
 wire \s$4375 ;
 wire \s$4377 ;
 wire \s$4379 ;
 wire \s$4381 ;
 wire \s$4383 ;
 wire \s$4385 ;
 wire \s$4387 ;
 wire \s$4389 ;
 wire \s$439 ;
 wire \s$4391 ;
 wire \s$4393 ;
 wire \s$4395 ;
 wire \s$4397 ;
 wire \s$4399 ;
 wire \s$4401 ;
 wire \s$4403 ;
 wire \s$4405 ;
 wire \s$4407 ;
 wire \s$441 ;
 wire \s$443 ;
 wire \s$445 ;
 wire \s$447 ;
 wire \s$449 ;
 wire \s$45 ;
 wire \s$451 ;
 wire \s$453 ;
 wire \s$455 ;
 wire \s$457 ;
 wire \s$459 ;
 wire \s$461 ;
 wire \s$463 ;
 wire \s$465 ;
 wire \s$467 ;
 wire \s$469 ;
 wire \s$47 ;
 wire \s$471 ;
 wire \s$473 ;
 wire \s$475 ;
 wire \s$477 ;
 wire \s$479 ;
 wire \s$481 ;
 wire \s$483 ;
 wire \s$485 ;
 wire \s$487 ;
 wire \s$489 ;
 wire \s$49 ;
 wire \s$491 ;
 wire \s$493 ;
 wire \s$495 ;
 wire \s$497 ;
 wire \s$499 ;
 wire \s$5 ;
 wire \s$501 ;
 wire \s$503 ;
 wire \s$505 ;
 wire \s$507 ;
 wire \s$509 ;
 wire \s$51 ;
 wire \s$511 ;
 wire \s$513 ;
 wire \s$515 ;
 wire \s$517 ;
 wire \s$519 ;
 wire \s$521 ;
 wire \s$523 ;
 wire \s$525 ;
 wire \s$527 ;
 wire \s$529 ;
 wire \s$53 ;
 wire \s$531 ;
 wire \s$533 ;
 wire \s$535 ;
 wire \s$537 ;
 wire \s$539 ;
 wire \s$541 ;
 wire \s$543 ;
 wire \s$545 ;
 wire \s$547 ;
 wire \s$549 ;
 wire \s$55 ;
 wire \s$551 ;
 wire \s$553 ;
 wire \s$555 ;
 wire \s$557 ;
 wire \s$559 ;
 wire \s$561 ;
 wire \s$563 ;
 wire \s$565 ;
 wire \s$567 ;
 wire \s$569 ;
 wire \s$57 ;
 wire \s$571 ;
 wire \s$573 ;
 wire \s$575 ;
 wire \s$577 ;
 wire \s$579 ;
 wire \s$581 ;
 wire \s$583 ;
 wire \s$585 ;
 wire \s$587 ;
 wire \s$589 ;
 wire \s$59 ;
 wire \s$591 ;
 wire \s$593 ;
 wire \s$595 ;
 wire \s$597 ;
 wire \s$599 ;
 wire \s$601 ;
 wire \s$603 ;
 wire \s$605 ;
 wire \s$607 ;
 wire \s$609 ;
 wire \s$61 ;
 wire \s$611 ;
 wire \s$613 ;
 wire \s$615 ;
 wire \s$617 ;
 wire \s$619 ;
 wire \s$621 ;
 wire \s$623 ;
 wire \s$625 ;
 wire \s$627 ;
 wire \s$629 ;
 wire \s$63 ;
 wire \s$631 ;
 wire \s$633 ;
 wire \s$635 ;
 wire \s$637 ;
 wire \s$639 ;
 wire \s$641 ;
 wire \s$643 ;
 wire \s$645 ;
 wire \s$647 ;
 wire \s$649 ;
 wire \s$65 ;
 wire \s$651 ;
 wire \s$653 ;
 wire \s$655 ;
 wire \s$657 ;
 wire \s$659 ;
 wire \s$661 ;
 wire \s$663 ;
 wire \s$665 ;
 wire \s$667 ;
 wire \s$669 ;
 wire \s$67 ;
 wire \s$671 ;
 wire \s$673 ;
 wire \s$675 ;
 wire \s$677 ;
 wire \s$679 ;
 wire \s$681 ;
 wire \s$683 ;
 wire \s$685 ;
 wire \s$687 ;
 wire \s$689 ;
 wire \s$69 ;
 wire \s$691 ;
 wire \s$693 ;
 wire \s$695 ;
 wire \s$697 ;
 wire \s$699 ;
 wire \s$7 ;
 wire \s$701 ;
 wire \s$703 ;
 wire \s$705 ;
 wire \s$707 ;
 wire \s$709 ;
 wire \s$71 ;
 wire \s$711 ;
 wire \s$713 ;
 wire \s$715 ;
 wire \s$717 ;
 wire \s$719 ;
 wire \s$721 ;
 wire \s$723 ;
 wire \s$725 ;
 wire \s$727 ;
 wire \s$729 ;
 wire \s$73 ;
 wire \s$731 ;
 wire \s$733 ;
 wire \s$735 ;
 wire \s$737 ;
 wire \s$739 ;
 wire \s$741 ;
 wire \s$743 ;
 wire \s$745 ;
 wire \s$747 ;
 wire \s$749 ;
 wire \s$75 ;
 wire \s$751 ;
 wire \s$753 ;
 wire \s$755 ;
 wire \s$757 ;
 wire \s$759 ;
 wire \s$761 ;
 wire \s$763 ;
 wire \s$765 ;
 wire \s$767 ;
 wire \s$769 ;
 wire \s$77 ;
 wire \s$771 ;
 wire \s$773 ;
 wire \s$775 ;
 wire \s$777 ;
 wire \s$779 ;
 wire \s$781 ;
 wire \s$783 ;
 wire \s$785 ;
 wire \s$787 ;
 wire \s$789 ;
 wire \s$79 ;
 wire \s$791 ;
 wire \s$793 ;
 wire \s$795 ;
 wire \s$797 ;
 wire \s$799 ;
 wire \s$801 ;
 wire \s$803 ;
 wire \s$805 ;
 wire \s$807 ;
 wire \s$809 ;
 wire \s$81 ;
 wire \s$811 ;
 wire \s$813 ;
 wire \s$815 ;
 wire \s$817 ;
 wire \s$819 ;
 wire \s$821 ;
 wire \s$823 ;
 wire \s$825 ;
 wire \s$827 ;
 wire \s$829 ;
 wire \s$83 ;
 wire \s$831 ;
 wire \s$833 ;
 wire \s$835 ;
 wire \s$837 ;
 wire \s$839 ;
 wire \s$841 ;
 wire \s$843 ;
 wire \s$845 ;
 wire \s$847 ;
 wire \s$849 ;
 wire \s$85 ;
 wire \s$851 ;
 wire \s$853 ;
 wire \s$855 ;
 wire \s$857 ;
 wire \s$859 ;
 wire \s$861 ;
 wire \s$863 ;
 wire \s$865 ;
 wire \s$867 ;
 wire \s$869 ;
 wire \s$87 ;
 wire \s$871 ;
 wire \s$873 ;
 wire \s$875 ;
 wire \s$877 ;
 wire \s$879 ;
 wire \s$881 ;
 wire \s$883 ;
 wire \s$885 ;
 wire \s$887 ;
 wire \s$889 ;
 wire \s$89 ;
 wire \s$891 ;
 wire \s$893 ;
 wire \s$895 ;
 wire \s$897 ;
 wire \s$899 ;
 wire \s$9 ;
 wire \s$901 ;
 wire \s$903 ;
 wire \s$905 ;
 wire \s$907 ;
 wire \s$909 ;
 wire \s$91 ;
 wire \s$911 ;
 wire \s$913 ;
 wire \s$915 ;
 wire \s$917 ;
 wire \s$919 ;
 wire \s$921 ;
 wire \s$923 ;
 wire \s$925 ;
 wire \s$927 ;
 wire \s$929 ;
 wire \s$93 ;
 wire \s$931 ;
 wire \s$933 ;
 wire \s$935 ;
 wire \s$937 ;
 wire \s$939 ;
 wire \s$941 ;
 wire \s$943 ;
 wire \s$945 ;
 wire \s$947 ;
 wire \s$949 ;
 wire \s$95 ;
 wire \s$951 ;
 wire \s$953 ;
 wire \s$955 ;
 wire \s$957 ;
 wire \s$959 ;
 wire \s$961 ;
 wire \s$963 ;
 wire \s$965 ;
 wire \s$967 ;
 wire \s$969 ;
 wire \s$97 ;
 wire \s$971 ;
 wire \s$973 ;
 wire \s$975 ;
 wire \s$977 ;
 wire \s$979 ;
 wire \s$981 ;
 wire \s$983 ;
 wire \s$985 ;
 wire \s$987 ;
 wire \s$989 ;
 wire \s$99 ;
 wire \s$991 ;
 wire \s$993 ;
 wire \s$995 ;
 wire \s$997 ;
 wire \s$999 ;
 wire sel_0;
 wire \sel_0$4477 ;
 wire \sel_0$4547 ;
 wire \sel_0$4617 ;
 wire \sel_0$4687 ;
 wire \sel_0$4757 ;
 wire \sel_0$4827 ;
 wire \sel_0$4897 ;
 wire \sel_0$4967 ;
 wire \sel_0$5037 ;
 wire \sel_0$5107 ;
 wire \sel_0$5177 ;
 wire \sel_0$5247 ;
 wire \sel_0$5317 ;
 wire \sel_0$5387 ;
 wire \sel_0$5457 ;
 wire \sel_0$5527 ;
 wire \sel_0$5597 ;
 wire \sel_0$5667 ;
 wire \sel_0$5737 ;
 wire \sel_0$5807 ;
 wire \sel_0$5877 ;
 wire \sel_0$5947 ;
 wire \sel_0$6017 ;
 wire \sel_0$6087 ;
 wire \sel_0$6157 ;
 wire \sel_0$6227 ;
 wire \sel_0$6297 ;
 wire \sel_0$6367 ;
 wire \sel_0$6437 ;
 wire \sel_0$6507 ;
 wire \sel_0$6577 ;
 wire \sel_0$6647 ;
 wire sel_1;
 wire \sel_1$4478 ;
 wire \sel_1$4548 ;
 wire \sel_1$4618 ;
 wire \sel_1$4688 ;
 wire \sel_1$4758 ;
 wire \sel_1$4828 ;
 wire \sel_1$4898 ;
 wire \sel_1$4968 ;
 wire \sel_1$5038 ;
 wire \sel_1$5108 ;
 wire \sel_1$5178 ;
 wire \sel_1$5248 ;
 wire \sel_1$5318 ;
 wire \sel_1$5388 ;
 wire \sel_1$5458 ;
 wire \sel_1$5528 ;
 wire \sel_1$5598 ;
 wire \sel_1$5668 ;
 wire \sel_1$5738 ;
 wire \sel_1$5808 ;
 wire \sel_1$5878 ;
 wire \sel_1$5948 ;
 wire \sel_1$6018 ;
 wire \sel_1$6088 ;
 wire \sel_1$6158 ;
 wire \sel_1$6228 ;
 wire \sel_1$6298 ;
 wire \sel_1$6368 ;
 wire \sel_1$6438 ;
 wire \sel_1$6508 ;
 wire \sel_1$6578 ;
 wire \sel_1$6648 ;
 wire t;
 wire \t$4410 ;
 wire \t$4411 ;
 wire \t$4412 ;
 wire \t$4413 ;
 wire \t$4414 ;
 wire \t$4415 ;
 wire \t$4416 ;
 wire \t$4417 ;
 wire \t$4418 ;
 wire \t$4419 ;
 wire \t$4420 ;
 wire \t$4421 ;
 wire \t$4422 ;
 wire \t$4423 ;
 wire \t$4424 ;
 wire \t$4425 ;
 wire \t$4426 ;
 wire \t$4427 ;
 wire \t$4428 ;
 wire \t$4429 ;
 wire \t$4430 ;
 wire \t$4431 ;
 wire \t$4432 ;
 wire \t$4433 ;
 wire \t$4434 ;
 wire \t$4435 ;
 wire \t$4436 ;
 wire \t$4437 ;
 wire \t$4438 ;
 wire \t$4439 ;
 wire \t$4440 ;
 wire \t$4441 ;
 wire \t$4442 ;
 wire \t$4443 ;
 wire \t$4444 ;
 wire \t$4445 ;
 wire \t$4446 ;
 wire \t$4447 ;
 wire \t$4448 ;
 wire \t$4449 ;
 wire \t$4450 ;
 wire \t$4451 ;
 wire \t$4452 ;
 wire \t$4453 ;
 wire \t$4454 ;
 wire \t$4455 ;
 wire \t$4456 ;
 wire \t$4457 ;
 wire \t$4458 ;
 wire \t$4459 ;
 wire \t$4460 ;
 wire \t$4461 ;
 wire \t$4462 ;
 wire \t$4463 ;
 wire \t$4464 ;
 wire \t$4465 ;
 wire \t$4466 ;
 wire \t$4467 ;
 wire \t$4468 ;
 wire \t$4469 ;
 wire \t$4470 ;
 wire \t$4471 ;
 wire \t$4472 ;
 wire \t$4473 ;
 wire \t$4474 ;
 wire \t$4476 ;
 wire \t$4479 ;
 wire \t$4480 ;
 wire \t$4481 ;
 wire \t$4482 ;
 wire \t$4483 ;
 wire \t$4484 ;
 wire \t$4485 ;
 wire \t$4486 ;
 wire \t$4487 ;
 wire \t$4488 ;
 wire \t$4489 ;
 wire \t$4490 ;
 wire \t$4491 ;
 wire \t$4492 ;
 wire \t$4493 ;
 wire \t$4494 ;
 wire \t$4495 ;
 wire \t$4496 ;
 wire \t$4497 ;
 wire \t$4498 ;
 wire \t$4499 ;
 wire \t$4500 ;
 wire \t$4501 ;
 wire \t$4502 ;
 wire \t$4503 ;
 wire \t$4504 ;
 wire \t$4505 ;
 wire \t$4506 ;
 wire \t$4507 ;
 wire \t$4508 ;
 wire \t$4509 ;
 wire \t$4510 ;
 wire \t$4511 ;
 wire \t$4512 ;
 wire \t$4513 ;
 wire \t$4514 ;
 wire \t$4515 ;
 wire \t$4516 ;
 wire \t$4517 ;
 wire \t$4518 ;
 wire \t$4519 ;
 wire \t$4520 ;
 wire \t$4521 ;
 wire \t$4522 ;
 wire \t$4523 ;
 wire \t$4524 ;
 wire \t$4525 ;
 wire \t$4526 ;
 wire \t$4527 ;
 wire \t$4528 ;
 wire \t$4529 ;
 wire \t$4530 ;
 wire \t$4531 ;
 wire \t$4532 ;
 wire \t$4533 ;
 wire \t$4534 ;
 wire \t$4535 ;
 wire \t$4536 ;
 wire \t$4537 ;
 wire \t$4538 ;
 wire \t$4539 ;
 wire \t$4540 ;
 wire \t$4541 ;
 wire \t$4542 ;
 wire \t$4543 ;
 wire \t$4546 ;
 wire \t$4549 ;
 wire \t$4550 ;
 wire \t$4551 ;
 wire \t$4552 ;
 wire \t$4553 ;
 wire \t$4554 ;
 wire \t$4555 ;
 wire \t$4556 ;
 wire \t$4557 ;
 wire \t$4558 ;
 wire \t$4559 ;
 wire \t$4560 ;
 wire \t$4561 ;
 wire \t$4562 ;
 wire \t$4563 ;
 wire \t$4564 ;
 wire \t$4565 ;
 wire \t$4566 ;
 wire \t$4567 ;
 wire \t$4568 ;
 wire \t$4569 ;
 wire \t$4570 ;
 wire \t$4571 ;
 wire \t$4572 ;
 wire \t$4573 ;
 wire \t$4574 ;
 wire \t$4575 ;
 wire \t$4576 ;
 wire \t$4577 ;
 wire \t$4578 ;
 wire \t$4579 ;
 wire \t$4580 ;
 wire \t$4581 ;
 wire \t$4582 ;
 wire \t$4583 ;
 wire \t$4584 ;
 wire \t$4585 ;
 wire \t$4586 ;
 wire \t$4587 ;
 wire \t$4588 ;
 wire \t$4589 ;
 wire \t$4590 ;
 wire \t$4591 ;
 wire \t$4592 ;
 wire \t$4593 ;
 wire \t$4594 ;
 wire \t$4595 ;
 wire \t$4596 ;
 wire \t$4597 ;
 wire \t$4598 ;
 wire \t$4599 ;
 wire \t$4600 ;
 wire \t$4601 ;
 wire \t$4602 ;
 wire \t$4603 ;
 wire \t$4604 ;
 wire \t$4605 ;
 wire \t$4606 ;
 wire \t$4607 ;
 wire \t$4608 ;
 wire \t$4609 ;
 wire \t$4610 ;
 wire \t$4611 ;
 wire \t$4612 ;
 wire \t$4613 ;
 wire \t$4616 ;
 wire \t$4619 ;
 wire \t$4620 ;
 wire \t$4621 ;
 wire \t$4622 ;
 wire \t$4623 ;
 wire \t$4624 ;
 wire \t$4625 ;
 wire \t$4626 ;
 wire \t$4627 ;
 wire \t$4628 ;
 wire \t$4629 ;
 wire \t$4630 ;
 wire \t$4631 ;
 wire \t$4632 ;
 wire \t$4633 ;
 wire \t$4634 ;
 wire \t$4635 ;
 wire \t$4636 ;
 wire \t$4637 ;
 wire \t$4638 ;
 wire \t$4639 ;
 wire \t$4640 ;
 wire \t$4641 ;
 wire \t$4642 ;
 wire \t$4643 ;
 wire \t$4644 ;
 wire \t$4645 ;
 wire \t$4646 ;
 wire \t$4647 ;
 wire \t$4648 ;
 wire \t$4649 ;
 wire \t$4650 ;
 wire \t$4651 ;
 wire \t$4652 ;
 wire \t$4653 ;
 wire \t$4654 ;
 wire \t$4655 ;
 wire \t$4656 ;
 wire \t$4657 ;
 wire \t$4658 ;
 wire \t$4659 ;
 wire \t$4660 ;
 wire \t$4661 ;
 wire \t$4662 ;
 wire \t$4663 ;
 wire \t$4664 ;
 wire \t$4665 ;
 wire \t$4666 ;
 wire \t$4667 ;
 wire \t$4668 ;
 wire \t$4669 ;
 wire \t$4670 ;
 wire \t$4671 ;
 wire \t$4672 ;
 wire \t$4673 ;
 wire \t$4674 ;
 wire \t$4675 ;
 wire \t$4676 ;
 wire \t$4677 ;
 wire \t$4678 ;
 wire \t$4679 ;
 wire \t$4680 ;
 wire \t$4681 ;
 wire \t$4682 ;
 wire \t$4683 ;
 wire \t$4686 ;
 wire \t$4689 ;
 wire \t$4690 ;
 wire \t$4691 ;
 wire \t$4692 ;
 wire \t$4693 ;
 wire \t$4694 ;
 wire \t$4695 ;
 wire \t$4696 ;
 wire \t$4697 ;
 wire \t$4698 ;
 wire \t$4699 ;
 wire \t$4700 ;
 wire \t$4701 ;
 wire \t$4702 ;
 wire \t$4703 ;
 wire \t$4704 ;
 wire \t$4705 ;
 wire \t$4706 ;
 wire \t$4707 ;
 wire \t$4708 ;
 wire \t$4709 ;
 wire \t$4710 ;
 wire \t$4711 ;
 wire \t$4712 ;
 wire \t$4713 ;
 wire \t$4714 ;
 wire \t$4715 ;
 wire \t$4716 ;
 wire \t$4717 ;
 wire \t$4718 ;
 wire \t$4719 ;
 wire \t$4720 ;
 wire \t$4721 ;
 wire \t$4722 ;
 wire \t$4723 ;
 wire \t$4724 ;
 wire \t$4725 ;
 wire \t$4726 ;
 wire \t$4727 ;
 wire \t$4728 ;
 wire \t$4729 ;
 wire \t$4730 ;
 wire \t$4731 ;
 wire \t$4732 ;
 wire \t$4733 ;
 wire \t$4734 ;
 wire \t$4735 ;
 wire \t$4736 ;
 wire \t$4737 ;
 wire \t$4738 ;
 wire \t$4739 ;
 wire \t$4740 ;
 wire \t$4741 ;
 wire \t$4742 ;
 wire \t$4743 ;
 wire \t$4744 ;
 wire \t$4745 ;
 wire \t$4746 ;
 wire \t$4747 ;
 wire \t$4748 ;
 wire \t$4749 ;
 wire \t$4750 ;
 wire \t$4751 ;
 wire \t$4752 ;
 wire \t$4753 ;
 wire \t$4756 ;
 wire \t$4759 ;
 wire \t$4760 ;
 wire \t$4761 ;
 wire \t$4762 ;
 wire \t$4763 ;
 wire \t$4764 ;
 wire \t$4765 ;
 wire \t$4766 ;
 wire \t$4767 ;
 wire \t$4768 ;
 wire \t$4769 ;
 wire \t$4770 ;
 wire \t$4771 ;
 wire \t$4772 ;
 wire \t$4773 ;
 wire \t$4774 ;
 wire \t$4775 ;
 wire \t$4776 ;
 wire \t$4777 ;
 wire \t$4778 ;
 wire \t$4779 ;
 wire \t$4780 ;
 wire \t$4781 ;
 wire \t$4782 ;
 wire \t$4783 ;
 wire \t$4784 ;
 wire \t$4785 ;
 wire \t$4786 ;
 wire \t$4787 ;
 wire \t$4788 ;
 wire \t$4789 ;
 wire \t$4790 ;
 wire \t$4791 ;
 wire \t$4792 ;
 wire \t$4793 ;
 wire \t$4794 ;
 wire \t$4795 ;
 wire \t$4796 ;
 wire \t$4797 ;
 wire \t$4798 ;
 wire \t$4799 ;
 wire \t$4800 ;
 wire \t$4801 ;
 wire \t$4802 ;
 wire \t$4803 ;
 wire \t$4804 ;
 wire \t$4805 ;
 wire \t$4806 ;
 wire \t$4807 ;
 wire \t$4808 ;
 wire \t$4809 ;
 wire \t$4810 ;
 wire \t$4811 ;
 wire \t$4812 ;
 wire \t$4813 ;
 wire \t$4814 ;
 wire \t$4815 ;
 wire \t$4816 ;
 wire \t$4817 ;
 wire \t$4818 ;
 wire \t$4819 ;
 wire \t$4820 ;
 wire \t$4821 ;
 wire \t$4822 ;
 wire \t$4823 ;
 wire \t$4826 ;
 wire \t$4829 ;
 wire \t$4830 ;
 wire \t$4831 ;
 wire \t$4832 ;
 wire \t$4833 ;
 wire \t$4834 ;
 wire \t$4835 ;
 wire \t$4836 ;
 wire \t$4837 ;
 wire \t$4838 ;
 wire \t$4839 ;
 wire \t$4840 ;
 wire \t$4841 ;
 wire \t$4842 ;
 wire \t$4843 ;
 wire \t$4844 ;
 wire \t$4845 ;
 wire \t$4846 ;
 wire \t$4847 ;
 wire \t$4848 ;
 wire \t$4849 ;
 wire \t$4850 ;
 wire \t$4851 ;
 wire \t$4852 ;
 wire \t$4853 ;
 wire \t$4854 ;
 wire \t$4855 ;
 wire \t$4856 ;
 wire \t$4857 ;
 wire \t$4858 ;
 wire \t$4859 ;
 wire \t$4860 ;
 wire \t$4861 ;
 wire \t$4862 ;
 wire \t$4863 ;
 wire \t$4864 ;
 wire \t$4865 ;
 wire \t$4866 ;
 wire \t$4867 ;
 wire \t$4868 ;
 wire \t$4869 ;
 wire \t$4870 ;
 wire \t$4871 ;
 wire \t$4872 ;
 wire \t$4873 ;
 wire \t$4874 ;
 wire \t$4875 ;
 wire \t$4876 ;
 wire \t$4877 ;
 wire \t$4878 ;
 wire \t$4879 ;
 wire \t$4880 ;
 wire \t$4881 ;
 wire \t$4882 ;
 wire \t$4883 ;
 wire \t$4884 ;
 wire \t$4885 ;
 wire \t$4886 ;
 wire \t$4887 ;
 wire \t$4888 ;
 wire \t$4889 ;
 wire \t$4890 ;
 wire \t$4891 ;
 wire \t$4892 ;
 wire \t$4893 ;
 wire \t$4896 ;
 wire \t$4899 ;
 wire \t$4900 ;
 wire \t$4901 ;
 wire \t$4902 ;
 wire \t$4903 ;
 wire \t$4904 ;
 wire \t$4905 ;
 wire \t$4906 ;
 wire \t$4907 ;
 wire \t$4908 ;
 wire \t$4909 ;
 wire \t$4910 ;
 wire \t$4911 ;
 wire \t$4912 ;
 wire \t$4913 ;
 wire \t$4914 ;
 wire \t$4915 ;
 wire \t$4916 ;
 wire \t$4917 ;
 wire \t$4918 ;
 wire \t$4919 ;
 wire \t$4920 ;
 wire \t$4921 ;
 wire \t$4922 ;
 wire \t$4923 ;
 wire \t$4924 ;
 wire \t$4925 ;
 wire \t$4926 ;
 wire \t$4927 ;
 wire \t$4928 ;
 wire \t$4929 ;
 wire \t$4930 ;
 wire \t$4931 ;
 wire \t$4932 ;
 wire \t$4933 ;
 wire \t$4934 ;
 wire \t$4935 ;
 wire \t$4936 ;
 wire \t$4937 ;
 wire \t$4938 ;
 wire \t$4939 ;
 wire \t$4940 ;
 wire \t$4941 ;
 wire \t$4942 ;
 wire \t$4943 ;
 wire \t$4944 ;
 wire \t$4945 ;
 wire \t$4946 ;
 wire \t$4947 ;
 wire \t$4948 ;
 wire \t$4949 ;
 wire \t$4950 ;
 wire \t$4951 ;
 wire \t$4952 ;
 wire \t$4953 ;
 wire \t$4954 ;
 wire \t$4955 ;
 wire \t$4956 ;
 wire \t$4957 ;
 wire \t$4958 ;
 wire \t$4959 ;
 wire \t$4960 ;
 wire \t$4961 ;
 wire \t$4962 ;
 wire \t$4963 ;
 wire \t$4966 ;
 wire \t$4969 ;
 wire \t$4970 ;
 wire \t$4971 ;
 wire \t$4972 ;
 wire \t$4973 ;
 wire \t$4974 ;
 wire \t$4975 ;
 wire \t$4976 ;
 wire \t$4977 ;
 wire \t$4978 ;
 wire \t$4979 ;
 wire \t$4980 ;
 wire \t$4981 ;
 wire \t$4982 ;
 wire \t$4983 ;
 wire \t$4984 ;
 wire \t$4985 ;
 wire \t$4986 ;
 wire \t$4987 ;
 wire \t$4988 ;
 wire \t$4989 ;
 wire \t$4990 ;
 wire \t$4991 ;
 wire \t$4992 ;
 wire \t$4993 ;
 wire \t$4994 ;
 wire \t$4995 ;
 wire \t$4996 ;
 wire \t$4997 ;
 wire \t$4998 ;
 wire \t$4999 ;
 wire \t$5000 ;
 wire \t$5001 ;
 wire \t$5002 ;
 wire \t$5003 ;
 wire \t$5004 ;
 wire \t$5005 ;
 wire \t$5006 ;
 wire \t$5007 ;
 wire \t$5008 ;
 wire \t$5009 ;
 wire \t$5010 ;
 wire \t$5011 ;
 wire \t$5012 ;
 wire \t$5013 ;
 wire \t$5014 ;
 wire \t$5015 ;
 wire \t$5016 ;
 wire \t$5017 ;
 wire \t$5018 ;
 wire \t$5019 ;
 wire \t$5020 ;
 wire \t$5021 ;
 wire \t$5022 ;
 wire \t$5023 ;
 wire \t$5024 ;
 wire \t$5025 ;
 wire \t$5026 ;
 wire \t$5027 ;
 wire \t$5028 ;
 wire \t$5029 ;
 wire \t$5030 ;
 wire \t$5031 ;
 wire \t$5032 ;
 wire \t$5033 ;
 wire \t$5036 ;
 wire \t$5039 ;
 wire \t$5040 ;
 wire \t$5041 ;
 wire \t$5042 ;
 wire \t$5043 ;
 wire \t$5044 ;
 wire \t$5045 ;
 wire \t$5046 ;
 wire \t$5047 ;
 wire \t$5048 ;
 wire \t$5049 ;
 wire \t$5050 ;
 wire \t$5051 ;
 wire \t$5052 ;
 wire \t$5053 ;
 wire \t$5054 ;
 wire \t$5055 ;
 wire \t$5056 ;
 wire \t$5057 ;
 wire \t$5058 ;
 wire \t$5059 ;
 wire \t$5060 ;
 wire \t$5061 ;
 wire \t$5062 ;
 wire \t$5063 ;
 wire \t$5064 ;
 wire \t$5065 ;
 wire \t$5066 ;
 wire \t$5067 ;
 wire \t$5068 ;
 wire \t$5069 ;
 wire \t$5070 ;
 wire \t$5071 ;
 wire \t$5072 ;
 wire \t$5073 ;
 wire \t$5074 ;
 wire \t$5075 ;
 wire \t$5076 ;
 wire \t$5077 ;
 wire \t$5078 ;
 wire \t$5079 ;
 wire \t$5080 ;
 wire \t$5081 ;
 wire \t$5082 ;
 wire \t$5083 ;
 wire \t$5084 ;
 wire \t$5085 ;
 wire \t$5086 ;
 wire \t$5087 ;
 wire \t$5088 ;
 wire \t$5089 ;
 wire \t$5090 ;
 wire \t$5091 ;
 wire \t$5092 ;
 wire \t$5093 ;
 wire \t$5094 ;
 wire \t$5095 ;
 wire \t$5096 ;
 wire \t$5097 ;
 wire \t$5098 ;
 wire \t$5099 ;
 wire \t$5100 ;
 wire \t$5101 ;
 wire \t$5102 ;
 wire \t$5103 ;
 wire \t$5106 ;
 wire \t$5109 ;
 wire \t$5110 ;
 wire \t$5111 ;
 wire \t$5112 ;
 wire \t$5113 ;
 wire \t$5114 ;
 wire \t$5115 ;
 wire \t$5116 ;
 wire \t$5117 ;
 wire \t$5118 ;
 wire \t$5119 ;
 wire \t$5120 ;
 wire \t$5121 ;
 wire \t$5122 ;
 wire \t$5123 ;
 wire \t$5124 ;
 wire \t$5125 ;
 wire \t$5126 ;
 wire \t$5127 ;
 wire \t$5128 ;
 wire \t$5129 ;
 wire \t$5130 ;
 wire \t$5131 ;
 wire \t$5132 ;
 wire \t$5133 ;
 wire \t$5134 ;
 wire \t$5135 ;
 wire \t$5136 ;
 wire \t$5137 ;
 wire \t$5138 ;
 wire \t$5139 ;
 wire \t$5140 ;
 wire \t$5141 ;
 wire \t$5142 ;
 wire \t$5143 ;
 wire \t$5144 ;
 wire \t$5145 ;
 wire \t$5146 ;
 wire \t$5147 ;
 wire \t$5148 ;
 wire \t$5149 ;
 wire \t$5150 ;
 wire \t$5151 ;
 wire \t$5152 ;
 wire \t$5153 ;
 wire \t$5154 ;
 wire \t$5155 ;
 wire \t$5156 ;
 wire \t$5157 ;
 wire \t$5158 ;
 wire \t$5159 ;
 wire \t$5160 ;
 wire \t$5161 ;
 wire \t$5162 ;
 wire \t$5163 ;
 wire \t$5164 ;
 wire \t$5165 ;
 wire \t$5166 ;
 wire \t$5167 ;
 wire \t$5168 ;
 wire \t$5169 ;
 wire \t$5170 ;
 wire \t$5171 ;
 wire \t$5172 ;
 wire \t$5173 ;
 wire \t$5176 ;
 wire \t$5179 ;
 wire \t$5180 ;
 wire \t$5181 ;
 wire \t$5182 ;
 wire \t$5183 ;
 wire \t$5184 ;
 wire \t$5185 ;
 wire \t$5186 ;
 wire \t$5187 ;
 wire \t$5188 ;
 wire \t$5189 ;
 wire \t$5190 ;
 wire \t$5191 ;
 wire \t$5192 ;
 wire \t$5193 ;
 wire \t$5194 ;
 wire \t$5195 ;
 wire \t$5196 ;
 wire \t$5197 ;
 wire \t$5198 ;
 wire \t$5199 ;
 wire \t$5200 ;
 wire \t$5201 ;
 wire \t$5202 ;
 wire \t$5203 ;
 wire \t$5204 ;
 wire \t$5205 ;
 wire \t$5206 ;
 wire \t$5207 ;
 wire \t$5208 ;
 wire \t$5209 ;
 wire \t$5210 ;
 wire \t$5211 ;
 wire \t$5212 ;
 wire \t$5213 ;
 wire \t$5214 ;
 wire \t$5215 ;
 wire \t$5216 ;
 wire \t$5217 ;
 wire \t$5218 ;
 wire \t$5219 ;
 wire \t$5220 ;
 wire \t$5221 ;
 wire \t$5222 ;
 wire \t$5223 ;
 wire \t$5224 ;
 wire \t$5225 ;
 wire \t$5226 ;
 wire \t$5227 ;
 wire \t$5228 ;
 wire \t$5229 ;
 wire \t$5230 ;
 wire \t$5231 ;
 wire \t$5232 ;
 wire \t$5233 ;
 wire \t$5234 ;
 wire \t$5235 ;
 wire \t$5236 ;
 wire \t$5237 ;
 wire \t$5238 ;
 wire \t$5239 ;
 wire \t$5240 ;
 wire \t$5241 ;
 wire \t$5242 ;
 wire \t$5243 ;
 wire \t$5246 ;
 wire \t$5249 ;
 wire \t$5250 ;
 wire \t$5251 ;
 wire \t$5252 ;
 wire \t$5253 ;
 wire \t$5254 ;
 wire \t$5255 ;
 wire \t$5256 ;
 wire \t$5257 ;
 wire \t$5258 ;
 wire \t$5259 ;
 wire \t$5260 ;
 wire \t$5261 ;
 wire \t$5262 ;
 wire \t$5263 ;
 wire \t$5264 ;
 wire \t$5265 ;
 wire \t$5266 ;
 wire \t$5267 ;
 wire \t$5268 ;
 wire \t$5269 ;
 wire \t$5270 ;
 wire \t$5271 ;
 wire \t$5272 ;
 wire \t$5273 ;
 wire \t$5274 ;
 wire \t$5275 ;
 wire \t$5276 ;
 wire \t$5277 ;
 wire \t$5278 ;
 wire \t$5279 ;
 wire \t$5280 ;
 wire \t$5281 ;
 wire \t$5282 ;
 wire \t$5283 ;
 wire \t$5284 ;
 wire \t$5285 ;
 wire \t$5286 ;
 wire \t$5287 ;
 wire \t$5288 ;
 wire \t$5289 ;
 wire \t$5290 ;
 wire \t$5291 ;
 wire \t$5292 ;
 wire \t$5293 ;
 wire \t$5294 ;
 wire \t$5295 ;
 wire \t$5296 ;
 wire \t$5297 ;
 wire \t$5298 ;
 wire \t$5299 ;
 wire \t$5300 ;
 wire \t$5301 ;
 wire \t$5302 ;
 wire \t$5303 ;
 wire \t$5304 ;
 wire \t$5305 ;
 wire \t$5306 ;
 wire \t$5307 ;
 wire \t$5308 ;
 wire \t$5309 ;
 wire \t$5310 ;
 wire \t$5311 ;
 wire \t$5312 ;
 wire \t$5313 ;
 wire \t$5316 ;
 wire \t$5319 ;
 wire \t$5320 ;
 wire \t$5321 ;
 wire \t$5322 ;
 wire \t$5323 ;
 wire \t$5324 ;
 wire \t$5325 ;
 wire \t$5326 ;
 wire \t$5327 ;
 wire \t$5328 ;
 wire \t$5329 ;
 wire \t$5330 ;
 wire \t$5331 ;
 wire \t$5332 ;
 wire \t$5333 ;
 wire \t$5334 ;
 wire \t$5335 ;
 wire \t$5336 ;
 wire \t$5337 ;
 wire \t$5338 ;
 wire \t$5339 ;
 wire \t$5340 ;
 wire \t$5341 ;
 wire \t$5342 ;
 wire \t$5343 ;
 wire \t$5344 ;
 wire \t$5345 ;
 wire \t$5346 ;
 wire \t$5347 ;
 wire \t$5348 ;
 wire \t$5349 ;
 wire \t$5350 ;
 wire \t$5351 ;
 wire \t$5352 ;
 wire \t$5353 ;
 wire \t$5354 ;
 wire \t$5355 ;
 wire \t$5356 ;
 wire \t$5357 ;
 wire \t$5358 ;
 wire \t$5359 ;
 wire \t$5360 ;
 wire \t$5361 ;
 wire \t$5362 ;
 wire \t$5363 ;
 wire \t$5364 ;
 wire \t$5365 ;
 wire \t$5366 ;
 wire \t$5367 ;
 wire \t$5368 ;
 wire \t$5369 ;
 wire \t$5370 ;
 wire \t$5371 ;
 wire \t$5372 ;
 wire \t$5373 ;
 wire \t$5374 ;
 wire \t$5375 ;
 wire \t$5376 ;
 wire \t$5377 ;
 wire \t$5378 ;
 wire \t$5379 ;
 wire \t$5380 ;
 wire \t$5381 ;
 wire \t$5382 ;
 wire \t$5383 ;
 wire \t$5386 ;
 wire \t$5389 ;
 wire \t$5390 ;
 wire \t$5391 ;
 wire \t$5392 ;
 wire \t$5393 ;
 wire \t$5394 ;
 wire \t$5395 ;
 wire \t$5396 ;
 wire \t$5397 ;
 wire \t$5398 ;
 wire \t$5399 ;
 wire \t$5400 ;
 wire \t$5401 ;
 wire \t$5402 ;
 wire \t$5403 ;
 wire \t$5404 ;
 wire \t$5405 ;
 wire \t$5406 ;
 wire \t$5407 ;
 wire \t$5408 ;
 wire \t$5409 ;
 wire \t$5410 ;
 wire \t$5411 ;
 wire \t$5412 ;
 wire \t$5413 ;
 wire \t$5414 ;
 wire \t$5415 ;
 wire \t$5416 ;
 wire \t$5417 ;
 wire \t$5418 ;
 wire \t$5419 ;
 wire \t$5420 ;
 wire \t$5421 ;
 wire \t$5422 ;
 wire \t$5423 ;
 wire \t$5424 ;
 wire \t$5425 ;
 wire \t$5426 ;
 wire \t$5427 ;
 wire \t$5428 ;
 wire \t$5429 ;
 wire \t$5430 ;
 wire \t$5431 ;
 wire \t$5432 ;
 wire \t$5433 ;
 wire \t$5434 ;
 wire \t$5435 ;
 wire \t$5436 ;
 wire \t$5437 ;
 wire \t$5438 ;
 wire \t$5439 ;
 wire \t$5440 ;
 wire \t$5441 ;
 wire \t$5442 ;
 wire \t$5443 ;
 wire \t$5444 ;
 wire \t$5445 ;
 wire \t$5446 ;
 wire \t$5447 ;
 wire \t$5448 ;
 wire \t$5449 ;
 wire \t$5450 ;
 wire \t$5451 ;
 wire \t$5452 ;
 wire \t$5453 ;
 wire \t$5456 ;
 wire \t$5459 ;
 wire \t$5460 ;
 wire \t$5461 ;
 wire \t$5462 ;
 wire \t$5463 ;
 wire \t$5464 ;
 wire \t$5465 ;
 wire \t$5466 ;
 wire \t$5467 ;
 wire \t$5468 ;
 wire \t$5469 ;
 wire \t$5470 ;
 wire \t$5471 ;
 wire \t$5472 ;
 wire \t$5473 ;
 wire \t$5474 ;
 wire \t$5475 ;
 wire \t$5476 ;
 wire \t$5477 ;
 wire \t$5478 ;
 wire \t$5479 ;
 wire \t$5480 ;
 wire \t$5481 ;
 wire \t$5482 ;
 wire \t$5483 ;
 wire \t$5484 ;
 wire \t$5485 ;
 wire \t$5486 ;
 wire \t$5487 ;
 wire \t$5488 ;
 wire \t$5489 ;
 wire \t$5490 ;
 wire \t$5491 ;
 wire \t$5492 ;
 wire \t$5493 ;
 wire \t$5494 ;
 wire \t$5495 ;
 wire \t$5496 ;
 wire \t$5497 ;
 wire \t$5498 ;
 wire \t$5499 ;
 wire \t$5500 ;
 wire \t$5501 ;
 wire \t$5502 ;
 wire \t$5503 ;
 wire \t$5504 ;
 wire \t$5505 ;
 wire \t$5506 ;
 wire \t$5507 ;
 wire \t$5508 ;
 wire \t$5509 ;
 wire \t$5510 ;
 wire \t$5511 ;
 wire \t$5512 ;
 wire \t$5513 ;
 wire \t$5514 ;
 wire \t$5515 ;
 wire \t$5516 ;
 wire \t$5517 ;
 wire \t$5518 ;
 wire \t$5519 ;
 wire \t$5520 ;
 wire \t$5521 ;
 wire \t$5522 ;
 wire \t$5523 ;
 wire \t$5526 ;
 wire \t$5529 ;
 wire \t$5530 ;
 wire \t$5531 ;
 wire \t$5532 ;
 wire \t$5533 ;
 wire \t$5534 ;
 wire \t$5535 ;
 wire \t$5536 ;
 wire \t$5537 ;
 wire \t$5538 ;
 wire \t$5539 ;
 wire \t$5540 ;
 wire \t$5541 ;
 wire \t$5542 ;
 wire \t$5543 ;
 wire \t$5544 ;
 wire \t$5545 ;
 wire \t$5546 ;
 wire \t$5547 ;
 wire \t$5548 ;
 wire \t$5549 ;
 wire \t$5550 ;
 wire \t$5551 ;
 wire \t$5552 ;
 wire \t$5553 ;
 wire \t$5554 ;
 wire \t$5555 ;
 wire \t$5556 ;
 wire \t$5557 ;
 wire \t$5558 ;
 wire \t$5559 ;
 wire \t$5560 ;
 wire \t$5561 ;
 wire \t$5562 ;
 wire \t$5563 ;
 wire \t$5564 ;
 wire \t$5565 ;
 wire \t$5566 ;
 wire \t$5567 ;
 wire \t$5568 ;
 wire \t$5569 ;
 wire \t$5570 ;
 wire \t$5571 ;
 wire \t$5572 ;
 wire \t$5573 ;
 wire \t$5574 ;
 wire \t$5575 ;
 wire \t$5576 ;
 wire \t$5577 ;
 wire \t$5578 ;
 wire \t$5579 ;
 wire \t$5580 ;
 wire \t$5581 ;
 wire \t$5582 ;
 wire \t$5583 ;
 wire \t$5584 ;
 wire \t$5585 ;
 wire \t$5586 ;
 wire \t$5587 ;
 wire \t$5588 ;
 wire \t$5589 ;
 wire \t$5590 ;
 wire \t$5591 ;
 wire \t$5592 ;
 wire \t$5593 ;
 wire \t$5596 ;
 wire \t$5599 ;
 wire \t$5600 ;
 wire \t$5601 ;
 wire \t$5602 ;
 wire \t$5603 ;
 wire \t$5604 ;
 wire \t$5605 ;
 wire \t$5606 ;
 wire \t$5607 ;
 wire \t$5608 ;
 wire \t$5609 ;
 wire \t$5610 ;
 wire \t$5611 ;
 wire \t$5612 ;
 wire \t$5613 ;
 wire \t$5614 ;
 wire \t$5615 ;
 wire \t$5616 ;
 wire \t$5617 ;
 wire \t$5618 ;
 wire \t$5619 ;
 wire \t$5620 ;
 wire \t$5621 ;
 wire \t$5622 ;
 wire \t$5623 ;
 wire \t$5624 ;
 wire \t$5625 ;
 wire \t$5626 ;
 wire \t$5627 ;
 wire \t$5628 ;
 wire \t$5629 ;
 wire \t$5630 ;
 wire \t$5631 ;
 wire \t$5632 ;
 wire \t$5633 ;
 wire \t$5634 ;
 wire \t$5635 ;
 wire \t$5636 ;
 wire \t$5637 ;
 wire \t$5638 ;
 wire \t$5639 ;
 wire \t$5640 ;
 wire \t$5641 ;
 wire \t$5642 ;
 wire \t$5643 ;
 wire \t$5644 ;
 wire \t$5645 ;
 wire \t$5646 ;
 wire \t$5647 ;
 wire \t$5648 ;
 wire \t$5649 ;
 wire \t$5650 ;
 wire \t$5651 ;
 wire \t$5652 ;
 wire \t$5653 ;
 wire \t$5654 ;
 wire \t$5655 ;
 wire \t$5656 ;
 wire \t$5657 ;
 wire \t$5658 ;
 wire \t$5659 ;
 wire \t$5660 ;
 wire \t$5661 ;
 wire \t$5662 ;
 wire \t$5663 ;
 wire \t$5666 ;
 wire \t$5669 ;
 wire \t$5670 ;
 wire \t$5671 ;
 wire \t$5672 ;
 wire \t$5673 ;
 wire \t$5674 ;
 wire \t$5675 ;
 wire \t$5676 ;
 wire \t$5677 ;
 wire \t$5678 ;
 wire \t$5679 ;
 wire \t$5680 ;
 wire \t$5681 ;
 wire \t$5682 ;
 wire \t$5683 ;
 wire \t$5684 ;
 wire \t$5685 ;
 wire \t$5686 ;
 wire \t$5687 ;
 wire \t$5688 ;
 wire \t$5689 ;
 wire \t$5690 ;
 wire \t$5691 ;
 wire \t$5692 ;
 wire \t$5693 ;
 wire \t$5694 ;
 wire \t$5695 ;
 wire \t$5696 ;
 wire \t$5697 ;
 wire \t$5698 ;
 wire \t$5699 ;
 wire \t$5700 ;
 wire \t$5701 ;
 wire \t$5702 ;
 wire \t$5703 ;
 wire \t$5704 ;
 wire \t$5705 ;
 wire \t$5706 ;
 wire \t$5707 ;
 wire \t$5708 ;
 wire \t$5709 ;
 wire \t$5710 ;
 wire \t$5711 ;
 wire \t$5712 ;
 wire \t$5713 ;
 wire \t$5714 ;
 wire \t$5715 ;
 wire \t$5716 ;
 wire \t$5717 ;
 wire \t$5718 ;
 wire \t$5719 ;
 wire \t$5720 ;
 wire \t$5721 ;
 wire \t$5722 ;
 wire \t$5723 ;
 wire \t$5724 ;
 wire \t$5725 ;
 wire \t$5726 ;
 wire \t$5727 ;
 wire \t$5728 ;
 wire \t$5729 ;
 wire \t$5730 ;
 wire \t$5731 ;
 wire \t$5732 ;
 wire \t$5733 ;
 wire \t$5736 ;
 wire \t$5739 ;
 wire \t$5740 ;
 wire \t$5741 ;
 wire \t$5742 ;
 wire \t$5743 ;
 wire \t$5744 ;
 wire \t$5745 ;
 wire \t$5746 ;
 wire \t$5747 ;
 wire \t$5748 ;
 wire \t$5749 ;
 wire \t$5750 ;
 wire \t$5751 ;
 wire \t$5752 ;
 wire \t$5753 ;
 wire \t$5754 ;
 wire \t$5755 ;
 wire \t$5756 ;
 wire \t$5757 ;
 wire \t$5758 ;
 wire \t$5759 ;
 wire \t$5760 ;
 wire \t$5761 ;
 wire \t$5762 ;
 wire \t$5763 ;
 wire \t$5764 ;
 wire \t$5765 ;
 wire \t$5766 ;
 wire \t$5767 ;
 wire \t$5768 ;
 wire \t$5769 ;
 wire \t$5770 ;
 wire \t$5771 ;
 wire \t$5772 ;
 wire \t$5773 ;
 wire \t$5774 ;
 wire \t$5775 ;
 wire \t$5776 ;
 wire \t$5777 ;
 wire \t$5778 ;
 wire \t$5779 ;
 wire \t$5780 ;
 wire \t$5781 ;
 wire \t$5782 ;
 wire \t$5783 ;
 wire \t$5784 ;
 wire \t$5785 ;
 wire \t$5786 ;
 wire \t$5787 ;
 wire \t$5788 ;
 wire \t$5789 ;
 wire \t$5790 ;
 wire \t$5791 ;
 wire \t$5792 ;
 wire \t$5793 ;
 wire \t$5794 ;
 wire \t$5795 ;
 wire \t$5796 ;
 wire \t$5797 ;
 wire \t$5798 ;
 wire \t$5799 ;
 wire \t$5800 ;
 wire \t$5801 ;
 wire \t$5802 ;
 wire \t$5803 ;
 wire \t$5806 ;
 wire \t$5809 ;
 wire \t$5810 ;
 wire \t$5811 ;
 wire \t$5812 ;
 wire \t$5813 ;
 wire \t$5814 ;
 wire \t$5815 ;
 wire \t$5816 ;
 wire \t$5817 ;
 wire \t$5818 ;
 wire \t$5819 ;
 wire \t$5820 ;
 wire \t$5821 ;
 wire \t$5822 ;
 wire \t$5823 ;
 wire \t$5824 ;
 wire \t$5825 ;
 wire \t$5826 ;
 wire \t$5827 ;
 wire \t$5828 ;
 wire \t$5829 ;
 wire \t$5830 ;
 wire \t$5831 ;
 wire \t$5832 ;
 wire \t$5833 ;
 wire \t$5834 ;
 wire \t$5835 ;
 wire \t$5836 ;
 wire \t$5837 ;
 wire \t$5838 ;
 wire \t$5839 ;
 wire \t$5840 ;
 wire \t$5841 ;
 wire \t$5842 ;
 wire \t$5843 ;
 wire \t$5844 ;
 wire \t$5845 ;
 wire \t$5846 ;
 wire \t$5847 ;
 wire \t$5848 ;
 wire \t$5849 ;
 wire \t$5850 ;
 wire \t$5851 ;
 wire \t$5852 ;
 wire \t$5853 ;
 wire \t$5854 ;
 wire \t$5855 ;
 wire \t$5856 ;
 wire \t$5857 ;
 wire \t$5858 ;
 wire \t$5859 ;
 wire \t$5860 ;
 wire \t$5861 ;
 wire \t$5862 ;
 wire \t$5863 ;
 wire \t$5864 ;
 wire \t$5865 ;
 wire \t$5866 ;
 wire \t$5867 ;
 wire \t$5868 ;
 wire \t$5869 ;
 wire \t$5870 ;
 wire \t$5871 ;
 wire \t$5872 ;
 wire \t$5873 ;
 wire \t$5876 ;
 wire \t$5879 ;
 wire \t$5880 ;
 wire \t$5881 ;
 wire \t$5882 ;
 wire \t$5883 ;
 wire \t$5884 ;
 wire \t$5885 ;
 wire \t$5886 ;
 wire \t$5887 ;
 wire \t$5888 ;
 wire \t$5889 ;
 wire \t$5890 ;
 wire \t$5891 ;
 wire \t$5892 ;
 wire \t$5893 ;
 wire \t$5894 ;
 wire \t$5895 ;
 wire \t$5896 ;
 wire \t$5897 ;
 wire \t$5898 ;
 wire \t$5899 ;
 wire \t$5900 ;
 wire \t$5901 ;
 wire \t$5902 ;
 wire \t$5903 ;
 wire \t$5904 ;
 wire \t$5905 ;
 wire \t$5906 ;
 wire \t$5907 ;
 wire \t$5908 ;
 wire \t$5909 ;
 wire \t$5910 ;
 wire \t$5911 ;
 wire \t$5912 ;
 wire \t$5913 ;
 wire \t$5914 ;
 wire \t$5915 ;
 wire \t$5916 ;
 wire \t$5917 ;
 wire \t$5918 ;
 wire \t$5919 ;
 wire \t$5920 ;
 wire \t$5921 ;
 wire \t$5922 ;
 wire \t$5923 ;
 wire \t$5924 ;
 wire \t$5925 ;
 wire \t$5926 ;
 wire \t$5927 ;
 wire \t$5928 ;
 wire \t$5929 ;
 wire \t$5930 ;
 wire \t$5931 ;
 wire \t$5932 ;
 wire \t$5933 ;
 wire \t$5934 ;
 wire \t$5935 ;
 wire \t$5936 ;
 wire \t$5937 ;
 wire \t$5938 ;
 wire \t$5939 ;
 wire \t$5940 ;
 wire \t$5941 ;
 wire \t$5942 ;
 wire \t$5943 ;
 wire \t$5946 ;
 wire \t$5949 ;
 wire \t$5950 ;
 wire \t$5951 ;
 wire \t$5952 ;
 wire \t$5953 ;
 wire \t$5954 ;
 wire \t$5955 ;
 wire \t$5956 ;
 wire \t$5957 ;
 wire \t$5958 ;
 wire \t$5959 ;
 wire \t$5960 ;
 wire \t$5961 ;
 wire \t$5962 ;
 wire \t$5963 ;
 wire \t$5964 ;
 wire \t$5965 ;
 wire \t$5966 ;
 wire \t$5967 ;
 wire \t$5968 ;
 wire \t$5969 ;
 wire \t$5970 ;
 wire \t$5971 ;
 wire \t$5972 ;
 wire \t$5973 ;
 wire \t$5974 ;
 wire \t$5975 ;
 wire \t$5976 ;
 wire \t$5977 ;
 wire \t$5978 ;
 wire \t$5979 ;
 wire \t$5980 ;
 wire \t$5981 ;
 wire \t$5982 ;
 wire \t$5983 ;
 wire \t$5984 ;
 wire \t$5985 ;
 wire \t$5986 ;
 wire \t$5987 ;
 wire \t$5988 ;
 wire \t$5989 ;
 wire \t$5990 ;
 wire \t$5991 ;
 wire \t$5992 ;
 wire \t$5993 ;
 wire \t$5994 ;
 wire \t$5995 ;
 wire \t$5996 ;
 wire \t$5997 ;
 wire \t$5998 ;
 wire \t$5999 ;
 wire \t$6000 ;
 wire \t$6001 ;
 wire \t$6002 ;
 wire \t$6003 ;
 wire \t$6004 ;
 wire \t$6005 ;
 wire \t$6006 ;
 wire \t$6007 ;
 wire \t$6008 ;
 wire \t$6009 ;
 wire \t$6010 ;
 wire \t$6011 ;
 wire \t$6012 ;
 wire \t$6013 ;
 wire \t$6016 ;
 wire \t$6019 ;
 wire \t$6020 ;
 wire \t$6021 ;
 wire \t$6022 ;
 wire \t$6023 ;
 wire \t$6024 ;
 wire \t$6025 ;
 wire \t$6026 ;
 wire \t$6027 ;
 wire \t$6028 ;
 wire \t$6029 ;
 wire \t$6030 ;
 wire \t$6031 ;
 wire \t$6032 ;
 wire \t$6033 ;
 wire \t$6034 ;
 wire \t$6035 ;
 wire \t$6036 ;
 wire \t$6037 ;
 wire \t$6038 ;
 wire \t$6039 ;
 wire \t$6040 ;
 wire \t$6041 ;
 wire \t$6042 ;
 wire \t$6043 ;
 wire \t$6044 ;
 wire \t$6045 ;
 wire \t$6046 ;
 wire \t$6047 ;
 wire \t$6048 ;
 wire \t$6049 ;
 wire \t$6050 ;
 wire \t$6051 ;
 wire \t$6052 ;
 wire \t$6053 ;
 wire \t$6054 ;
 wire \t$6055 ;
 wire \t$6056 ;
 wire \t$6057 ;
 wire \t$6058 ;
 wire \t$6059 ;
 wire \t$6060 ;
 wire \t$6061 ;
 wire \t$6062 ;
 wire \t$6063 ;
 wire \t$6064 ;
 wire \t$6065 ;
 wire \t$6066 ;
 wire \t$6067 ;
 wire \t$6068 ;
 wire \t$6069 ;
 wire \t$6070 ;
 wire \t$6071 ;
 wire \t$6072 ;
 wire \t$6073 ;
 wire \t$6074 ;
 wire \t$6075 ;
 wire \t$6076 ;
 wire \t$6077 ;
 wire \t$6078 ;
 wire \t$6079 ;
 wire \t$6080 ;
 wire \t$6081 ;
 wire \t$6082 ;
 wire \t$6083 ;
 wire \t$6086 ;
 wire \t$6089 ;
 wire \t$6090 ;
 wire \t$6091 ;
 wire \t$6092 ;
 wire \t$6093 ;
 wire \t$6094 ;
 wire \t$6095 ;
 wire \t$6096 ;
 wire \t$6097 ;
 wire \t$6098 ;
 wire \t$6099 ;
 wire \t$6100 ;
 wire \t$6101 ;
 wire \t$6102 ;
 wire \t$6103 ;
 wire \t$6104 ;
 wire \t$6105 ;
 wire \t$6106 ;
 wire \t$6107 ;
 wire \t$6108 ;
 wire \t$6109 ;
 wire \t$6110 ;
 wire \t$6111 ;
 wire \t$6112 ;
 wire \t$6113 ;
 wire \t$6114 ;
 wire \t$6115 ;
 wire \t$6116 ;
 wire \t$6117 ;
 wire \t$6118 ;
 wire \t$6119 ;
 wire \t$6120 ;
 wire \t$6121 ;
 wire \t$6122 ;
 wire \t$6123 ;
 wire \t$6124 ;
 wire \t$6125 ;
 wire \t$6126 ;
 wire \t$6127 ;
 wire \t$6128 ;
 wire \t$6129 ;
 wire \t$6130 ;
 wire \t$6131 ;
 wire \t$6132 ;
 wire \t$6133 ;
 wire \t$6134 ;
 wire \t$6135 ;
 wire \t$6136 ;
 wire \t$6137 ;
 wire \t$6138 ;
 wire \t$6139 ;
 wire \t$6140 ;
 wire \t$6141 ;
 wire \t$6142 ;
 wire \t$6143 ;
 wire \t$6144 ;
 wire \t$6145 ;
 wire \t$6146 ;
 wire \t$6147 ;
 wire \t$6148 ;
 wire \t$6149 ;
 wire \t$6150 ;
 wire \t$6151 ;
 wire \t$6152 ;
 wire \t$6153 ;
 wire \t$6156 ;
 wire \t$6159 ;
 wire \t$6160 ;
 wire \t$6161 ;
 wire \t$6162 ;
 wire \t$6163 ;
 wire \t$6164 ;
 wire \t$6165 ;
 wire \t$6166 ;
 wire \t$6167 ;
 wire \t$6168 ;
 wire \t$6169 ;
 wire \t$6170 ;
 wire \t$6171 ;
 wire \t$6172 ;
 wire \t$6173 ;
 wire \t$6174 ;
 wire \t$6175 ;
 wire \t$6176 ;
 wire \t$6177 ;
 wire \t$6178 ;
 wire \t$6179 ;
 wire \t$6180 ;
 wire \t$6181 ;
 wire \t$6182 ;
 wire \t$6183 ;
 wire \t$6184 ;
 wire \t$6185 ;
 wire \t$6186 ;
 wire \t$6187 ;
 wire \t$6188 ;
 wire \t$6189 ;
 wire \t$6190 ;
 wire \t$6191 ;
 wire \t$6192 ;
 wire \t$6193 ;
 wire \t$6194 ;
 wire \t$6195 ;
 wire \t$6196 ;
 wire \t$6197 ;
 wire \t$6198 ;
 wire \t$6199 ;
 wire \t$6200 ;
 wire \t$6201 ;
 wire \t$6202 ;
 wire \t$6203 ;
 wire \t$6204 ;
 wire \t$6205 ;
 wire \t$6206 ;
 wire \t$6207 ;
 wire \t$6208 ;
 wire \t$6209 ;
 wire \t$6210 ;
 wire \t$6211 ;
 wire \t$6212 ;
 wire \t$6213 ;
 wire \t$6214 ;
 wire \t$6215 ;
 wire \t$6216 ;
 wire \t$6217 ;
 wire \t$6218 ;
 wire \t$6219 ;
 wire \t$6220 ;
 wire \t$6221 ;
 wire \t$6222 ;
 wire \t$6223 ;
 wire \t$6226 ;
 wire \t$6229 ;
 wire \t$6230 ;
 wire \t$6231 ;
 wire \t$6232 ;
 wire \t$6233 ;
 wire \t$6234 ;
 wire \t$6235 ;
 wire \t$6236 ;
 wire \t$6237 ;
 wire \t$6238 ;
 wire \t$6239 ;
 wire \t$6240 ;
 wire \t$6241 ;
 wire \t$6242 ;
 wire \t$6243 ;
 wire \t$6244 ;
 wire \t$6245 ;
 wire \t$6246 ;
 wire \t$6247 ;
 wire \t$6248 ;
 wire \t$6249 ;
 wire \t$6250 ;
 wire \t$6251 ;
 wire \t$6252 ;
 wire \t$6253 ;
 wire \t$6254 ;
 wire \t$6255 ;
 wire \t$6256 ;
 wire \t$6257 ;
 wire \t$6258 ;
 wire \t$6259 ;
 wire \t$6260 ;
 wire \t$6261 ;
 wire \t$6262 ;
 wire \t$6263 ;
 wire \t$6264 ;
 wire \t$6265 ;
 wire \t$6266 ;
 wire \t$6267 ;
 wire \t$6268 ;
 wire \t$6269 ;
 wire \t$6270 ;
 wire \t$6271 ;
 wire \t$6272 ;
 wire \t$6273 ;
 wire \t$6274 ;
 wire \t$6275 ;
 wire \t$6276 ;
 wire \t$6277 ;
 wire \t$6278 ;
 wire \t$6279 ;
 wire \t$6280 ;
 wire \t$6281 ;
 wire \t$6282 ;
 wire \t$6283 ;
 wire \t$6284 ;
 wire \t$6285 ;
 wire \t$6286 ;
 wire \t$6287 ;
 wire \t$6288 ;
 wire \t$6289 ;
 wire \t$6290 ;
 wire \t$6291 ;
 wire \t$6292 ;
 wire \t$6293 ;
 wire \t$6296 ;
 wire \t$6299 ;
 wire \t$6300 ;
 wire \t$6301 ;
 wire \t$6302 ;
 wire \t$6303 ;
 wire \t$6304 ;
 wire \t$6305 ;
 wire \t$6306 ;
 wire \t$6307 ;
 wire \t$6308 ;
 wire \t$6309 ;
 wire \t$6310 ;
 wire \t$6311 ;
 wire \t$6312 ;
 wire \t$6313 ;
 wire \t$6314 ;
 wire \t$6315 ;
 wire \t$6316 ;
 wire \t$6317 ;
 wire \t$6318 ;
 wire \t$6319 ;
 wire \t$6320 ;
 wire \t$6321 ;
 wire \t$6322 ;
 wire \t$6323 ;
 wire \t$6324 ;
 wire \t$6325 ;
 wire \t$6326 ;
 wire \t$6327 ;
 wire \t$6328 ;
 wire \t$6329 ;
 wire \t$6330 ;
 wire \t$6331 ;
 wire \t$6332 ;
 wire \t$6333 ;
 wire \t$6334 ;
 wire \t$6335 ;
 wire \t$6336 ;
 wire \t$6337 ;
 wire \t$6338 ;
 wire \t$6339 ;
 wire \t$6340 ;
 wire \t$6341 ;
 wire \t$6342 ;
 wire \t$6343 ;
 wire \t$6344 ;
 wire \t$6345 ;
 wire \t$6346 ;
 wire \t$6347 ;
 wire \t$6348 ;
 wire \t$6349 ;
 wire \t$6350 ;
 wire \t$6351 ;
 wire \t$6352 ;
 wire \t$6353 ;
 wire \t$6354 ;
 wire \t$6355 ;
 wire \t$6356 ;
 wire \t$6357 ;
 wire \t$6358 ;
 wire \t$6359 ;
 wire \t$6360 ;
 wire \t$6361 ;
 wire \t$6362 ;
 wire \t$6363 ;
 wire \t$6366 ;
 wire \t$6369 ;
 wire \t$6370 ;
 wire \t$6371 ;
 wire \t$6372 ;
 wire \t$6373 ;
 wire \t$6374 ;
 wire \t$6375 ;
 wire \t$6376 ;
 wire \t$6377 ;
 wire \t$6378 ;
 wire \t$6379 ;
 wire \t$6380 ;
 wire \t$6381 ;
 wire \t$6382 ;
 wire \t$6383 ;
 wire \t$6384 ;
 wire \t$6385 ;
 wire \t$6386 ;
 wire \t$6387 ;
 wire \t$6388 ;
 wire \t$6389 ;
 wire \t$6390 ;
 wire \t$6391 ;
 wire \t$6392 ;
 wire \t$6393 ;
 wire \t$6394 ;
 wire \t$6395 ;
 wire \t$6396 ;
 wire \t$6397 ;
 wire \t$6398 ;
 wire \t$6399 ;
 wire \t$6400 ;
 wire \t$6401 ;
 wire \t$6402 ;
 wire \t$6403 ;
 wire \t$6404 ;
 wire \t$6405 ;
 wire \t$6406 ;
 wire \t$6407 ;
 wire \t$6408 ;
 wire \t$6409 ;
 wire \t$6410 ;
 wire \t$6411 ;
 wire \t$6412 ;
 wire \t$6413 ;
 wire \t$6414 ;
 wire \t$6415 ;
 wire \t$6416 ;
 wire \t$6417 ;
 wire \t$6418 ;
 wire \t$6419 ;
 wire \t$6420 ;
 wire \t$6421 ;
 wire \t$6422 ;
 wire \t$6423 ;
 wire \t$6424 ;
 wire \t$6425 ;
 wire \t$6426 ;
 wire \t$6427 ;
 wire \t$6428 ;
 wire \t$6429 ;
 wire \t$6430 ;
 wire \t$6431 ;
 wire \t$6432 ;
 wire \t$6433 ;
 wire \t$6436 ;
 wire \t$6439 ;
 wire \t$6440 ;
 wire \t$6441 ;
 wire \t$6442 ;
 wire \t$6443 ;
 wire \t$6444 ;
 wire \t$6445 ;
 wire \t$6446 ;
 wire \t$6447 ;
 wire \t$6448 ;
 wire \t$6449 ;
 wire \t$6450 ;
 wire \t$6451 ;
 wire \t$6452 ;
 wire \t$6453 ;
 wire \t$6454 ;
 wire \t$6455 ;
 wire \t$6456 ;
 wire \t$6457 ;
 wire \t$6458 ;
 wire \t$6459 ;
 wire \t$6460 ;
 wire \t$6461 ;
 wire \t$6462 ;
 wire \t$6463 ;
 wire \t$6464 ;
 wire \t$6465 ;
 wire \t$6466 ;
 wire \t$6467 ;
 wire \t$6468 ;
 wire \t$6469 ;
 wire \t$6470 ;
 wire \t$6471 ;
 wire \t$6472 ;
 wire \t$6473 ;
 wire \t$6474 ;
 wire \t$6475 ;
 wire \t$6476 ;
 wire \t$6477 ;
 wire \t$6478 ;
 wire \t$6479 ;
 wire \t$6480 ;
 wire \t$6481 ;
 wire \t$6482 ;
 wire \t$6483 ;
 wire \t$6484 ;
 wire \t$6485 ;
 wire \t$6486 ;
 wire \t$6487 ;
 wire \t$6488 ;
 wire \t$6489 ;
 wire \t$6490 ;
 wire \t$6491 ;
 wire \t$6492 ;
 wire \t$6493 ;
 wire \t$6494 ;
 wire \t$6495 ;
 wire \t$6496 ;
 wire \t$6497 ;
 wire \t$6498 ;
 wire \t$6499 ;
 wire \t$6500 ;
 wire \t$6501 ;
 wire \t$6502 ;
 wire \t$6503 ;
 wire \t$6506 ;
 wire \t$6509 ;
 wire \t$6510 ;
 wire \t$6511 ;
 wire \t$6512 ;
 wire \t$6513 ;
 wire \t$6514 ;
 wire \t$6515 ;
 wire \t$6516 ;
 wire \t$6517 ;
 wire \t$6518 ;
 wire \t$6519 ;
 wire \t$6520 ;
 wire \t$6521 ;
 wire \t$6522 ;
 wire \t$6523 ;
 wire \t$6524 ;
 wire \t$6525 ;
 wire \t$6526 ;
 wire \t$6527 ;
 wire \t$6528 ;
 wire \t$6529 ;
 wire \t$6530 ;
 wire \t$6531 ;
 wire \t$6532 ;
 wire \t$6533 ;
 wire \t$6534 ;
 wire \t$6535 ;
 wire \t$6536 ;
 wire \t$6537 ;
 wire \t$6538 ;
 wire \t$6539 ;
 wire \t$6540 ;
 wire \t$6541 ;
 wire \t$6542 ;
 wire \t$6543 ;
 wire \t$6544 ;
 wire \t$6545 ;
 wire \t$6546 ;
 wire \t$6547 ;
 wire \t$6548 ;
 wire \t$6549 ;
 wire \t$6550 ;
 wire \t$6551 ;
 wire \t$6552 ;
 wire \t$6553 ;
 wire \t$6554 ;
 wire \t$6555 ;
 wire \t$6556 ;
 wire \t$6557 ;
 wire \t$6558 ;
 wire \t$6559 ;
 wire \t$6560 ;
 wire \t$6561 ;
 wire \t$6562 ;
 wire \t$6563 ;
 wire \t$6564 ;
 wire \t$6565 ;
 wire \t$6566 ;
 wire \t$6567 ;
 wire \t$6568 ;
 wire \t$6569 ;
 wire \t$6570 ;
 wire \t$6571 ;
 wire \t$6572 ;
 wire \t$6573 ;
 wire \t$6576 ;
 wire \t$6579 ;
 wire \t$6580 ;
 wire \t$6581 ;
 wire \t$6582 ;
 wire \t$6583 ;
 wire \t$6584 ;
 wire \t$6585 ;
 wire \t$6586 ;
 wire \t$6587 ;
 wire \t$6588 ;
 wire \t$6589 ;
 wire \t$6590 ;
 wire \t$6591 ;
 wire \t$6592 ;
 wire \t$6593 ;
 wire \t$6594 ;
 wire \t$6595 ;
 wire \t$6596 ;
 wire \t$6597 ;
 wire \t$6598 ;
 wire \t$6599 ;
 wire \t$6600 ;
 wire \t$6601 ;
 wire \t$6602 ;
 wire \t$6603 ;
 wire \t$6604 ;
 wire \t$6605 ;
 wire \t$6606 ;
 wire \t$6607 ;
 wire \t$6608 ;
 wire \t$6609 ;
 wire \t$6610 ;
 wire \t$6611 ;
 wire \t$6612 ;
 wire \t$6613 ;
 wire \t$6614 ;
 wire \t$6615 ;
 wire \t$6616 ;
 wire \t$6617 ;
 wire \t$6618 ;
 wire \t$6619 ;
 wire \t$6620 ;
 wire \t$6621 ;
 wire \t$6622 ;
 wire \t$6623 ;
 wire \t$6624 ;
 wire \t$6625 ;
 wire \t$6626 ;
 wire \t$6627 ;
 wire \t$6628 ;
 wire \t$6629 ;
 wire \t$6630 ;
 wire \t$6631 ;
 wire \t$6632 ;
 wire \t$6633 ;
 wire \t$6634 ;
 wire \t$6635 ;
 wire \t$6636 ;
 wire \t$6637 ;
 wire \t$6638 ;
 wire \t$6639 ;
 wire \t$6640 ;
 wire \t$6641 ;
 wire \t$6642 ;
 wire \t$6643 ;
 wire \t$6646 ;
 wire \t$6649 ;
 wire \t$6650 ;
 wire \t$6651 ;
 wire \t$6652 ;
 wire \t$6653 ;
 wire \t$6654 ;
 wire \t$6655 ;
 wire \t$6656 ;
 wire \t$6657 ;
 wire \t$6658 ;
 wire \t$6659 ;
 wire \t$6660 ;
 wire \t$6661 ;
 wire \t$6662 ;
 wire \t$6663 ;
 wire \t$6664 ;
 wire \t$6665 ;
 wire \t$6666 ;
 wire \t$6667 ;
 wire \t$6668 ;
 wire \t$6669 ;
 wire \t$6670 ;
 wire \t$6671 ;
 wire \t$6672 ;
 wire \t$6673 ;
 wire \t$6674 ;
 wire \t$6675 ;
 wire \t$6676 ;
 wire \t$6677 ;
 wire \t$6678 ;
 wire \t$6679 ;
 wire \t$6680 ;
 wire \t$6681 ;
 wire \t$6682 ;
 wire \t$6683 ;
 wire \t$6684 ;
 wire \t$6685 ;
 wire \t$6686 ;
 wire \t$6687 ;
 wire \t$6688 ;
 wire \t$6689 ;
 wire \t$6690 ;
 wire \t$6691 ;
 wire \t$6692 ;
 wire \t$6693 ;
 wire \t$6694 ;
 wire \t$6695 ;
 wire \t$6696 ;
 wire \t$6697 ;
 wire \t$6698 ;
 wire \t$6699 ;
 wire \t$6700 ;
 wire \t$6701 ;
 wire \t$6702 ;
 wire \t$6703 ;
 wire \t$6704 ;
 wire \t$6705 ;
 wire \t$6706 ;
 wire \t$6707 ;
 wire \t$6708 ;
 wire \t$6709 ;
 wire \t$6710 ;
 wire \t$6711 ;
 wire \t$6712 ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sky130_fd_sc_hd__inv_1 \U$$0  (.A(net1753),
    .Y(\notblock[0] ));
 sky130_fd_sc_hd__inv_1 \U$$1  (.A(net1),
    .Y(\notblock[1] ));
 sky130_fd_sc_hd__a22o_1 \U$$10  (.A1(net1127),
    .A2(net447),
    .B1(net1035),
    .B2(net689),
    .X(\t$4412 ));
 sky130_fd_sc_hd__a22o_1 \U$$100  (.A1(net1703),
    .A2(net444),
    .B1(net1695),
    .B2(net686),
    .X(\t$4457 ));
 sky130_fd_sc_hd__xor2_1 \U$$1000  (.A(\t$4916 ),
    .B(net1183),
    .X(booth_b14_m17));
 sky130_fd_sc_hd__a22o_1 \U$$1001  (.A1(net1149),
    .A2(net388),
    .B1(net1143),
    .B2(net654),
    .X(\t$4917 ));
 sky130_fd_sc_hd__xor2_1 \U$$1002  (.A(\t$4917 ),
    .B(net1186),
    .X(booth_b14_m18));
 sky130_fd_sc_hd__a22o_1 \U$$1003  (.A1(net1143),
    .A2(net387),
    .B1(net1133),
    .B2(net653),
    .X(\t$4918 ));
 sky130_fd_sc_hd__xor2_1 \U$$1004  (.A(\t$4918 ),
    .B(net1185),
    .X(booth_b14_m19));
 sky130_fd_sc_hd__a22o_1 \U$$1005  (.A1(net1133),
    .A2(net387),
    .B1(net1117),
    .B2(net653),
    .X(\t$4919 ));
 sky130_fd_sc_hd__xor2_1 \U$$1006  (.A(\t$4919 ),
    .B(net1185),
    .X(booth_b14_m20));
 sky130_fd_sc_hd__a22o_1 \U$$1007  (.A1(net1117),
    .A2(net389),
    .B1(net1108),
    .B2(net655),
    .X(\t$4920 ));
 sky130_fd_sc_hd__xor2_1 \U$$1008  (.A(\t$4920 ),
    .B(net1187),
    .X(booth_b14_m21));
 sky130_fd_sc_hd__a22o_1 \U$$1009  (.A1(net1108),
    .A2(net388),
    .B1(net1100),
    .B2(net654),
    .X(\t$4921 ));
 sky130_fd_sc_hd__xor2_1 \U$$101  (.A(\t$4457 ),
    .B(net1570),
    .X(booth_b0_m47));
 sky130_fd_sc_hd__xor2_1 \U$$1010  (.A(\t$4921 ),
    .B(net1186),
    .X(booth_b14_m22));
 sky130_fd_sc_hd__a22o_1 \U$$1011  (.A1(net1100),
    .A2(net388),
    .B1(net1091),
    .B2(net654),
    .X(\t$4922 ));
 sky130_fd_sc_hd__xor2_1 \U$$1012  (.A(\t$4922 ),
    .B(net1186),
    .X(booth_b14_m23));
 sky130_fd_sc_hd__a22o_1 \U$$1013  (.A1(net1091),
    .A2(net387),
    .B1(net1083),
    .B2(net653),
    .X(\t$4923 ));
 sky130_fd_sc_hd__xor2_1 \U$$1014  (.A(\t$4923 ),
    .B(net1185),
    .X(booth_b14_m24));
 sky130_fd_sc_hd__a22o_1 \U$$1015  (.A1(net1081),
    .A2(net387),
    .B1(net1072),
    .B2(net653),
    .X(\t$4924 ));
 sky130_fd_sc_hd__xor2_1 \U$$1016  (.A(\t$4924 ),
    .B(net1185),
    .X(booth_b14_m25));
 sky130_fd_sc_hd__a22o_1 \U$$1017  (.A1(net1071),
    .A2(net386),
    .B1(net1063),
    .B2(net652),
    .X(\t$4925 ));
 sky130_fd_sc_hd__xor2_1 \U$$1018  (.A(\t$4925 ),
    .B(net1183),
    .X(booth_b14_m26));
 sky130_fd_sc_hd__a22o_1 \U$$1019  (.A1(net1063),
    .A2(net386),
    .B1(net1055),
    .B2(net652),
    .X(\t$4926 ));
 sky130_fd_sc_hd__a22o_1 \U$$102  (.A1(net1695),
    .A2(net444),
    .B1(net1687),
    .B2(net686),
    .X(\t$4458 ));
 sky130_fd_sc_hd__xor2_1 \U$$1020  (.A(\t$4926 ),
    .B(net1184),
    .X(booth_b14_m27));
 sky130_fd_sc_hd__a22o_1 \U$$1021  (.A1(net1055),
    .A2(net386),
    .B1(net1047),
    .B2(net652),
    .X(\t$4927 ));
 sky130_fd_sc_hd__xor2_1 \U$$1022  (.A(\t$4927 ),
    .B(net1184),
    .X(booth_b14_m28));
 sky130_fd_sc_hd__a22o_1 \U$$1023  (.A1(net1047),
    .A2(net386),
    .B1(net1039),
    .B2(net652),
    .X(\t$4928 ));
 sky130_fd_sc_hd__xor2_1 \U$$1024  (.A(\t$4928 ),
    .B(net1184),
    .X(booth_b14_m29));
 sky130_fd_sc_hd__a22o_1 \U$$1025  (.A1(net1039),
    .A2(net386),
    .B1(net1023),
    .B2(net652),
    .X(\t$4929 ));
 sky130_fd_sc_hd__xor2_1 \U$$1026  (.A(\t$4929 ),
    .B(net1184),
    .X(booth_b14_m30));
 sky130_fd_sc_hd__a22o_1 \U$$1027  (.A1(net1023),
    .A2(net388),
    .B1(net1015),
    .B2(net654),
    .X(\t$4930 ));
 sky130_fd_sc_hd__xor2_1 \U$$1028  (.A(\t$4930 ),
    .B(net1186),
    .X(booth_b14_m31));
 sky130_fd_sc_hd__a22o_1 \U$$1029  (.A1(net1015),
    .A2(net386),
    .B1(net998),
    .B2(net652),
    .X(\t$4931 ));
 sky130_fd_sc_hd__xor2_1 \U$$103  (.A(\t$4458 ),
    .B(net1570),
    .X(booth_b0_m48));
 sky130_fd_sc_hd__xor2_1 \U$$1030  (.A(\t$4931 ),
    .B(net1184),
    .X(booth_b14_m32));
 sky130_fd_sc_hd__a22o_1 \U$$1031  (.A1(net998),
    .A2(net386),
    .B1(net990),
    .B2(net652),
    .X(\t$4932 ));
 sky130_fd_sc_hd__xor2_1 \U$$1032  (.A(\t$4932 ),
    .B(net1184),
    .X(booth_b14_m33));
 sky130_fd_sc_hd__a22o_1 \U$$1033  (.A1(net990),
    .A2(net386),
    .B1(net982),
    .B2(net652),
    .X(\t$4933 ));
 sky130_fd_sc_hd__xor2_1 \U$$1034  (.A(\t$4933 ),
    .B(net1184),
    .X(booth_b14_m34));
 sky130_fd_sc_hd__a22o_1 \U$$1035  (.A1(net983),
    .A2(net390),
    .B1(net974),
    .B2(net656),
    .X(\t$4934 ));
 sky130_fd_sc_hd__xor2_1 \U$$1036  (.A(\t$4934 ),
    .B(net1184),
    .X(booth_b14_m35));
 sky130_fd_sc_hd__a22o_1 \U$$1037  (.A1(net977),
    .A2(net388),
    .B1(net969),
    .B2(net654),
    .X(\t$4935 ));
 sky130_fd_sc_hd__xor2_1 \U$$1038  (.A(\t$4935 ),
    .B(net1186),
    .X(booth_b14_m36));
 sky130_fd_sc_hd__a22o_1 \U$$1039  (.A1(net969),
    .A2(net389),
    .B1(net961),
    .B2(net655),
    .X(\t$4936 ));
 sky130_fd_sc_hd__a22o_1 \U$$104  (.A1(net1690),
    .A2(net449),
    .B1(net1682),
    .B2(net691),
    .X(\t$4459 ));
 sky130_fd_sc_hd__xor2_1 \U$$1040  (.A(\t$4936 ),
    .B(net1186),
    .X(booth_b14_m37));
 sky130_fd_sc_hd__a22o_1 \U$$1041  (.A1(net961),
    .A2(net388),
    .B1(net955),
    .B2(net654),
    .X(\t$4937 ));
 sky130_fd_sc_hd__xor2_1 \U$$1042  (.A(\t$4937 ),
    .B(net1186),
    .X(booth_b14_m38));
 sky130_fd_sc_hd__a22o_1 \U$$1043  (.A1(net955),
    .A2(net388),
    .B1(net944),
    .B2(net654),
    .X(\t$4938 ));
 sky130_fd_sc_hd__xor2_1 \U$$1044  (.A(\t$4938 ),
    .B(net1186),
    .X(booth_b14_m39));
 sky130_fd_sc_hd__a22o_1 \U$$1045  (.A1(net944),
    .A2(net388),
    .B1(net928),
    .B2(net654),
    .X(\t$4939 ));
 sky130_fd_sc_hd__xor2_1 \U$$1046  (.A(\t$4939 ),
    .B(net1186),
    .X(booth_b14_m40));
 sky130_fd_sc_hd__a22o_1 \U$$1047  (.A1(net928),
    .A2(net388),
    .B1(net1749),
    .B2(net654),
    .X(\t$4940 ));
 sky130_fd_sc_hd__xor2_1 \U$$1048  (.A(\t$4940 ),
    .B(net1186),
    .X(booth_b14_m41));
 sky130_fd_sc_hd__a22o_1 \U$$1049  (.A1(net1749),
    .A2(net392),
    .B1(net1741),
    .B2(net658),
    .X(\t$4941 ));
 sky130_fd_sc_hd__xor2_1 \U$$105  (.A(\t$4459 ),
    .B(net1576),
    .X(booth_b0_m49));
 sky130_fd_sc_hd__xor2_1 \U$$1050  (.A(\t$4941 ),
    .B(net1187),
    .X(booth_b14_m42));
 sky130_fd_sc_hd__a22o_1 \U$$1051  (.A1(net1741),
    .A2(net388),
    .B1(net1733),
    .B2(net654),
    .X(\t$4942 ));
 sky130_fd_sc_hd__xor2_1 \U$$1052  (.A(\t$4942 ),
    .B(net1187),
    .X(booth_b14_m43));
 sky130_fd_sc_hd__a22o_1 \U$$1053  (.A1(net1733),
    .A2(net391),
    .B1(net1724),
    .B2(net657),
    .X(\t$4943 ));
 sky130_fd_sc_hd__xor2_1 \U$$1054  (.A(\t$4943 ),
    .B(net1187),
    .X(booth_b14_m44));
 sky130_fd_sc_hd__a22o_1 \U$$1055  (.A1(net1720),
    .A2(net390),
    .B1(net1711),
    .B2(net656),
    .X(\t$4944 ));
 sky130_fd_sc_hd__xor2_1 \U$$1056  (.A(\t$4944 ),
    .B(net1190),
    .X(booth_b14_m45));
 sky130_fd_sc_hd__a22o_1 \U$$1057  (.A1(net1711),
    .A2(net390),
    .B1(net1703),
    .B2(net656),
    .X(\t$4945 ));
 sky130_fd_sc_hd__xor2_1 \U$$1058  (.A(\t$4945 ),
    .B(net1190),
    .X(booth_b14_m46));
 sky130_fd_sc_hd__a22o_1 \U$$1059  (.A1(net1703),
    .A2(net390),
    .B1(net1695),
    .B2(net656),
    .X(\t$4946 ));
 sky130_fd_sc_hd__a22o_1 \U$$106  (.A1(net1679),
    .A2(net445),
    .B1(net1654),
    .B2(net687),
    .X(\t$4460 ));
 sky130_fd_sc_hd__xor2_1 \U$$1060  (.A(\t$4946 ),
    .B(net1190),
    .X(booth_b14_m47));
 sky130_fd_sc_hd__a22o_1 \U$$1061  (.A1(net1695),
    .A2(net390),
    .B1(net1687),
    .B2(net656),
    .X(\t$4947 ));
 sky130_fd_sc_hd__xor2_1 \U$$1062  (.A(\t$4947 ),
    .B(net1190),
    .X(booth_b14_m48));
 sky130_fd_sc_hd__a22o_1 \U$$1063  (.A1(net1687),
    .A2(net390),
    .B1(net1679),
    .B2(net656),
    .X(\t$4948 ));
 sky130_fd_sc_hd__xor2_1 \U$$1064  (.A(\t$4948 ),
    .B(net1190),
    .X(booth_b14_m49));
 sky130_fd_sc_hd__a22o_1 \U$$1065  (.A1(net1682),
    .A2(net391),
    .B1(net1657),
    .B2(net657),
    .X(\t$4949 ));
 sky130_fd_sc_hd__xor2_1 \U$$1066  (.A(\t$4949 ),
    .B(net1191),
    .X(booth_b14_m50));
 sky130_fd_sc_hd__a22o_1 \U$$1067  (.A1(net1657),
    .A2(net391),
    .B1(net1649),
    .B2(net657),
    .X(\t$4950 ));
 sky130_fd_sc_hd__xor2_1 \U$$1068  (.A(\t$4950 ),
    .B(net1191),
    .X(booth_b14_m51));
 sky130_fd_sc_hd__a22o_1 \U$$1069  (.A1(net1649),
    .A2(net391),
    .B1(net1641),
    .B2(net657),
    .X(\t$4951 ));
 sky130_fd_sc_hd__xor2_1 \U$$107  (.A(\t$4460 ),
    .B(net1570),
    .X(booth_b0_m50));
 sky130_fd_sc_hd__xor2_1 \U$$1070  (.A(\t$4951 ),
    .B(net1191),
    .X(booth_b14_m52));
 sky130_fd_sc_hd__a22o_1 \U$$1071  (.A1(net1641),
    .A2(net392),
    .B1(net1633),
    .B2(net658),
    .X(\t$4952 ));
 sky130_fd_sc_hd__xor2_1 \U$$1072  (.A(\t$4952 ),
    .B(net1191),
    .X(booth_b14_m53));
 sky130_fd_sc_hd__a22o_1 \U$$1073  (.A1(net1633),
    .A2(net392),
    .B1(net1623),
    .B2(net658),
    .X(\t$4953 ));
 sky130_fd_sc_hd__xor2_1 \U$$1074  (.A(\t$4953 ),
    .B(net1191),
    .X(booth_b14_m54));
 sky130_fd_sc_hd__a22o_1 \U$$1075  (.A1(net1623),
    .A2(net391),
    .B1(net1615),
    .B2(net657),
    .X(\t$4954 ));
 sky130_fd_sc_hd__xor2_1 \U$$1076  (.A(\t$4954 ),
    .B(net1191),
    .X(booth_b14_m55));
 sky130_fd_sc_hd__a22o_1 \U$$1077  (.A1(net1615),
    .A2(net392),
    .B1(net1607),
    .B2(net658),
    .X(\t$4955 ));
 sky130_fd_sc_hd__xor2_1 \U$$1078  (.A(\t$4955 ),
    .B(net1191),
    .X(booth_b14_m56));
 sky130_fd_sc_hd__a22o_1 \U$$1079  (.A1(net1604),
    .A2(net390),
    .B1(net1595),
    .B2(net656),
    .X(\t$4956 ));
 sky130_fd_sc_hd__a22o_1 \U$$108  (.A1(net1658),
    .A2(net449),
    .B1(net1649),
    .B2(net691),
    .X(\t$4461 ));
 sky130_fd_sc_hd__xor2_1 \U$$1080  (.A(\t$4956 ),
    .B(net1188),
    .X(booth_b14_m57));
 sky130_fd_sc_hd__a22o_1 \U$$1081  (.A1(net1596),
    .A2(net390),
    .B1(net1587),
    .B2(net656),
    .X(\t$4957 ));
 sky130_fd_sc_hd__xor2_1 \U$$1082  (.A(\t$4957 ),
    .B(net1189),
    .X(booth_b14_m58));
 sky130_fd_sc_hd__a22o_1 \U$$1083  (.A1(net1586),
    .A2(net390),
    .B1(net1578),
    .B2(net656),
    .X(\t$4958 ));
 sky130_fd_sc_hd__xor2_1 \U$$1084  (.A(\t$4958 ),
    .B(net1188),
    .X(booth_b14_m59));
 sky130_fd_sc_hd__a22o_1 \U$$1085  (.A1(net1578),
    .A2(net391),
    .B1(net1551),
    .B2(net657),
    .X(\t$4959 ));
 sky130_fd_sc_hd__xor2_1 \U$$1086  (.A(\t$4959 ),
    .B(net1188),
    .X(booth_b14_m60));
 sky130_fd_sc_hd__a22o_1 \U$$1087  (.A1(net1551),
    .A2(net391),
    .B1(net1543),
    .B2(net657),
    .X(\t$4960 ));
 sky130_fd_sc_hd__xor2_1 \U$$1088  (.A(\t$4960 ),
    .B(net1188),
    .X(booth_b14_m61));
 sky130_fd_sc_hd__a22o_1 \U$$1089  (.A1(net1543),
    .A2(net391),
    .B1(net1535),
    .B2(net657),
    .X(\t$4961 ));
 sky130_fd_sc_hd__xor2_1 \U$$109  (.A(\t$4461 ),
    .B(net1576),
    .X(booth_b0_m51));
 sky130_fd_sc_hd__xor2_1 \U$$1090  (.A(\t$4961 ),
    .B(net1188),
    .X(booth_b14_m62));
 sky130_fd_sc_hd__a22o_1 \U$$1091  (.A1(net1535),
    .A2(net391),
    .B1(net1527),
    .B2(net657),
    .X(\t$4962 ));
 sky130_fd_sc_hd__xor2_1 \U$$1092  (.A(\t$4962 ),
    .B(net1188),
    .X(booth_b14_m63));
 sky130_fd_sc_hd__a22o_1 \U$$1093  (.A1(net1530),
    .A2(net390),
    .B1(net1754),
    .B2(net656),
    .X(\t$4963 ));
 sky130_fd_sc_hd__xor2_1 \U$$1094  (.A(\t$4963 ),
    .B(net1189),
    .X(booth_b14_m64));
 sky130_fd_sc_hd__inv_1 \U$$1095  (.A(net1188),
    .Y(\notsign$4964 ));
 sky130_fd_sc_hd__inv_1 \U$$1096  (.A(net1188),
    .Y(\notblock$4965[0] ));
 sky130_fd_sc_hd__inv_1 \U$$1097  (.A(net8),
    .Y(\notblock$4965[1] ));
 sky130_fd_sc_hd__inv_1 \U$$1098  (.A(net1012),
    .Y(\notblock$4965[2] ));
 sky130_fd_sc_hd__and2_1 \U$$1099  (.A(net1012),
    .B(\notblock$4965[1] ),
    .X(\t$4966 ));
 sky130_fd_sc_hd__xor2_1 \U$$11  (.A(\t$4412 ),
    .B(net1573),
    .X(booth_b0_m2));
 sky130_fd_sc_hd__a22o_1 \U$$110  (.A1(net1650),
    .A2(net449),
    .B1(net1641),
    .B2(net691),
    .X(\t$4462 ));
 sky130_fd_sc_hd__a32o_2 \U$$1100  (.A1(\notblock$4965[2] ),
    .A2(net8),
    .A3(net1188),
    .B1(\t$4966 ),
    .B2(\notblock$4965[0] ),
    .X(\sel_0$4967 ));
 sky130_fd_sc_hd__xor2_4 \U$$1101  (.A(net8),
    .B(net1188),
    .X(\sel_1$4968 ));
 sky130_fd_sc_hd__a22o_1 \U$$1102  (.A1(net1755),
    .A2(net643),
    .B1(net1228),
    .B2(net916),
    .X(\t$4969 ));
 sky130_fd_sc_hd__xor2_1 \U$$1103  (.A(\t$4969 ),
    .B(net1006),
    .X(booth_b16_m0));
 sky130_fd_sc_hd__a22o_1 \U$$1104  (.A1(net1228),
    .A2(net644),
    .B1(net1123),
    .B2(net917),
    .X(\t$4970 ));
 sky130_fd_sc_hd__xor2_1 \U$$1105  (.A(\t$4970 ),
    .B(net1006),
    .X(booth_b16_m1));
 sky130_fd_sc_hd__a22o_1 \U$$1106  (.A1(net1123),
    .A2(net646),
    .B1(net1032),
    .B2(net919),
    .X(\t$4971 ));
 sky130_fd_sc_hd__xor2_1 \U$$1107  (.A(\t$4971 ),
    .B(net1009),
    .X(booth_b16_m2));
 sky130_fd_sc_hd__a22o_1 \U$$1108  (.A1(net1032),
    .A2(net646),
    .B1(net933),
    .B2(net919),
    .X(\t$4972 ));
 sky130_fd_sc_hd__xor2_1 \U$$1109  (.A(\t$4972 ),
    .B(net1009),
    .X(booth_b16_m3));
 sky130_fd_sc_hd__xor2_1 \U$$111  (.A(\t$4462 ),
    .B(net1576),
    .X(booth_b0_m52));
 sky130_fd_sc_hd__a22o_1 \U$$1110  (.A1(net936),
    .A2(net646),
    .B1(net1676),
    .B2(net919),
    .X(\t$4973 ));
 sky130_fd_sc_hd__xor2_1 \U$$1111  (.A(\t$4973 ),
    .B(net1009),
    .X(booth_b16_m4));
 sky130_fd_sc_hd__a22o_1 \U$$1112  (.A1(net1676),
    .A2(net646),
    .B1(net1564),
    .B2(net919),
    .X(\t$4974 ));
 sky130_fd_sc_hd__xor2_1 \U$$1113  (.A(\t$4974 ),
    .B(net1009),
    .X(booth_b16_m5));
 sky130_fd_sc_hd__a22o_1 \U$$1114  (.A1(net1564),
    .A2(net646),
    .B1(net1523),
    .B2(net919),
    .X(\t$4975 ));
 sky130_fd_sc_hd__xor2_1 \U$$1115  (.A(\t$4975 ),
    .B(net1009),
    .X(booth_b16_m6));
 sky130_fd_sc_hd__a22o_1 \U$$1116  (.A1(net1521),
    .A2(net646),
    .B1(net1513),
    .B2(net919),
    .X(\t$4976 ));
 sky130_fd_sc_hd__xor2_1 \U$$1117  (.A(\t$4976 ),
    .B(net1009),
    .X(booth_b16_m7));
 sky130_fd_sc_hd__a22o_1 \U$$1118  (.A1(net1513),
    .A2(net643),
    .B1(net1505),
    .B2(net916),
    .X(\t$4977 ));
 sky130_fd_sc_hd__xor2_1 \U$$1119  (.A(\t$4977 ),
    .B(net1006),
    .X(booth_b16_m8));
 sky130_fd_sc_hd__a22o_1 \U$$112  (.A1(net1642),
    .A2(net449),
    .B1(net1633),
    .B2(net691),
    .X(\t$4463 ));
 sky130_fd_sc_hd__a22o_1 \U$$1120  (.A1(net1505),
    .A2(net644),
    .B1(net1496),
    .B2(net917),
    .X(\t$4978 ));
 sky130_fd_sc_hd__xor2_1 \U$$1121  (.A(\t$4978 ),
    .B(net1008),
    .X(booth_b16_m9));
 sky130_fd_sc_hd__a22o_1 \U$$1122  (.A1(net1494),
    .A2(net643),
    .B1(net1219),
    .B2(net916),
    .X(\t$4979 ));
 sky130_fd_sc_hd__xor2_1 \U$$1123  (.A(\t$4979 ),
    .B(net1008),
    .X(booth_b16_m10));
 sky130_fd_sc_hd__a22o_1 \U$$1124  (.A1(net1219),
    .A2(net643),
    .B1(net1210),
    .B2(net916),
    .X(\t$4980 ));
 sky130_fd_sc_hd__xor2_1 \U$$1125  (.A(\t$4980 ),
    .B(net1006),
    .X(booth_b16_m11));
 sky130_fd_sc_hd__a22o_1 \U$$1126  (.A1(net1210),
    .A2(net643),
    .B1(net1201),
    .B2(net916),
    .X(\t$4981 ));
 sky130_fd_sc_hd__xor2_1 \U$$1127  (.A(\t$4981 ),
    .B(net1006),
    .X(booth_b16_m12));
 sky130_fd_sc_hd__a22o_1 \U$$1128  (.A1(net1201),
    .A2(net643),
    .B1(net1192),
    .B2(net916),
    .X(\t$4982 ));
 sky130_fd_sc_hd__xor2_1 \U$$1129  (.A(\t$4982 ),
    .B(net1006),
    .X(booth_b16_m13));
 sky130_fd_sc_hd__xor2_1 \U$$113  (.A(\t$4463 ),
    .B(net1576),
    .X(booth_b0_m53));
 sky130_fd_sc_hd__a22o_1 \U$$1130  (.A1(net1192),
    .A2(net643),
    .B1(net1173),
    .B2(net916),
    .X(\t$4983 ));
 sky130_fd_sc_hd__xor2_1 \U$$1131  (.A(\t$4983 ),
    .B(net1006),
    .X(booth_b16_m14));
 sky130_fd_sc_hd__a22o_1 \U$$1132  (.A1(net1173),
    .A2(net643),
    .B1(net1164),
    .B2(net916),
    .X(\t$4984 ));
 sky130_fd_sc_hd__xor2_1 \U$$1133  (.A(\t$4984 ),
    .B(net1006),
    .X(booth_b16_m15));
 sky130_fd_sc_hd__a22o_1 \U$$1134  (.A1(net1166),
    .A2(net645),
    .B1(net1157),
    .B2(net918),
    .X(\t$4985 ));
 sky130_fd_sc_hd__xor2_1 \U$$1135  (.A(\t$4985 ),
    .B(net1010),
    .X(booth_b16_m16));
 sky130_fd_sc_hd__a22o_1 \U$$1136  (.A1(net1161),
    .A2(net646),
    .B1(net1149),
    .B2(net919),
    .X(\t$4986 ));
 sky130_fd_sc_hd__xor2_1 \U$$1137  (.A(\t$4986 ),
    .B(net1009),
    .X(booth_b16_m17));
 sky130_fd_sc_hd__a22o_1 \U$$1138  (.A1(net1149),
    .A2(net646),
    .B1(net1143),
    .B2(net919),
    .X(\t$4987 ));
 sky130_fd_sc_hd__xor2_1 \U$$1139  (.A(\t$4987 ),
    .B(net1010),
    .X(booth_b16_m18));
 sky130_fd_sc_hd__a22o_1 \U$$114  (.A1(net1633),
    .A2(net449),
    .B1(net1623),
    .B2(net691),
    .X(\t$4464 ));
 sky130_fd_sc_hd__a22o_1 \U$$1140  (.A1(net1144),
    .A2(net647),
    .B1(net1133),
    .B2(net920),
    .X(\t$4988 ));
 sky130_fd_sc_hd__xor2_1 \U$$1141  (.A(\t$4988 ),
    .B(net1010),
    .X(booth_b16_m19));
 sky130_fd_sc_hd__a22o_1 \U$$1142  (.A1(net1133),
    .A2(net645),
    .B1(net1117),
    .B2(net918),
    .X(\t$4989 ));
 sky130_fd_sc_hd__xor2_1 \U$$1143  (.A(\t$4989 ),
    .B(net1009),
    .X(booth_b16_m20));
 sky130_fd_sc_hd__a22o_1 \U$$1144  (.A1(net1115),
    .A2(net645),
    .B1(net1106),
    .B2(net918),
    .X(\t$4990 ));
 sky130_fd_sc_hd__xor2_1 \U$$1145  (.A(\t$4990 ),
    .B(net1009),
    .X(booth_b16_m21));
 sky130_fd_sc_hd__a22o_1 \U$$1146  (.A1(net1106),
    .A2(net646),
    .B1(net1100),
    .B2(net919),
    .X(\t$4991 ));
 sky130_fd_sc_hd__xor2_1 \U$$1147  (.A(\t$4991 ),
    .B(net1009),
    .X(booth_b16_m22));
 sky130_fd_sc_hd__a22o_1 \U$$1148  (.A1(net1099),
    .A2(net643),
    .B1(net1089),
    .B2(net916),
    .X(\t$4992 ));
 sky130_fd_sc_hd__xor2_1 \U$$1149  (.A(\t$4992 ),
    .B(net1008),
    .X(booth_b16_m23));
 sky130_fd_sc_hd__xor2_1 \U$$115  (.A(\t$4464 ),
    .B(net1576),
    .X(booth_b0_m54));
 sky130_fd_sc_hd__a22o_1 \U$$1150  (.A1(net1088),
    .A2(net643),
    .B1(net1080),
    .B2(net916),
    .X(\t$4993 ));
 sky130_fd_sc_hd__xor2_1 \U$$1151  (.A(\t$4993 ),
    .B(net1006),
    .X(booth_b16_m24));
 sky130_fd_sc_hd__a22o_1 \U$$1152  (.A1(net1080),
    .A2(net644),
    .B1(net1071),
    .B2(net917),
    .X(\t$4994 ));
 sky130_fd_sc_hd__xor2_1 \U$$1153  (.A(\t$4994 ),
    .B(net1007),
    .X(booth_b16_m25));
 sky130_fd_sc_hd__a22o_1 \U$$1154  (.A1(net1071),
    .A2(net644),
    .B1(net1063),
    .B2(net917),
    .X(\t$4995 ));
 sky130_fd_sc_hd__xor2_1 \U$$1155  (.A(\t$4995 ),
    .B(net1006),
    .X(booth_b16_m26));
 sky130_fd_sc_hd__a22o_1 \U$$1156  (.A1(net1064),
    .A2(net648),
    .B1(net1056),
    .B2(net921),
    .X(\t$4996 ));
 sky130_fd_sc_hd__xor2_1 \U$$1157  (.A(\t$4996 ),
    .B(net1007),
    .X(booth_b16_m27));
 sky130_fd_sc_hd__a22o_1 \U$$1158  (.A1(net1055),
    .A2(net647),
    .B1(net1047),
    .B2(net920),
    .X(\t$4997 ));
 sky130_fd_sc_hd__xor2_1 \U$$1159  (.A(\t$4997 ),
    .B(net1007),
    .X(booth_b16_m28));
 sky130_fd_sc_hd__a22o_1 \U$$116  (.A1(net1623),
    .A2(net449),
    .B1(net1619),
    .B2(net691),
    .X(\t$4465 ));
 sky130_fd_sc_hd__a22o_1 \U$$1160  (.A1(net1047),
    .A2(net644),
    .B1(net1039),
    .B2(net917),
    .X(\t$4998 ));
 sky130_fd_sc_hd__xor2_1 \U$$1161  (.A(\t$4998 ),
    .B(net1007),
    .X(booth_b16_m29));
 sky130_fd_sc_hd__a22o_1 \U$$1162  (.A1(net1039),
    .A2(net644),
    .B1(net1023),
    .B2(net917),
    .X(\t$4999 ));
 sky130_fd_sc_hd__xor2_1 \U$$1163  (.A(\t$4999 ),
    .B(net1007),
    .X(booth_b16_m30));
 sky130_fd_sc_hd__a22o_1 \U$$1164  (.A1(net1023),
    .A2(net644),
    .B1(net1015),
    .B2(net917),
    .X(\t$5000 ));
 sky130_fd_sc_hd__xor2_1 \U$$1165  (.A(\t$5000 ),
    .B(net1007),
    .X(booth_b16_m31));
 sky130_fd_sc_hd__a22o_1 \U$$1166  (.A1(net1015),
    .A2(net644),
    .B1(net998),
    .B2(net917),
    .X(\t$5001 ));
 sky130_fd_sc_hd__xor2_1 \U$$1167  (.A(\t$5001 ),
    .B(net1007),
    .X(booth_b16_m32));
 sky130_fd_sc_hd__a22o_1 \U$$1168  (.A1(net999),
    .A2(net644),
    .B1(net991),
    .B2(net917),
    .X(\t$5002 ));
 sky130_fd_sc_hd__xor2_1 \U$$1169  (.A(\t$5002 ),
    .B(net1007),
    .X(booth_b16_m33));
 sky130_fd_sc_hd__xor2_1 \U$$117  (.A(\t$4465 ),
    .B(net1576),
    .X(booth_b0_m55));
 sky130_fd_sc_hd__a22o_1 \U$$1170  (.A1(net990),
    .A2(net645),
    .B1(net983),
    .B2(net918),
    .X(\t$5003 ));
 sky130_fd_sc_hd__xor2_1 \U$$1171  (.A(\t$5003 ),
    .B(net1010),
    .X(booth_b16_m34));
 sky130_fd_sc_hd__a22o_1 \U$$1172  (.A1(net987),
    .A2(net647),
    .B1(net977),
    .B2(net920),
    .X(\t$5004 ));
 sky130_fd_sc_hd__xor2_1 \U$$1173  (.A(\t$5004 ),
    .B(net1010),
    .X(booth_b16_m35));
 sky130_fd_sc_hd__a22o_1 \U$$1174  (.A1(net977),
    .A2(net645),
    .B1(net969),
    .B2(net918),
    .X(\t$5005 ));
 sky130_fd_sc_hd__xor2_1 \U$$1175  (.A(\t$5005 ),
    .B(net1010),
    .X(booth_b16_m36));
 sky130_fd_sc_hd__a22o_1 \U$$1176  (.A1(net969),
    .A2(net647),
    .B1(net961),
    .B2(net920),
    .X(\t$5006 ));
 sky130_fd_sc_hd__xor2_1 \U$$1177  (.A(\t$5006 ),
    .B(net1010),
    .X(booth_b16_m37));
 sky130_fd_sc_hd__a22o_1 \U$$1178  (.A1(net961),
    .A2(net645),
    .B1(net955),
    .B2(net918),
    .X(\t$5007 ));
 sky130_fd_sc_hd__xor2_1 \U$$1179  (.A(\t$5007 ),
    .B(net1010),
    .X(booth_b16_m38));
 sky130_fd_sc_hd__a22o_1 \U$$118  (.A1(net1615),
    .A2(net449),
    .B1(net1607),
    .B2(net691),
    .X(\t$4466 ));
 sky130_fd_sc_hd__a22o_1 \U$$1180  (.A1(net955),
    .A2(net645),
    .B1(net944),
    .B2(net918),
    .X(\t$5008 ));
 sky130_fd_sc_hd__xor2_1 \U$$1181  (.A(\t$5008 ),
    .B(net1010),
    .X(booth_b16_m39));
 sky130_fd_sc_hd__a22o_1 \U$$1182  (.A1(net944),
    .A2(net645),
    .B1(net928),
    .B2(net918),
    .X(\t$5009 ));
 sky130_fd_sc_hd__xor2_1 \U$$1183  (.A(\t$5009 ),
    .B(net1011),
    .X(booth_b16_m40));
 sky130_fd_sc_hd__a22o_1 \U$$1184  (.A1(net928),
    .A2(net645),
    .B1(net1749),
    .B2(net918),
    .X(\t$5010 ));
 sky130_fd_sc_hd__xor2_1 \U$$1185  (.A(\t$5010 ),
    .B(net1011),
    .X(booth_b16_m41));
 sky130_fd_sc_hd__a22o_1 \U$$1186  (.A1(net1749),
    .A2(net645),
    .B1(net1741),
    .B2(net918),
    .X(\t$5011 ));
 sky130_fd_sc_hd__xor2_1 \U$$1187  (.A(\t$5011 ),
    .B(net1011),
    .X(booth_b16_m42));
 sky130_fd_sc_hd__a22o_1 \U$$1188  (.A1(net1738),
    .A2(net648),
    .B1(net1730),
    .B2(net921),
    .X(\t$5012 ));
 sky130_fd_sc_hd__xor2_1 \U$$1189  (.A(\t$5012 ),
    .B(net1008),
    .X(booth_b16_m43));
 sky130_fd_sc_hd__xor2_1 \U$$119  (.A(\t$4466 ),
    .B(net1576),
    .X(booth_b0_m56));
 sky130_fd_sc_hd__a22o_1 \U$$1190  (.A1(net1730),
    .A2(net648),
    .B1(net1721),
    .B2(net921),
    .X(\t$5013 ));
 sky130_fd_sc_hd__xor2_1 \U$$1191  (.A(\t$5013 ),
    .B(net1008),
    .X(booth_b16_m44));
 sky130_fd_sc_hd__a22o_1 \U$$1192  (.A1(net1720),
    .A2(net648),
    .B1(net1711),
    .B2(net921),
    .X(\t$5014 ));
 sky130_fd_sc_hd__xor2_1 \U$$1193  (.A(\t$5014 ),
    .B(net1007),
    .X(booth_b16_m45));
 sky130_fd_sc_hd__a22o_1 \U$$1194  (.A1(net1711),
    .A2(net648),
    .B1(net1703),
    .B2(net921),
    .X(\t$5015 ));
 sky130_fd_sc_hd__xor2_1 \U$$1195  (.A(\t$5015 ),
    .B(net1007),
    .X(booth_b16_m46));
 sky130_fd_sc_hd__a22o_1 \U$$1196  (.A1(net1703),
    .A2(net648),
    .B1(net1695),
    .B2(net921),
    .X(\t$5016 ));
 sky130_fd_sc_hd__xor2_1 \U$$1197  (.A(\t$5016 ),
    .B(net1008),
    .X(booth_b16_m47));
 sky130_fd_sc_hd__a22o_1 \U$$1198  (.A1(net1698),
    .A2(net650),
    .B1(net1690),
    .B2(net923),
    .X(\t$5017 ));
 sky130_fd_sc_hd__xor2_1 \U$$1199  (.A(\t$5017 ),
    .B(net1014),
    .X(booth_b16_m48));
 sky130_fd_sc_hd__a22o_1 \U$$12  (.A1(net1035),
    .A2(net446),
    .B1(net937),
    .B2(net688),
    .X(\t$4413 ));
 sky130_fd_sc_hd__a22o_1 \U$$120  (.A1(net1607),
    .A2(net450),
    .B1(net1599),
    .B2(net692),
    .X(\t$4467 ));
 sky130_fd_sc_hd__a22o_1 \U$$1200  (.A1(net1690),
    .A2(net650),
    .B1(net1682),
    .B2(net923),
    .X(\t$5018 ));
 sky130_fd_sc_hd__xor2_1 \U$$1201  (.A(\t$5018 ),
    .B(net1014),
    .X(booth_b16_m49));
 sky130_fd_sc_hd__a22o_1 \U$$1202  (.A1(net1682),
    .A2(net650),
    .B1(net1657),
    .B2(net923),
    .X(\t$5019 ));
 sky130_fd_sc_hd__xor2_1 \U$$1203  (.A(\t$5019 ),
    .B(net1011),
    .X(booth_b16_m50));
 sky130_fd_sc_hd__a22o_1 \U$$1204  (.A1(net1657),
    .A2(net650),
    .B1(net1649),
    .B2(net923),
    .X(\t$5020 ));
 sky130_fd_sc_hd__xor2_1 \U$$1205  (.A(\t$5020 ),
    .B(net1014),
    .X(booth_b16_m51));
 sky130_fd_sc_hd__a22o_1 \U$$1206  (.A1(net1649),
    .A2(net650),
    .B1(net1641),
    .B2(net923),
    .X(\t$5021 ));
 sky130_fd_sc_hd__xor2_1 \U$$1207  (.A(\t$5021 ),
    .B(net1014),
    .X(booth_b16_m52));
 sky130_fd_sc_hd__a22o_1 \U$$1208  (.A1(net1641),
    .A2(net650),
    .B1(net1633),
    .B2(net923),
    .X(\t$5022 ));
 sky130_fd_sc_hd__xor2_1 \U$$1209  (.A(\t$5022 ),
    .B(net1014),
    .X(booth_b16_m53));
 sky130_fd_sc_hd__xor2_1 \U$$121  (.A(\t$4467 ),
    .B(net1576),
    .X(booth_b0_m57));
 sky130_fd_sc_hd__a22o_1 \U$$1210  (.A1(net1630),
    .A2(net650),
    .B1(net1621),
    .B2(net923),
    .X(\t$5023 ));
 sky130_fd_sc_hd__xor2_1 \U$$1211  (.A(\t$5023 ),
    .B(net1014),
    .X(booth_b16_m54));
 sky130_fd_sc_hd__a22o_1 \U$$1212  (.A1(net1620),
    .A2(net649),
    .B1(net1612),
    .B2(net922),
    .X(\t$5024 ));
 sky130_fd_sc_hd__xor2_1 \U$$1213  (.A(\t$5024 ),
    .B(net1012),
    .X(booth_b16_m55));
 sky130_fd_sc_hd__a22o_1 \U$$1214  (.A1(net1614),
    .A2(net649),
    .B1(net1606),
    .B2(net922),
    .X(\t$5025 ));
 sky130_fd_sc_hd__xor2_1 \U$$1215  (.A(\t$5025 ),
    .B(net1012),
    .X(booth_b16_m56));
 sky130_fd_sc_hd__a22o_1 \U$$1216  (.A1(net1604),
    .A2(net648),
    .B1(net1595),
    .B2(net921),
    .X(\t$5026 ));
 sky130_fd_sc_hd__xor2_1 \U$$1217  (.A(\t$5026 ),
    .B(net1012),
    .X(booth_b16_m57));
 sky130_fd_sc_hd__a22o_1 \U$$1218  (.A1(net1595),
    .A2(net649),
    .B1(net1586),
    .B2(net922),
    .X(\t$5027 ));
 sky130_fd_sc_hd__xor2_1 \U$$1219  (.A(\t$5027 ),
    .B(net1012),
    .X(booth_b16_m58));
 sky130_fd_sc_hd__a22o_1 \U$$122  (.A1(net1599),
    .A2(net449),
    .B1(net1590),
    .B2(net691),
    .X(\t$4468 ));
 sky130_fd_sc_hd__a22o_1 \U$$1220  (.A1(net1586),
    .A2(net649),
    .B1(net1578),
    .B2(net922),
    .X(\t$5028 ));
 sky130_fd_sc_hd__xor2_1 \U$$1221  (.A(\t$5028 ),
    .B(net1012),
    .X(booth_b16_m59));
 sky130_fd_sc_hd__a22o_1 \U$$1222  (.A1(net1578),
    .A2(net648),
    .B1(net1551),
    .B2(net921),
    .X(\t$5029 ));
 sky130_fd_sc_hd__xor2_1 \U$$1223  (.A(\t$5029 ),
    .B(net1012),
    .X(booth_b16_m60));
 sky130_fd_sc_hd__a22o_1 \U$$1224  (.A1(net1551),
    .A2(net648),
    .B1(net1543),
    .B2(net921),
    .X(\t$5030 ));
 sky130_fd_sc_hd__xor2_1 \U$$1225  (.A(\t$5030 ),
    .B(net1012),
    .X(booth_b16_m61));
 sky130_fd_sc_hd__a22o_1 \U$$1226  (.A1(net1546),
    .A2(net648),
    .B1(net1538),
    .B2(net921),
    .X(\t$5031 ));
 sky130_fd_sc_hd__xor2_1 \U$$1227  (.A(\t$5031 ),
    .B(net1012),
    .X(booth_b16_m62));
 sky130_fd_sc_hd__a22o_1 \U$$1228  (.A1(net1535),
    .A2(net649),
    .B1(net1527),
    .B2(net922),
    .X(\t$5032 ));
 sky130_fd_sc_hd__xor2_1 \U$$1229  (.A(\t$5032 ),
    .B(net1013),
    .X(booth_b16_m63));
 sky130_fd_sc_hd__xor2_1 \U$$123  (.A(\t$4468 ),
    .B(net1576),
    .X(booth_b0_m58));
 sky130_fd_sc_hd__a22o_1 \U$$1230  (.A1(net1527),
    .A2(net649),
    .B1(net1756),
    .B2(net922),
    .X(\t$5033 ));
 sky130_fd_sc_hd__xor2_1 \U$$1231  (.A(\t$5033 ),
    .B(net1013),
    .X(booth_b16_m64));
 sky130_fd_sc_hd__inv_1 \U$$1232  (.A(net1013),
    .Y(\notsign$5034 ));
 sky130_fd_sc_hd__inv_1 \U$$1233  (.A(net1013),
    .Y(\notblock$5035[0] ));
 sky130_fd_sc_hd__inv_1 \U$$1234  (.A(net10),
    .Y(\notblock$5035[1] ));
 sky130_fd_sc_hd__inv_1 \U$$1235  (.A(net1668),
    .Y(\notblock$5035[2] ));
 sky130_fd_sc_hd__and2_1 \U$$1236  (.A(net1668),
    .B(\notblock$5035[1] ),
    .X(\t$5036 ));
 sky130_fd_sc_hd__a32o_2 \U$$1237  (.A1(\notblock$5035[2] ),
    .A2(net10),
    .A3(net1013),
    .B1(\t$5036 ),
    .B2(\notblock$5035[0] ),
    .X(\sel_0$5037 ));
 sky130_fd_sc_hd__xor2_4 \U$$1238  (.A(net10),
    .B(net1013),
    .X(\sel_1$5038 ));
 sky130_fd_sc_hd__a22o_1 \U$$1239  (.A1(net1757),
    .A2(net637),
    .B1(net1228),
    .B2(net910),
    .X(\t$5039 ));
 sky130_fd_sc_hd__a22o_1 \U$$124  (.A1(net1586),
    .A2(net445),
    .B1(net1578),
    .B2(net687),
    .X(\t$4469 ));
 sky130_fd_sc_hd__xor2_1 \U$$1240  (.A(\t$5039 ),
    .B(net1664),
    .X(booth_b18_m0));
 sky130_fd_sc_hd__a22o_1 \U$$1241  (.A1(net1230),
    .A2(net637),
    .B1(net1123),
    .B2(net910),
    .X(\t$5040 ));
 sky130_fd_sc_hd__xor2_1 \U$$1242  (.A(\t$5040 ),
    .B(net1664),
    .X(booth_b18_m1));
 sky130_fd_sc_hd__a22o_1 \U$$1243  (.A1(net1126),
    .A2(net638),
    .B1(net1036),
    .B2(net911),
    .X(\t$5041 ));
 sky130_fd_sc_hd__xor2_1 \U$$1244  (.A(\t$5041 ),
    .B(net1664),
    .X(booth_b18_m2));
 sky130_fd_sc_hd__a22o_1 \U$$1245  (.A1(net1036),
    .A2(net638),
    .B1(net936),
    .B2(net911),
    .X(\t$5042 ));
 sky130_fd_sc_hd__xor2_1 \U$$1246  (.A(\t$5042 ),
    .B(net1665),
    .X(booth_b18_m3));
 sky130_fd_sc_hd__a22o_1 \U$$1247  (.A1(net936),
    .A2(net637),
    .B1(net1676),
    .B2(net910),
    .X(\t$5043 ));
 sky130_fd_sc_hd__xor2_1 \U$$1248  (.A(\t$5043 ),
    .B(net1664),
    .X(booth_b18_m4));
 sky130_fd_sc_hd__a22o_1 \U$$1249  (.A1(net1672),
    .A2(net637),
    .B1(net1561),
    .B2(net910),
    .X(\t$5044 ));
 sky130_fd_sc_hd__xor2_1 \U$$125  (.A(\t$4469 ),
    .B(net1572),
    .X(booth_b0_m59));
 sky130_fd_sc_hd__xor2_1 \U$$1250  (.A(\t$5044 ),
    .B(net1664),
    .X(booth_b18_m5));
 sky130_fd_sc_hd__a22o_1 \U$$1251  (.A1(net1561),
    .A2(net635),
    .B1(net1521),
    .B2(net908),
    .X(\t$5045 ));
 sky130_fd_sc_hd__xor2_1 \U$$1252  (.A(\t$5045 ),
    .B(net1662),
    .X(booth_b18_m6));
 sky130_fd_sc_hd__a22o_1 \U$$1253  (.A1(net1519),
    .A2(net636),
    .B1(net1513),
    .B2(net909),
    .X(\t$5046 ));
 sky130_fd_sc_hd__xor2_1 \U$$1254  (.A(\t$5046 ),
    .B(net1662),
    .X(booth_b18_m7));
 sky130_fd_sc_hd__a22o_1 \U$$1255  (.A1(net1511),
    .A2(net635),
    .B1(net1503),
    .B2(net908),
    .X(\t$5047 ));
 sky130_fd_sc_hd__xor2_1 \U$$1256  (.A(\t$5047 ),
    .B(net1662),
    .X(booth_b18_m8));
 sky130_fd_sc_hd__a22o_1 \U$$1257  (.A1(net1503),
    .A2(net635),
    .B1(net1494),
    .B2(net908),
    .X(\t$5048 ));
 sky130_fd_sc_hd__xor2_1 \U$$1258  (.A(\t$5048 ),
    .B(net1662),
    .X(booth_b18_m9));
 sky130_fd_sc_hd__a22o_1 \U$$1259  (.A1(net1494),
    .A2(net635),
    .B1(net1219),
    .B2(net908),
    .X(\t$5049 ));
 sky130_fd_sc_hd__a22o_1 \U$$126  (.A1(net1581),
    .A2(net445),
    .B1(net1552),
    .B2(net687),
    .X(\t$4470 ));
 sky130_fd_sc_hd__xor2_1 \U$$1260  (.A(\t$5049 ),
    .B(net1662),
    .X(booth_b18_m10));
 sky130_fd_sc_hd__a22o_1 \U$$1261  (.A1(net1219),
    .A2(net635),
    .B1(net1210),
    .B2(net908),
    .X(\t$5050 ));
 sky130_fd_sc_hd__xor2_1 \U$$1262  (.A(\t$5050 ),
    .B(net1662),
    .X(booth_b18_m11));
 sky130_fd_sc_hd__a22o_1 \U$$1263  (.A1(net1210),
    .A2(net635),
    .B1(net1201),
    .B2(net908),
    .X(\t$5051 ));
 sky130_fd_sc_hd__xor2_1 \U$$1264  (.A(\t$5051 ),
    .B(net1662),
    .X(booth_b18_m12));
 sky130_fd_sc_hd__a22o_1 \U$$1265  (.A1(net1201),
    .A2(net635),
    .B1(net1192),
    .B2(net908),
    .X(\t$5052 ));
 sky130_fd_sc_hd__xor2_1 \U$$1266  (.A(\t$5052 ),
    .B(net1662),
    .X(booth_b18_m13));
 sky130_fd_sc_hd__a22o_1 \U$$1267  (.A1(net1195),
    .A2(net637),
    .B1(net1175),
    .B2(net910),
    .X(\t$5053 ));
 sky130_fd_sc_hd__xor2_1 \U$$1268  (.A(\t$5053 ),
    .B(net1664),
    .X(booth_b18_m14));
 sky130_fd_sc_hd__a22o_1 \U$$1269  (.A1(net1179),
    .A2(net638),
    .B1(net1170),
    .B2(net911),
    .X(\t$5054 ));
 sky130_fd_sc_hd__xor2_1 \U$$127  (.A(\t$4470 ),
    .B(net1572),
    .X(booth_b0_m60));
 sky130_fd_sc_hd__xor2_1 \U$$1270  (.A(\t$5054 ),
    .B(net1665),
    .X(booth_b18_m15));
 sky130_fd_sc_hd__a22o_1 \U$$1271  (.A1(net1170),
    .A2(net638),
    .B1(net1161),
    .B2(net911),
    .X(\t$5055 ));
 sky130_fd_sc_hd__xor2_1 \U$$1272  (.A(\t$5055 ),
    .B(net1665),
    .X(booth_b18_m16));
 sky130_fd_sc_hd__a22o_1 \U$$1273  (.A1(net1161),
    .A2(net637),
    .B1(net1149),
    .B2(net910),
    .X(\t$5056 ));
 sky130_fd_sc_hd__xor2_1 \U$$1274  (.A(\t$5056 ),
    .B(net1665),
    .X(booth_b18_m17));
 sky130_fd_sc_hd__a22o_1 \U$$1275  (.A1(net1150),
    .A2(net637),
    .B1(net1143),
    .B2(net910),
    .X(\t$5057 ));
 sky130_fd_sc_hd__xor2_1 \U$$1276  (.A(\t$5057 ),
    .B(net1664),
    .X(booth_b18_m18));
 sky130_fd_sc_hd__a22o_1 \U$$1277  (.A1(net1139),
    .A2(net637),
    .B1(net1130),
    .B2(net910),
    .X(\t$5058 ));
 sky130_fd_sc_hd__xor2_1 \U$$1278  (.A(\t$5058 ),
    .B(net1664),
    .X(booth_b18_m19));
 sky130_fd_sc_hd__a22o_1 \U$$1279  (.A1(net1131),
    .A2(net637),
    .B1(net1115),
    .B2(net910),
    .X(\t$5059 ));
 sky130_fd_sc_hd__a22o_1 \U$$128  (.A1(net1551),
    .A2(net444),
    .B1(net1543),
    .B2(net686),
    .X(\t$4471 ));
 sky130_fd_sc_hd__xor2_1 \U$$1280  (.A(\t$5059 ),
    .B(net1664),
    .X(booth_b18_m20));
 sky130_fd_sc_hd__a22o_1 \U$$1281  (.A1(net1115),
    .A2(net635),
    .B1(net1106),
    .B2(net908),
    .X(\t$5060 ));
 sky130_fd_sc_hd__xor2_1 \U$$1282  (.A(\t$5060 ),
    .B(net1662),
    .X(booth_b18_m21));
 sky130_fd_sc_hd__a22o_1 \U$$1283  (.A1(net1105),
    .A2(net635),
    .B1(net1097),
    .B2(net908),
    .X(\t$5061 ));
 sky130_fd_sc_hd__xor2_1 \U$$1284  (.A(\t$5061 ),
    .B(net1667),
    .X(booth_b18_m22));
 sky130_fd_sc_hd__a22o_1 \U$$1285  (.A1(net1097),
    .A2(net635),
    .B1(net1088),
    .B2(net908),
    .X(\t$5062 ));
 sky130_fd_sc_hd__xor2_1 \U$$1286  (.A(\t$5062 ),
    .B(net1662),
    .X(booth_b18_m23));
 sky130_fd_sc_hd__a22o_1 \U$$1287  (.A1(net1090),
    .A2(net636),
    .B1(net1080),
    .B2(net909),
    .X(\t$5063 ));
 sky130_fd_sc_hd__xor2_1 \U$$1288  (.A(\t$5063 ),
    .B(net1663),
    .X(booth_b18_m24));
 sky130_fd_sc_hd__a22o_1 \U$$1289  (.A1(net1081),
    .A2(net636),
    .B1(net1072),
    .B2(net909),
    .X(\t$5064 ));
 sky130_fd_sc_hd__xor2_1 \U$$129  (.A(\t$4471 ),
    .B(net1570),
    .X(booth_b0_m61));
 sky130_fd_sc_hd__xor2_1 \U$$1290  (.A(\t$5064 ),
    .B(net1663),
    .X(booth_b18_m25));
 sky130_fd_sc_hd__a22o_1 \U$$1291  (.A1(net1073),
    .A2(net636),
    .B1(net1063),
    .B2(net909),
    .X(\t$5065 ));
 sky130_fd_sc_hd__xor2_1 \U$$1292  (.A(\t$5065 ),
    .B(net1663),
    .X(booth_b18_m26));
 sky130_fd_sc_hd__a22o_1 \U$$1293  (.A1(net1064),
    .A2(net639),
    .B1(net1055),
    .B2(net912),
    .X(\t$5066 ));
 sky130_fd_sc_hd__xor2_1 \U$$1294  (.A(\t$5066 ),
    .B(net1663),
    .X(booth_b18_m27));
 sky130_fd_sc_hd__a22o_1 \U$$1295  (.A1(net1056),
    .A2(net639),
    .B1(net1048),
    .B2(net912),
    .X(\t$5067 ));
 sky130_fd_sc_hd__xor2_1 \U$$1296  (.A(\t$5067 ),
    .B(net1663),
    .X(booth_b18_m28));
 sky130_fd_sc_hd__a22o_1 \U$$1297  (.A1(net1048),
    .A2(net636),
    .B1(net1040),
    .B2(net909),
    .X(\t$5068 ));
 sky130_fd_sc_hd__xor2_1 \U$$1298  (.A(\t$5068 ),
    .B(net1663),
    .X(booth_b18_m29));
 sky130_fd_sc_hd__a22o_1 \U$$1299  (.A1(net1040),
    .A2(net636),
    .B1(net1023),
    .B2(net909),
    .X(\t$5069 ));
 sky130_fd_sc_hd__xor2_1 \U$$13  (.A(\t$4413 ),
    .B(net1573),
    .X(booth_b0_m3));
 sky130_fd_sc_hd__a22o_1 \U$$130  (.A1(net1543),
    .A2(net444),
    .B1(net1535),
    .B2(net686),
    .X(\t$4472 ));
 sky130_fd_sc_hd__xor2_1 \U$$1300  (.A(\t$5069 ),
    .B(net1663),
    .X(booth_b18_m30));
 sky130_fd_sc_hd__a22o_1 \U$$1301  (.A1(net1024),
    .A2(net636),
    .B1(net1015),
    .B2(net909),
    .X(\t$5070 ));
 sky130_fd_sc_hd__xor2_1 \U$$1302  (.A(\t$5070 ),
    .B(net1663),
    .X(booth_b18_m31));
 sky130_fd_sc_hd__a22o_1 \U$$1303  (.A1(net1015),
    .A2(net639),
    .B1(net998),
    .B2(net912),
    .X(\t$5071 ));
 sky130_fd_sc_hd__xor2_1 \U$$1304  (.A(\t$5071 ),
    .B(net1666),
    .X(booth_b18_m32));
 sky130_fd_sc_hd__a22o_1 \U$$1305  (.A1(net1000),
    .A2(net638),
    .B1(net992),
    .B2(net911),
    .X(\t$5072 ));
 sky130_fd_sc_hd__xor2_1 \U$$1306  (.A(\t$5072 ),
    .B(net1666),
    .X(booth_b18_m33));
 sky130_fd_sc_hd__a22o_1 \U$$1307  (.A1(net992),
    .A2(net637),
    .B1(net987),
    .B2(net910),
    .X(\t$5073 ));
 sky130_fd_sc_hd__xor2_1 \U$$1308  (.A(\t$5073 ),
    .B(net1665),
    .X(booth_b18_m34));
 sky130_fd_sc_hd__a22o_1 \U$$1309  (.A1(net987),
    .A2(net639),
    .B1(net978),
    .B2(net912),
    .X(\t$5074 ));
 sky130_fd_sc_hd__xor2_1 \U$$131  (.A(\t$4472 ),
    .B(net1570),
    .X(booth_b0_m62));
 sky130_fd_sc_hd__xor2_1 \U$$1310  (.A(\t$5074 ),
    .B(net1666),
    .X(booth_b18_m35));
 sky130_fd_sc_hd__a22o_1 \U$$1311  (.A1(net978),
    .A2(net638),
    .B1(net972),
    .B2(net911),
    .X(\t$5075 ));
 sky130_fd_sc_hd__xor2_1 \U$$1312  (.A(\t$5075 ),
    .B(net1666),
    .X(booth_b18_m36));
 sky130_fd_sc_hd__a22o_1 \U$$1313  (.A1(net969),
    .A2(net638),
    .B1(net961),
    .B2(net911),
    .X(\t$5076 ));
 sky130_fd_sc_hd__xor2_1 \U$$1314  (.A(\t$5076 ),
    .B(net1666),
    .X(booth_b18_m37));
 sky130_fd_sc_hd__a22o_1 \U$$1315  (.A1(net957),
    .A2(net638),
    .B1(net949),
    .B2(net911),
    .X(\t$5077 ));
 sky130_fd_sc_hd__xor2_1 \U$$1316  (.A(\t$5077 ),
    .B(net1666),
    .X(booth_b18_m38));
 sky130_fd_sc_hd__a22o_1 \U$$1317  (.A1(net955),
    .A2(net638),
    .B1(net944),
    .B2(net911),
    .X(\t$5078 ));
 sky130_fd_sc_hd__xor2_1 \U$$1318  (.A(\t$5078 ),
    .B(net1666),
    .X(booth_b18_m39));
 sky130_fd_sc_hd__a22o_1 \U$$1319  (.A1(net944),
    .A2(net639),
    .B1(net928),
    .B2(net912),
    .X(\t$5079 ));
 sky130_fd_sc_hd__a22o_1 \U$$132  (.A1(net1535),
    .A2(net444),
    .B1(net1527),
    .B2(net686),
    .X(\t$4473 ));
 sky130_fd_sc_hd__xor2_1 \U$$1320  (.A(\t$5079 ),
    .B(net1666),
    .X(booth_b18_m40));
 sky130_fd_sc_hd__a22o_1 \U$$1321  (.A1(net925),
    .A2(net640),
    .B1(net1746),
    .B2(net913),
    .X(\t$5080 ));
 sky130_fd_sc_hd__xor2_1 \U$$1322  (.A(\t$5080 ),
    .B(net1669),
    .X(booth_b18_m41));
 sky130_fd_sc_hd__a22o_1 \U$$1323  (.A1(net1746),
    .A2(net640),
    .B1(net1738),
    .B2(net913),
    .X(\t$5081 ));
 sky130_fd_sc_hd__xor2_1 \U$$1324  (.A(\t$5081 ),
    .B(net1667),
    .X(booth_b18_m42));
 sky130_fd_sc_hd__a22o_1 \U$$1325  (.A1(net1737),
    .A2(net636),
    .B1(net1729),
    .B2(net909),
    .X(\t$5082 ));
 sky130_fd_sc_hd__xor2_1 \U$$1326  (.A(\t$5082 ),
    .B(net1663),
    .X(booth_b18_m43));
 sky130_fd_sc_hd__a22o_1 \U$$1327  (.A1(net1729),
    .A2(net636),
    .B1(net1720),
    .B2(net909),
    .X(\t$5083 ));
 sky130_fd_sc_hd__xor2_1 \U$$1328  (.A(\t$5083 ),
    .B(net1663),
    .X(booth_b18_m44));
 sky130_fd_sc_hd__a22o_1 \U$$1329  (.A1(net1721),
    .A2(net640),
    .B1(net1712),
    .B2(net913),
    .X(\t$5084 ));
 sky130_fd_sc_hd__xor2_1 \U$$133  (.A(\t$4473 ),
    .B(net1570),
    .X(booth_b0_m63));
 sky130_fd_sc_hd__xor2_1 \U$$1330  (.A(\t$5084 ),
    .B(net1669),
    .X(booth_b18_m45));
 sky130_fd_sc_hd__a22o_1 \U$$1331  (.A1(net1715),
    .A2(net642),
    .B1(net1706),
    .B2(net915),
    .X(\t$5085 ));
 sky130_fd_sc_hd__xor2_1 \U$$1332  (.A(\t$5085 ),
    .B(net1670),
    .X(booth_b18_m46));
 sky130_fd_sc_hd__a22o_1 \U$$1333  (.A1(net1706),
    .A2(net642),
    .B1(net1698),
    .B2(net915),
    .X(\t$5086 ));
 sky130_fd_sc_hd__xor2_1 \U$$1334  (.A(\t$5086 ),
    .B(net1670),
    .X(booth_b18_m47));
 sky130_fd_sc_hd__a22o_1 \U$$1335  (.A1(net1698),
    .A2(net642),
    .B1(net1690),
    .B2(net915),
    .X(\t$5087 ));
 sky130_fd_sc_hd__xor2_1 \U$$1336  (.A(\t$5087 ),
    .B(net1667),
    .X(booth_b18_m48));
 sky130_fd_sc_hd__a22o_1 \U$$1337  (.A1(net1692),
    .A2(net642),
    .B1(net1680),
    .B2(net915),
    .X(\t$5088 ));
 sky130_fd_sc_hd__xor2_1 \U$$1338  (.A(\t$5088 ),
    .B(net1670),
    .X(booth_b18_m49));
 sky130_fd_sc_hd__a22o_1 \U$$1339  (.A1(net1682),
    .A2(net642),
    .B1(net1657),
    .B2(net915),
    .X(\t$5089 ));
 sky130_fd_sc_hd__a22o_1 \U$$134  (.A1(net1527),
    .A2(net444),
    .B1(net1758),
    .B2(net686),
    .X(\t$4474 ));
 sky130_fd_sc_hd__xor2_1 \U$$1340  (.A(\t$5089 ),
    .B(net1670),
    .X(booth_b18_m50));
 sky130_fd_sc_hd__a22o_1 \U$$1341  (.A1(net1657),
    .A2(net642),
    .B1(net1649),
    .B2(net915),
    .X(\t$5090 ));
 sky130_fd_sc_hd__xor2_1 \U$$1342  (.A(\t$5090 ),
    .B(net1670),
    .X(booth_b18_m51));
 sky130_fd_sc_hd__a22o_1 \U$$1343  (.A1(net1646),
    .A2(net642),
    .B1(net1640),
    .B2(net915),
    .X(\t$5091 ));
 sky130_fd_sc_hd__xor2_1 \U$$1344  (.A(\t$5091 ),
    .B(net1670),
    .X(booth_b18_m52));
 sky130_fd_sc_hd__a22o_1 \U$$1345  (.A1(net1638),
    .A2(net640),
    .B1(net1629),
    .B2(net913),
    .X(\t$5092 ));
 sky130_fd_sc_hd__xor2_1 \U$$1346  (.A(\t$5092 ),
    .B(net1669),
    .X(booth_b18_m53));
 sky130_fd_sc_hd__a22o_1 \U$$1347  (.A1(net1629),
    .A2(net640),
    .B1(net1620),
    .B2(net913),
    .X(\t$5093 ));
 sky130_fd_sc_hd__xor2_1 \U$$1348  (.A(\t$5093 ),
    .B(net1669),
    .X(booth_b18_m54));
 sky130_fd_sc_hd__a22o_1 \U$$1349  (.A1(net1620),
    .A2(net640),
    .B1(net1612),
    .B2(net913),
    .X(\t$5094 ));
 sky130_fd_sc_hd__xor2_1 \U$$135  (.A(\t$4474 ),
    .B(net1571),
    .X(booth_b0_m64));
 sky130_fd_sc_hd__xor2_1 \U$$1350  (.A(\t$5094 ),
    .B(net1669),
    .X(booth_b18_m55));
 sky130_fd_sc_hd__a22o_1 \U$$1351  (.A1(net1612),
    .A2(net640),
    .B1(net1604),
    .B2(net913),
    .X(\t$5095 ));
 sky130_fd_sc_hd__xor2_1 \U$$1352  (.A(\t$5095 ),
    .B(net1669),
    .X(booth_b18_m56));
 sky130_fd_sc_hd__a22o_1 \U$$1353  (.A1(net1604),
    .A2(net640),
    .B1(net1595),
    .B2(net913),
    .X(\t$5096 ));
 sky130_fd_sc_hd__xor2_1 \U$$1354  (.A(\t$5096 ),
    .B(net1669),
    .X(booth_b18_m57));
 sky130_fd_sc_hd__a22o_1 \U$$1355  (.A1(net1595),
    .A2(net640),
    .B1(net1586),
    .B2(net913),
    .X(\t$5097 ));
 sky130_fd_sc_hd__xor2_1 \U$$1356  (.A(\t$5097 ),
    .B(net1669),
    .X(booth_b18_m58));
 sky130_fd_sc_hd__a22o_1 \U$$1357  (.A1(net1587),
    .A2(net640),
    .B1(net1581),
    .B2(net913),
    .X(\t$5098 ));
 sky130_fd_sc_hd__xor2_1 \U$$1358  (.A(\t$5098 ),
    .B(net1668),
    .X(booth_b18_m59));
 sky130_fd_sc_hd__a22o_1 \U$$1359  (.A1(net1581),
    .A2(net641),
    .B1(net1552),
    .B2(net914),
    .X(\t$5099 ));
 sky130_fd_sc_hd__inv_1 \U$$136  (.A(net1577),
    .Y(notsign));
 sky130_fd_sc_hd__xor2_1 \U$$1360  (.A(\t$5099 ),
    .B(net1668),
    .X(booth_b18_m60));
 sky130_fd_sc_hd__a22o_1 \U$$1361  (.A1(net1552),
    .A2(net641),
    .B1(net1546),
    .B2(net914),
    .X(\t$5100 ));
 sky130_fd_sc_hd__xor2_1 \U$$1362  (.A(\t$5100 ),
    .B(net1668),
    .X(booth_b18_m61));
 sky130_fd_sc_hd__a22o_1 \U$$1363  (.A1(net1544),
    .A2(net641),
    .B1(net1536),
    .B2(net914),
    .X(\t$5101 ));
 sky130_fd_sc_hd__xor2_1 \U$$1364  (.A(\t$5101 ),
    .B(net1670),
    .X(booth_b18_m62));
 sky130_fd_sc_hd__a22o_1 \U$$1365  (.A1(net1537),
    .A2(net641),
    .B1(net1528),
    .B2(net914),
    .X(\t$5102 ));
 sky130_fd_sc_hd__xor2_1 \U$$1366  (.A(\t$5102 ),
    .B(net1669),
    .X(booth_b18_m63));
 sky130_fd_sc_hd__a22o_1 \U$$1367  (.A1(net1528),
    .A2(net641),
    .B1(net1759),
    .B2(net914),
    .X(\t$5103 ));
 sky130_fd_sc_hd__xor2_1 \U$$1368  (.A(\t$5103 ),
    .B(net1668),
    .X(booth_b18_m64));
 sky130_fd_sc_hd__inv_1 \U$$1369  (.A(net1668),
    .Y(\notsign$5104 ));
 sky130_fd_sc_hd__inv_1 \U$$137  (.A(net1571),
    .Y(\notblock$4475[0] ));
 sky130_fd_sc_hd__inv_1 \U$$1370  (.A(net1668),
    .Y(\notblock$5105[0] ));
 sky130_fd_sc_hd__inv_1 \U$$1371  (.A(net13),
    .Y(\notblock$5105[1] ));
 sky130_fd_sc_hd__inv_1 \U$$1372  (.A(net1491),
    .Y(\notblock$5105[2] ));
 sky130_fd_sc_hd__and2_1 \U$$1373  (.A(net1491),
    .B(\notblock$5105[1] ),
    .X(\t$5106 ));
 sky130_fd_sc_hd__a32o_2 \U$$1374  (.A1(\notblock$5105[2] ),
    .A2(net13),
    .A3(net1668),
    .B1(\t$5106 ),
    .B2(\notblock$5105[0] ),
    .X(\sel_0$5107 ));
 sky130_fd_sc_hd__xor2_4 \U$$1375  (.A(net13),
    .B(net1668),
    .X(\sel_1$5108 ));
 sky130_fd_sc_hd__a22o_1 \U$$1376  (.A1(net1760),
    .A2(net630),
    .B1(net1230),
    .B2(net903),
    .X(\t$5109 ));
 sky130_fd_sc_hd__xor2_1 \U$$1377  (.A(\t$5109 ),
    .B(net1487),
    .X(booth_b20_m0));
 sky130_fd_sc_hd__a22o_1 \U$$1378  (.A1(net1230),
    .A2(net630),
    .B1(net1126),
    .B2(net903),
    .X(\t$5110 ));
 sky130_fd_sc_hd__xor2_1 \U$$1379  (.A(\t$5110 ),
    .B(net1487),
    .X(booth_b20_m1));
 sky130_fd_sc_hd__inv_1 \U$$138  (.A(net23),
    .Y(\notblock$4475[1] ));
 sky130_fd_sc_hd__a22o_1 \U$$1380  (.A1(net1126),
    .A2(net629),
    .B1(net1036),
    .B2(net902),
    .X(\t$5111 ));
 sky130_fd_sc_hd__xor2_1 \U$$1381  (.A(\t$5111 ),
    .B(net1487),
    .X(booth_b20_m2));
 sky130_fd_sc_hd__a22o_1 \U$$1382  (.A1(net1036),
    .A2(net629),
    .B1(net933),
    .B2(net902),
    .X(\t$5112 ));
 sky130_fd_sc_hd__xor2_1 \U$$1383  (.A(\t$5112 ),
    .B(net1487),
    .X(booth_b20_m3));
 sky130_fd_sc_hd__a22o_1 \U$$1384  (.A1(net933),
    .A2(net627),
    .B1(net1672),
    .B2(net900),
    .X(\t$5113 ));
 sky130_fd_sc_hd__xor2_1 \U$$1385  (.A(\t$5113 ),
    .B(net1485),
    .X(booth_b20_m4));
 sky130_fd_sc_hd__a22o_1 \U$$1386  (.A1(net1671),
    .A2(net628),
    .B1(net1560),
    .B2(net901),
    .X(\t$5114 ));
 sky130_fd_sc_hd__xor2_1 \U$$1387  (.A(\t$5114 ),
    .B(net1485),
    .X(booth_b20_m5));
 sky130_fd_sc_hd__a22o_1 \U$$1388  (.A1(net1560),
    .A2(net627),
    .B1(net1519),
    .B2(net900),
    .X(\t$5115 ));
 sky130_fd_sc_hd__xor2_1 \U$$1389  (.A(\t$5115 ),
    .B(net1485),
    .X(booth_b20_m6));
 sky130_fd_sc_hd__inv_1 \U$$139  (.A(net1387),
    .Y(\notblock$4475[2] ));
 sky130_fd_sc_hd__a22o_1 \U$$1390  (.A1(net1519),
    .A2(net627),
    .B1(net1511),
    .B2(net900),
    .X(\t$5116 ));
 sky130_fd_sc_hd__xor2_1 \U$$1391  (.A(\t$5116 ),
    .B(net1485),
    .X(booth_b20_m7));
 sky130_fd_sc_hd__a22o_1 \U$$1392  (.A1(net1511),
    .A2(net627),
    .B1(net1503),
    .B2(net900),
    .X(\t$5117 ));
 sky130_fd_sc_hd__xor2_1 \U$$1393  (.A(\t$5117 ),
    .B(net1485),
    .X(booth_b20_m8));
 sky130_fd_sc_hd__a22o_1 \U$$1394  (.A1(net1503),
    .A2(net627),
    .B1(net1494),
    .B2(net900),
    .X(\t$5118 ));
 sky130_fd_sc_hd__xor2_1 \U$$1395  (.A(\t$5118 ),
    .B(net1485),
    .X(booth_b20_m9));
 sky130_fd_sc_hd__a22o_1 \U$$1396  (.A1(net1494),
    .A2(net627),
    .B1(net1219),
    .B2(net900),
    .X(\t$5119 ));
 sky130_fd_sc_hd__xor2_1 \U$$1397  (.A(\t$5119 ),
    .B(net1485),
    .X(booth_b20_m10));
 sky130_fd_sc_hd__a22o_1 \U$$1398  (.A1(net1219),
    .A2(net627),
    .B1(net1210),
    .B2(net900),
    .X(\t$5120 ));
 sky130_fd_sc_hd__xor2_1 \U$$1399  (.A(\t$5120 ),
    .B(net1485),
    .X(booth_b20_m11));
 sky130_fd_sc_hd__a22o_1 \U$$14  (.A1(net937),
    .A2(net447),
    .B1(net1675),
    .B2(net689),
    .X(\t$4414 ));
 sky130_fd_sc_hd__and2_1 \U$$140  (.A(net1387),
    .B(\notblock$4475[1] ),
    .X(\t$4476 ));
 sky130_fd_sc_hd__a22o_1 \U$$1400  (.A1(net1212),
    .A2(net629),
    .B1(net1203),
    .B2(net902),
    .X(\t$5121 ));
 sky130_fd_sc_hd__xor2_1 \U$$1401  (.A(\t$5121 ),
    .B(net1487),
    .X(booth_b20_m12));
 sky130_fd_sc_hd__a22o_1 \U$$1402  (.A1(net1206),
    .A2(net629),
    .B1(net1198),
    .B2(net902),
    .X(\t$5122 ));
 sky130_fd_sc_hd__xor2_1 \U$$1403  (.A(\t$5122 ),
    .B(net1488),
    .X(booth_b20_m13));
 sky130_fd_sc_hd__a22o_1 \U$$1404  (.A1(net1198),
    .A2(net629),
    .B1(net1179),
    .B2(net902),
    .X(\t$5123 ));
 sky130_fd_sc_hd__xor2_1 \U$$1405  (.A(\t$5123 ),
    .B(net1488),
    .X(booth_b20_m14));
 sky130_fd_sc_hd__a22o_1 \U$$1406  (.A1(net1179),
    .A2(net629),
    .B1(net1170),
    .B2(net902),
    .X(\t$5124 ));
 sky130_fd_sc_hd__xor2_1 \U$$1407  (.A(\t$5124 ),
    .B(net1488),
    .X(booth_b20_m15));
 sky130_fd_sc_hd__a22o_1 \U$$1408  (.A1(net1170),
    .A2(net629),
    .B1(net1161),
    .B2(net902),
    .X(\t$5125 ));
 sky130_fd_sc_hd__xor2_1 \U$$1409  (.A(\t$5125 ),
    .B(net1487),
    .X(booth_b20_m16));
 sky130_fd_sc_hd__a32o_4 \U$$141  (.A1(\notblock$4475[2] ),
    .A2(net23),
    .A3(net1571),
    .B1(\t$4476 ),
    .B2(\notblock$4475[0] ),
    .X(\sel_0$4477 ));
 sky130_fd_sc_hd__a22o_1 \U$$1410  (.A1(net1157),
    .A2(net629),
    .B1(net1147),
    .B2(net902),
    .X(\t$5126 ));
 sky130_fd_sc_hd__xor2_1 \U$$1411  (.A(\t$5126 ),
    .B(net1487),
    .X(booth_b20_m17));
 sky130_fd_sc_hd__a22o_1 \U$$1412  (.A1(net1146),
    .A2(net629),
    .B1(net1139),
    .B2(net902),
    .X(\t$5127 ));
 sky130_fd_sc_hd__xor2_1 \U$$1413  (.A(\t$5127 ),
    .B(net1487),
    .X(booth_b20_m18));
 sky130_fd_sc_hd__a22o_1 \U$$1414  (.A1(net1139),
    .A2(net627),
    .B1(net1131),
    .B2(net900),
    .X(\t$5128 ));
 sky130_fd_sc_hd__xor2_1 \U$$1415  (.A(\t$5128 ),
    .B(net1486),
    .X(booth_b20_m19));
 sky130_fd_sc_hd__a22o_1 \U$$1416  (.A1(net1130),
    .A2(net627),
    .B1(net1114),
    .B2(net900),
    .X(\t$5129 ));
 sky130_fd_sc_hd__xor2_1 \U$$1417  (.A(\t$5129 ),
    .B(net1486),
    .X(booth_b20_m20));
 sky130_fd_sc_hd__a22o_1 \U$$1418  (.A1(net1114),
    .A2(net627),
    .B1(net1105),
    .B2(net900),
    .X(\t$5130 ));
 sky130_fd_sc_hd__xor2_1 \U$$1419  (.A(\t$5130 ),
    .B(net1485),
    .X(booth_b20_m21));
 sky130_fd_sc_hd__xor2_4 \U$$142  (.A(net23),
    .B(net1571),
    .X(\sel_1$4478 ));
 sky130_fd_sc_hd__a22o_1 \U$$1420  (.A1(net1107),
    .A2(net628),
    .B1(net1098),
    .B2(net901),
    .X(\t$5131 ));
 sky130_fd_sc_hd__xor2_1 \U$$1421  (.A(\t$5131 ),
    .B(net1486),
    .X(booth_b20_m22));
 sky130_fd_sc_hd__a22o_1 \U$$1422  (.A1(net1097),
    .A2(net631),
    .B1(net1088),
    .B2(net904),
    .X(\t$5132 ));
 sky130_fd_sc_hd__xor2_1 \U$$1423  (.A(\t$5132 ),
    .B(net1485),
    .X(booth_b20_m23));
 sky130_fd_sc_hd__a22o_1 \U$$1424  (.A1(net1089),
    .A2(net628),
    .B1(net1081),
    .B2(net901),
    .X(\t$5133 ));
 sky130_fd_sc_hd__xor2_1 \U$$1425  (.A(\t$5133 ),
    .B(net1486),
    .X(booth_b20_m24));
 sky130_fd_sc_hd__a22o_1 \U$$1426  (.A1(net1081),
    .A2(net628),
    .B1(net1072),
    .B2(net901),
    .X(\t$5134 ));
 sky130_fd_sc_hd__xor2_1 \U$$1427  (.A(\t$5134 ),
    .B(net1486),
    .X(booth_b20_m25));
 sky130_fd_sc_hd__a22o_1 \U$$1428  (.A1(net1072),
    .A2(net628),
    .B1(net1064),
    .B2(net901),
    .X(\t$5135 ));
 sky130_fd_sc_hd__xor2_1 \U$$1429  (.A(\t$5135 ),
    .B(net1486),
    .X(booth_b20_m26));
 sky130_fd_sc_hd__a22o_1 \U$$143  (.A1(net1761),
    .A2(net624),
    .B1(net1231),
    .B2(net897),
    .X(\t$4479 ));
 sky130_fd_sc_hd__a22o_1 \U$$1430  (.A1(net1064),
    .A2(net628),
    .B1(net1056),
    .B2(net901),
    .X(\t$5136 ));
 sky130_fd_sc_hd__xor2_1 \U$$1431  (.A(\t$5136 ),
    .B(net1486),
    .X(booth_b20_m27));
 sky130_fd_sc_hd__a22o_1 \U$$1432  (.A1(net1056),
    .A2(net628),
    .B1(net1048),
    .B2(net901),
    .X(\t$5137 ));
 sky130_fd_sc_hd__xor2_1 \U$$1433  (.A(\t$5137 ),
    .B(net1486),
    .X(booth_b20_m28));
 sky130_fd_sc_hd__a22o_1 \U$$1434  (.A1(net1048),
    .A2(net628),
    .B1(net1040),
    .B2(net901),
    .X(\t$5138 ));
 sky130_fd_sc_hd__xor2_1 \U$$1435  (.A(\t$5138 ),
    .B(net1486),
    .X(booth_b20_m29));
 sky130_fd_sc_hd__a22o_1 \U$$1436  (.A1(net1041),
    .A2(net631),
    .B1(net1025),
    .B2(net904),
    .X(\t$5139 ));
 sky130_fd_sc_hd__xor2_1 \U$$1437  (.A(\t$5139 ),
    .B(net1487),
    .X(booth_b20_m30));
 sky130_fd_sc_hd__a22o_1 \U$$1438  (.A1(net1025),
    .A2(net630),
    .B1(net1017),
    .B2(net903),
    .X(\t$5140 ));
 sky130_fd_sc_hd__xor2_1 \U$$1439  (.A(\t$5140 ),
    .B(net1489),
    .X(booth_b20_m31));
 sky130_fd_sc_hd__xor2_1 \U$$144  (.A(\t$4479 ),
    .B(net1390),
    .X(booth_b2_m0));
 sky130_fd_sc_hd__a22o_1 \U$$1440  (.A1(net1017),
    .A2(net629),
    .B1(net1000),
    .B2(net902),
    .X(\t$5141 ));
 sky130_fd_sc_hd__xor2_1 \U$$1441  (.A(\t$5141 ),
    .B(net1488),
    .X(booth_b20_m32));
 sky130_fd_sc_hd__a22o_1 \U$$1442  (.A1(net1000),
    .A2(net630),
    .B1(net992),
    .B2(net903),
    .X(\t$5142 ));
 sky130_fd_sc_hd__xor2_1 \U$$1443  (.A(\t$5142 ),
    .B(net1488),
    .X(booth_b20_m33));
 sky130_fd_sc_hd__a22o_1 \U$$1444  (.A1(net993),
    .A2(net630),
    .B1(net987),
    .B2(net903),
    .X(\t$5143 ));
 sky130_fd_sc_hd__xor2_1 \U$$1445  (.A(\t$5143 ),
    .B(net1489),
    .X(booth_b20_m34));
 sky130_fd_sc_hd__a22o_1 \U$$1446  (.A1(net987),
    .A2(net630),
    .B1(net977),
    .B2(net903),
    .X(\t$5144 ));
 sky130_fd_sc_hd__xor2_1 \U$$1447  (.A(\t$5144 ),
    .B(net1489),
    .X(booth_b20_m35));
 sky130_fd_sc_hd__a22o_1 \U$$1448  (.A1(net977),
    .A2(net630),
    .B1(net969),
    .B2(net903),
    .X(\t$5145 ));
 sky130_fd_sc_hd__xor2_1 \U$$1449  (.A(\t$5145 ),
    .B(net1489),
    .X(booth_b20_m36));
 sky130_fd_sc_hd__a22o_1 \U$$145  (.A1(net1231),
    .A2(net624),
    .B1(net1127),
    .B2(net897),
    .X(\t$4480 ));
 sky130_fd_sc_hd__a22o_1 \U$$1450  (.A1(net969),
    .A2(net630),
    .B1(net961),
    .B2(net903),
    .X(\t$5146 ));
 sky130_fd_sc_hd__xor2_1 \U$$1451  (.A(\t$5146 ),
    .B(net1489),
    .X(booth_b20_m37));
 sky130_fd_sc_hd__a22o_1 \U$$1452  (.A1(net961),
    .A2(net631),
    .B1(net955),
    .B2(net904),
    .X(\t$5147 ));
 sky130_fd_sc_hd__xor2_1 \U$$1453  (.A(\t$5147 ),
    .B(net1489),
    .X(booth_b20_m38));
 sky130_fd_sc_hd__a22o_1 \U$$1454  (.A1(net949),
    .A2(net632),
    .B1(net941),
    .B2(net905),
    .X(\t$5148 ));
 sky130_fd_sc_hd__xor2_1 \U$$1455  (.A(\t$5148 ),
    .B(net1490),
    .X(booth_b20_m39));
 sky130_fd_sc_hd__a22o_1 \U$$1456  (.A1(net941),
    .A2(net632),
    .B1(net925),
    .B2(net905),
    .X(\t$5149 ));
 sky130_fd_sc_hd__xor2_1 \U$$1457  (.A(\t$5149 ),
    .B(net1490),
    .X(booth_b20_m40));
 sky130_fd_sc_hd__a22o_1 \U$$1458  (.A1(net925),
    .A2(net628),
    .B1(net1745),
    .B2(net901),
    .X(\t$5150 ));
 sky130_fd_sc_hd__xor2_1 \U$$1459  (.A(\t$5150 ),
    .B(net1490),
    .X(booth_b20_m41));
 sky130_fd_sc_hd__xor2_1 \U$$146  (.A(\t$4480 ),
    .B(net1390),
    .X(booth_b2_m1));
 sky130_fd_sc_hd__a22o_1 \U$$1460  (.A1(net1745),
    .A2(net631),
    .B1(net1737),
    .B2(net904),
    .X(\t$5151 ));
 sky130_fd_sc_hd__xor2_1 \U$$1461  (.A(\t$5151 ),
    .B(net1490),
    .X(booth_b20_m42));
 sky130_fd_sc_hd__a22o_1 \U$$1462  (.A1(net1738),
    .A2(net632),
    .B1(net1730),
    .B2(net905),
    .X(\t$5152 ));
 sky130_fd_sc_hd__xor2_1 \U$$1463  (.A(\t$5152 ),
    .B(net1492),
    .X(booth_b20_m43));
 sky130_fd_sc_hd__a22o_1 \U$$1464  (.A1(net1733),
    .A2(net634),
    .B1(net1724),
    .B2(net907),
    .X(\t$5153 ));
 sky130_fd_sc_hd__xor2_1 \U$$1465  (.A(\t$5153 ),
    .B(net1493),
    .X(booth_b20_m44));
 sky130_fd_sc_hd__a22o_1 \U$$1466  (.A1(net1724),
    .A2(net634),
    .B1(net1715),
    .B2(net907),
    .X(\t$5154 ));
 sky130_fd_sc_hd__xor2_1 \U$$1467  (.A(\t$5154 ),
    .B(net1493),
    .X(booth_b20_m45));
 sky130_fd_sc_hd__a22o_1 \U$$1468  (.A1(net1715),
    .A2(net630),
    .B1(net1706),
    .B2(net903),
    .X(\t$5155 ));
 sky130_fd_sc_hd__xor2_1 \U$$1469  (.A(\t$5155 ),
    .B(net1489),
    .X(booth_b20_m46));
 sky130_fd_sc_hd__a22o_1 \U$$147  (.A1(net1127),
    .A2(net624),
    .B1(net1035),
    .B2(net897),
    .X(\t$4481 ));
 sky130_fd_sc_hd__a22o_1 \U$$1470  (.A1(net1710),
    .A2(net634),
    .B1(net1702),
    .B2(net907),
    .X(\t$5156 ));
 sky130_fd_sc_hd__xor2_1 \U$$1471  (.A(\t$5156 ),
    .B(net1493),
    .X(booth_b20_m47));
 sky130_fd_sc_hd__a22o_1 \U$$1472  (.A1(net1702),
    .A2(net634),
    .B1(net1692),
    .B2(net907),
    .X(\t$5157 ));
 sky130_fd_sc_hd__xor2_1 \U$$1473  (.A(\t$5157 ),
    .B(net1493),
    .X(booth_b20_m48));
 sky130_fd_sc_hd__a22o_1 \U$$1474  (.A1(net1690),
    .A2(net634),
    .B1(net1682),
    .B2(net907),
    .X(\t$5158 ));
 sky130_fd_sc_hd__xor2_1 \U$$1475  (.A(\t$5158 ),
    .B(net1493),
    .X(booth_b20_m49));
 sky130_fd_sc_hd__a22o_1 \U$$1476  (.A1(net1683),
    .A2(net634),
    .B1(net1657),
    .B2(net907),
    .X(\t$5159 ));
 sky130_fd_sc_hd__xor2_1 \U$$1477  (.A(\t$5159 ),
    .B(net1493),
    .X(booth_b20_m50));
 sky130_fd_sc_hd__a22o_1 \U$$1478  (.A1(net1654),
    .A2(net632),
    .B1(net1646),
    .B2(net905),
    .X(\t$5160 ));
 sky130_fd_sc_hd__xor2_1 \U$$1479  (.A(\t$5160 ),
    .B(net1492),
    .X(booth_b20_m51));
 sky130_fd_sc_hd__xor2_1 \U$$148  (.A(\t$4481 ),
    .B(net1390),
    .X(booth_b2_m2));
 sky130_fd_sc_hd__a22o_1 \U$$1480  (.A1(net1646),
    .A2(net632),
    .B1(net1640),
    .B2(net905),
    .X(\t$5161 ));
 sky130_fd_sc_hd__xor2_1 \U$$1481  (.A(\t$5161 ),
    .B(net1492),
    .X(booth_b20_m52));
 sky130_fd_sc_hd__a22o_1 \U$$1482  (.A1(net1638),
    .A2(net632),
    .B1(net1629),
    .B2(net905),
    .X(\t$5162 ));
 sky130_fd_sc_hd__xor2_1 \U$$1483  (.A(\t$5162 ),
    .B(net1492),
    .X(booth_b20_m53));
 sky130_fd_sc_hd__a22o_1 \U$$1484  (.A1(net1629),
    .A2(net632),
    .B1(net1620),
    .B2(net905),
    .X(\t$5163 ));
 sky130_fd_sc_hd__xor2_1 \U$$1485  (.A(\t$5163 ),
    .B(net1492),
    .X(booth_b20_m54));
 sky130_fd_sc_hd__a22o_1 \U$$1486  (.A1(net1620),
    .A2(net632),
    .B1(net1612),
    .B2(net905),
    .X(\t$5164 ));
 sky130_fd_sc_hd__xor2_1 \U$$1487  (.A(\t$5164 ),
    .B(net1492),
    .X(booth_b20_m55));
 sky130_fd_sc_hd__a22o_1 \U$$1488  (.A1(net1612),
    .A2(net633),
    .B1(net1604),
    .B2(net906),
    .X(\t$5165 ));
 sky130_fd_sc_hd__xor2_1 \U$$1489  (.A(\t$5165 ),
    .B(net1492),
    .X(booth_b20_m56));
 sky130_fd_sc_hd__a22o_1 \U$$149  (.A1(net1035),
    .A2(net624),
    .B1(net937),
    .B2(net897),
    .X(\t$4482 ));
 sky130_fd_sc_hd__a22o_1 \U$$1490  (.A1(net1606),
    .A2(net632),
    .B1(net1596),
    .B2(net905),
    .X(\t$5166 ));
 sky130_fd_sc_hd__xor2_1 \U$$1491  (.A(\t$5166 ),
    .B(net1492),
    .X(booth_b20_m57));
 sky130_fd_sc_hd__a22o_1 \U$$1492  (.A1(net1596),
    .A2(net632),
    .B1(net1587),
    .B2(net905),
    .X(\t$5167 ));
 sky130_fd_sc_hd__xor2_1 \U$$1493  (.A(\t$5167 ),
    .B(net1492),
    .X(booth_b20_m58));
 sky130_fd_sc_hd__a22o_1 \U$$1494  (.A1(net1588),
    .A2(net633),
    .B1(net1579),
    .B2(net906),
    .X(\t$5168 ));
 sky130_fd_sc_hd__xor2_1 \U$$1495  (.A(\t$5168 ),
    .B(net1491),
    .X(booth_b20_m59));
 sky130_fd_sc_hd__a22o_1 \U$$1496  (.A1(net1579),
    .A2(net633),
    .B1(net1553),
    .B2(net906),
    .X(\t$5169 ));
 sky130_fd_sc_hd__xor2_1 \U$$1497  (.A(\t$5169 ),
    .B(net1493),
    .X(booth_b20_m60));
 sky130_fd_sc_hd__a22o_1 \U$$1498  (.A1(net1553),
    .A2(net633),
    .B1(net1544),
    .B2(net906),
    .X(\t$5170 ));
 sky130_fd_sc_hd__xor2_1 \U$$1499  (.A(\t$5170 ),
    .B(net1493),
    .X(booth_b20_m61));
 sky130_fd_sc_hd__xor2_1 \U$$15  (.A(\t$4414 ),
    .B(net1573),
    .X(booth_b0_m4));
 sky130_fd_sc_hd__xor2_1 \U$$150  (.A(\t$4482 ),
    .B(net1390),
    .X(booth_b2_m3));
 sky130_fd_sc_hd__a22o_1 \U$$1500  (.A1(net1544),
    .A2(net633),
    .B1(net1536),
    .B2(net906),
    .X(\t$5171 ));
 sky130_fd_sc_hd__xor2_1 \U$$1501  (.A(\t$5171 ),
    .B(net1491),
    .X(booth_b20_m62));
 sky130_fd_sc_hd__a22o_1 \U$$1502  (.A1(net1536),
    .A2(net633),
    .B1(net1528),
    .B2(net906),
    .X(\t$5172 ));
 sky130_fd_sc_hd__xor2_1 \U$$1503  (.A(\t$5172 ),
    .B(net1491),
    .X(booth_b20_m63));
 sky130_fd_sc_hd__a22o_1 \U$$1504  (.A1(net1528),
    .A2(net633),
    .B1(net1762),
    .B2(net906),
    .X(\t$5173 ));
 sky130_fd_sc_hd__xor2_1 \U$$1505  (.A(\t$5173 ),
    .B(net1491),
    .X(booth_b20_m64));
 sky130_fd_sc_hd__inv_1 \U$$1506  (.A(net1491),
    .Y(\notsign$5174 ));
 sky130_fd_sc_hd__inv_1 \U$$1507  (.A(net1491),
    .Y(\notblock$5175[0] ));
 sky130_fd_sc_hd__inv_1 \U$$1508  (.A(net15),
    .Y(\notblock$5175[1] ));
 sky130_fd_sc_hd__inv_1 \U$$1509  (.A(net1481),
    .Y(\notblock$5175[2] ));
 sky130_fd_sc_hd__a22o_1 \U$$151  (.A1(net937),
    .A2(net624),
    .B1(net1675),
    .B2(net897),
    .X(\t$4483 ));
 sky130_fd_sc_hd__and2_1 \U$$1510  (.A(net1481),
    .B(\notblock$5175[1] ),
    .X(\t$5176 ));
 sky130_fd_sc_hd__a32o_4 \U$$1511  (.A1(\notblock$5175[2] ),
    .A2(net15),
    .A3(net1491),
    .B1(\t$5176 ),
    .B2(\notblock$5175[0] ),
    .X(\sel_0$5177 ));
 sky130_fd_sc_hd__xor2_4 \U$$1512  (.A(net15),
    .B(net1491),
    .X(\sel_1$5178 ));
 sky130_fd_sc_hd__a22o_1 \U$$1513  (.A1(net1763),
    .A2(net613),
    .B1(net1230),
    .B2(net886),
    .X(\t$5179 ));
 sky130_fd_sc_hd__xor2_1 \U$$1514  (.A(\t$5179 ),
    .B(net1478),
    .X(booth_b22_m0));
 sky130_fd_sc_hd__a22o_1 \U$$1515  (.A1(net1230),
    .A2(net613),
    .B1(net1126),
    .B2(net886),
    .X(\t$5180 ));
 sky130_fd_sc_hd__xor2_1 \U$$1516  (.A(\t$5180 ),
    .B(net1478),
    .X(booth_b22_m1));
 sky130_fd_sc_hd__a22o_1 \U$$1517  (.A1(net1123),
    .A2(net610),
    .B1(net1032),
    .B2(net883),
    .X(\t$5181 ));
 sky130_fd_sc_hd__xor2_1 \U$$1518  (.A(\t$5181 ),
    .B(net1475),
    .X(booth_b22_m2));
 sky130_fd_sc_hd__a22o_1 \U$$1519  (.A1(net1031),
    .A2(net611),
    .B1(net932),
    .B2(net884),
    .X(\t$5182 ));
 sky130_fd_sc_hd__xor2_1 \U$$152  (.A(\t$4483 ),
    .B(net1390),
    .X(booth_b2_m4));
 sky130_fd_sc_hd__xor2_1 \U$$1520  (.A(\t$5182 ),
    .B(net1475),
    .X(booth_b22_m3));
 sky130_fd_sc_hd__a22o_1 \U$$1521  (.A1(net932),
    .A2(net610),
    .B1(net1671),
    .B2(net883),
    .X(\t$5183 ));
 sky130_fd_sc_hd__xor2_1 \U$$1522  (.A(\t$5183 ),
    .B(net1475),
    .X(booth_b22_m4));
 sky130_fd_sc_hd__a22o_1 \U$$1523  (.A1(net1671),
    .A2(net610),
    .B1(net1560),
    .B2(net883),
    .X(\t$5184 ));
 sky130_fd_sc_hd__xor2_1 \U$$1524  (.A(\t$5184 ),
    .B(net1475),
    .X(booth_b22_m5));
 sky130_fd_sc_hd__a22o_1 \U$$1525  (.A1(net1560),
    .A2(net610),
    .B1(net1519),
    .B2(net883),
    .X(\t$5185 ));
 sky130_fd_sc_hd__xor2_1 \U$$1526  (.A(\t$5185 ),
    .B(net1475),
    .X(booth_b22_m6));
 sky130_fd_sc_hd__a22o_1 \U$$1527  (.A1(net1519),
    .A2(net610),
    .B1(net1511),
    .B2(net883),
    .X(\t$5186 ));
 sky130_fd_sc_hd__xor2_1 \U$$1528  (.A(\t$5186 ),
    .B(net1475),
    .X(booth_b22_m7));
 sky130_fd_sc_hd__a22o_1 \U$$1529  (.A1(net1511),
    .A2(net610),
    .B1(net1503),
    .B2(net883),
    .X(\t$5187 ));
 sky130_fd_sc_hd__a22o_1 \U$$153  (.A1(net1675),
    .A2(net624),
    .B1(net1565),
    .B2(net897),
    .X(\t$4484 ));
 sky130_fd_sc_hd__xor2_1 \U$$1530  (.A(\t$5187 ),
    .B(net1475),
    .X(booth_b22_m8));
 sky130_fd_sc_hd__a22o_1 \U$$1531  (.A1(net1503),
    .A2(net611),
    .B1(net1494),
    .B2(net884),
    .X(\t$5188 ));
 sky130_fd_sc_hd__xor2_1 \U$$1532  (.A(\t$5188 ),
    .B(net1476),
    .X(booth_b22_m9));
 sky130_fd_sc_hd__a22o_1 \U$$1533  (.A1(net1497),
    .A2(net613),
    .B1(net1221),
    .B2(net886),
    .X(\t$5189 ));
 sky130_fd_sc_hd__xor2_1 \U$$1534  (.A(\t$5189 ),
    .B(net1478),
    .X(booth_b22_m10));
 sky130_fd_sc_hd__a22o_1 \U$$1535  (.A1(net1224),
    .A2(net614),
    .B1(net1216),
    .B2(net887),
    .X(\t$5190 ));
 sky130_fd_sc_hd__xor2_1 \U$$1536  (.A(\t$5190 ),
    .B(net1479),
    .X(booth_b22_m11));
 sky130_fd_sc_hd__a22o_1 \U$$1537  (.A1(net1216),
    .A2(net613),
    .B1(net1206),
    .B2(net886),
    .X(\t$5191 ));
 sky130_fd_sc_hd__xor2_1 \U$$1538  (.A(\t$5191 ),
    .B(net1479),
    .X(booth_b22_m12));
 sky130_fd_sc_hd__a22o_1 \U$$1539  (.A1(net1206),
    .A2(net614),
    .B1(net1198),
    .B2(net887),
    .X(\t$5192 ));
 sky130_fd_sc_hd__xor2_1 \U$$154  (.A(\t$4484 ),
    .B(net1390),
    .X(booth_b2_m5));
 sky130_fd_sc_hd__xor2_1 \U$$1540  (.A(\t$5192 ),
    .B(net1479),
    .X(booth_b22_m13));
 sky130_fd_sc_hd__a22o_1 \U$$1541  (.A1(net1198),
    .A2(net613),
    .B1(net1179),
    .B2(net886),
    .X(\t$5193 ));
 sky130_fd_sc_hd__xor2_1 \U$$1542  (.A(\t$5193 ),
    .B(net1478),
    .X(booth_b22_m14));
 sky130_fd_sc_hd__a22o_1 \U$$1543  (.A1(net1179),
    .A2(net613),
    .B1(net1170),
    .B2(net886),
    .X(\t$5194 ));
 sky130_fd_sc_hd__xor2_1 \U$$1544  (.A(\t$5194 ),
    .B(net1478),
    .X(booth_b22_m15));
 sky130_fd_sc_hd__a22o_1 \U$$1545  (.A1(net1166),
    .A2(net613),
    .B1(net1157),
    .B2(net886),
    .X(\t$5195 ));
 sky130_fd_sc_hd__xor2_1 \U$$1546  (.A(\t$5195 ),
    .B(net1478),
    .X(booth_b22_m16));
 sky130_fd_sc_hd__a22o_1 \U$$1547  (.A1(net1157),
    .A2(net610),
    .B1(net1147),
    .B2(net883),
    .X(\t$5196 ));
 sky130_fd_sc_hd__xor2_1 \U$$1548  (.A(\t$5196 ),
    .B(net1476),
    .X(booth_b22_m17));
 sky130_fd_sc_hd__a22o_1 \U$$1549  (.A1(net1146),
    .A2(net611),
    .B1(net1139),
    .B2(net884),
    .X(\t$5197 ));
 sky130_fd_sc_hd__a22o_1 \U$$155  (.A1(net1564),
    .A2(net624),
    .B1(net1523),
    .B2(net897),
    .X(\t$4485 ));
 sky130_fd_sc_hd__xor2_1 \U$$1550  (.A(\t$5197 ),
    .B(net1476),
    .X(booth_b22_m18));
 sky130_fd_sc_hd__a22o_1 \U$$1551  (.A1(net1138),
    .A2(net610),
    .B1(net1130),
    .B2(net883),
    .X(\t$5198 ));
 sky130_fd_sc_hd__xor2_1 \U$$1552  (.A(\t$5198 ),
    .B(net1475),
    .X(booth_b22_m19));
 sky130_fd_sc_hd__a22o_1 \U$$1553  (.A1(net1132),
    .A2(net610),
    .B1(net1116),
    .B2(net883),
    .X(\t$5199 ));
 sky130_fd_sc_hd__xor2_1 \U$$1554  (.A(\t$5199 ),
    .B(net1475),
    .X(booth_b22_m20));
 sky130_fd_sc_hd__a22o_1 \U$$1555  (.A1(net1114),
    .A2(net610),
    .B1(net1105),
    .B2(net883),
    .X(\t$5200 ));
 sky130_fd_sc_hd__xor2_1 \U$$1556  (.A(\t$5200 ),
    .B(net1475),
    .X(booth_b22_m21));
 sky130_fd_sc_hd__a22o_1 \U$$1557  (.A1(net1107),
    .A2(net612),
    .B1(net1098),
    .B2(net885),
    .X(\t$5201 ));
 sky130_fd_sc_hd__xor2_1 \U$$1558  (.A(\t$5201 ),
    .B(net1477),
    .X(booth_b22_m22));
 sky130_fd_sc_hd__a22o_1 \U$$1559  (.A1(net1099),
    .A2(net611),
    .B1(net1089),
    .B2(net884),
    .X(\t$5202 ));
 sky130_fd_sc_hd__xor2_1 \U$$156  (.A(\t$4485 ),
    .B(net1390),
    .X(booth_b2_m6));
 sky130_fd_sc_hd__xor2_1 \U$$1560  (.A(\t$5202 ),
    .B(net1476),
    .X(booth_b22_m23));
 sky130_fd_sc_hd__a22o_1 \U$$1561  (.A1(net1089),
    .A2(net611),
    .B1(net1081),
    .B2(net884),
    .X(\t$5203 ));
 sky130_fd_sc_hd__xor2_1 \U$$1562  (.A(\t$5203 ),
    .B(net1476),
    .X(booth_b22_m24));
 sky130_fd_sc_hd__a22o_1 \U$$1563  (.A1(net1082),
    .A2(net612),
    .B1(net1073),
    .B2(net885),
    .X(\t$5204 ));
 sky130_fd_sc_hd__xor2_1 \U$$1564  (.A(\t$5204 ),
    .B(net1477),
    .X(booth_b22_m25));
 sky130_fd_sc_hd__a22o_1 \U$$1565  (.A1(net1073),
    .A2(net612),
    .B1(net1064),
    .B2(net885),
    .X(\t$5205 ));
 sky130_fd_sc_hd__xor2_1 \U$$1566  (.A(\t$5205 ),
    .B(net1477),
    .X(booth_b22_m26));
 sky130_fd_sc_hd__a22o_1 \U$$1567  (.A1(net1064),
    .A2(net612),
    .B1(net1056),
    .B2(net885),
    .X(\t$5206 ));
 sky130_fd_sc_hd__xor2_1 \U$$1568  (.A(\t$5206 ),
    .B(net1477),
    .X(booth_b22_m27));
 sky130_fd_sc_hd__a22o_1 \U$$1569  (.A1(net1057),
    .A2(net613),
    .B1(net1049),
    .B2(net886),
    .X(\t$5207 ));
 sky130_fd_sc_hd__a22o_1 \U$$157  (.A1(net1523),
    .A2(net624),
    .B1(net1515),
    .B2(net897),
    .X(\t$4486 ));
 sky130_fd_sc_hd__xor2_1 \U$$1570  (.A(\t$5207 ),
    .B(net1478),
    .X(booth_b22_m28));
 sky130_fd_sc_hd__a22o_1 \U$$1571  (.A1(net1049),
    .A2(net615),
    .B1(net1041),
    .B2(net888),
    .X(\t$5208 ));
 sky130_fd_sc_hd__xor2_1 \U$$1572  (.A(\t$5208 ),
    .B(net1480),
    .X(booth_b22_m29));
 sky130_fd_sc_hd__a22o_1 \U$$1573  (.A1(net1041),
    .A2(net614),
    .B1(net1025),
    .B2(net887),
    .X(\t$5209 ));
 sky130_fd_sc_hd__xor2_1 \U$$1574  (.A(\t$5209 ),
    .B(net1479),
    .X(booth_b22_m30));
 sky130_fd_sc_hd__a22o_1 \U$$1575  (.A1(net1025),
    .A2(net614),
    .B1(net1017),
    .B2(net887),
    .X(\t$5210 ));
 sky130_fd_sc_hd__xor2_1 \U$$1576  (.A(\t$5210 ),
    .B(net1479),
    .X(booth_b22_m31));
 sky130_fd_sc_hd__a22o_1 \U$$1577  (.A1(net1018),
    .A2(net614),
    .B1(net1001),
    .B2(net887),
    .X(\t$5211 ));
 sky130_fd_sc_hd__xor2_1 \U$$1578  (.A(\t$5211 ),
    .B(net1479),
    .X(booth_b22_m32));
 sky130_fd_sc_hd__a22o_1 \U$$1579  (.A1(net1001),
    .A2(net614),
    .B1(net993),
    .B2(net887),
    .X(\t$5212 ));
 sky130_fd_sc_hd__xor2_1 \U$$158  (.A(\t$4486 ),
    .B(net1390),
    .X(booth_b2_m7));
 sky130_fd_sc_hd__xor2_1 \U$$1580  (.A(\t$5212 ),
    .B(net1479),
    .X(booth_b22_m33));
 sky130_fd_sc_hd__a22o_1 \U$$1581  (.A1(net992),
    .A2(net613),
    .B1(net987),
    .B2(net886),
    .X(\t$5213 ));
 sky130_fd_sc_hd__xor2_1 \U$$1582  (.A(\t$5213 ),
    .B(net1478),
    .X(booth_b22_m34));
 sky130_fd_sc_hd__a22o_1 \U$$1583  (.A1(net987),
    .A2(net613),
    .B1(net977),
    .B2(net886),
    .X(\t$5214 ));
 sky130_fd_sc_hd__xor2_1 \U$$1584  (.A(\t$5214 ),
    .B(net1478),
    .X(booth_b22_m35));
 sky130_fd_sc_hd__a22o_1 \U$$1585  (.A1(net977),
    .A2(net618),
    .B1(net965),
    .B2(net891),
    .X(\t$5215 ));
 sky130_fd_sc_hd__xor2_1 \U$$1586  (.A(\t$5215 ),
    .B(net1484),
    .X(booth_b22_m36));
 sky130_fd_sc_hd__a22o_1 \U$$1587  (.A1(net965),
    .A2(net615),
    .B1(net957),
    .B2(net888),
    .X(\t$5216 ));
 sky130_fd_sc_hd__xor2_1 \U$$1588  (.A(\t$5216 ),
    .B(net1480),
    .X(booth_b22_m37));
 sky130_fd_sc_hd__a22o_1 \U$$1589  (.A1(net957),
    .A2(net612),
    .B1(net949),
    .B2(net885),
    .X(\t$5217 ));
 sky130_fd_sc_hd__a22o_1 \U$$159  (.A1(net1515),
    .A2(net623),
    .B1(net1508),
    .B2(net896),
    .X(\t$4487 ));
 sky130_fd_sc_hd__xor2_1 \U$$1590  (.A(\t$5217 ),
    .B(net1477),
    .X(booth_b22_m38));
 sky130_fd_sc_hd__a22o_1 \U$$1591  (.A1(net948),
    .A2(net612),
    .B1(net941),
    .B2(net885),
    .X(\t$5218 ));
 sky130_fd_sc_hd__xor2_1 \U$$1592  (.A(\t$5218 ),
    .B(net1477),
    .X(booth_b22_m39));
 sky130_fd_sc_hd__a22o_1 \U$$1593  (.A1(net940),
    .A2(net612),
    .B1(net924),
    .B2(net885),
    .X(\t$5219 ));
 sky130_fd_sc_hd__xor2_1 \U$$1594  (.A(\t$5219 ),
    .B(net1477),
    .X(booth_b22_m40));
 sky130_fd_sc_hd__a22o_1 \U$$1595  (.A1(net925),
    .A2(net616),
    .B1(net1746),
    .B2(net889),
    .X(\t$5220 ));
 sky130_fd_sc_hd__xor2_1 \U$$1596  (.A(\t$5220 ),
    .B(net1483),
    .X(booth_b22_m41));
 sky130_fd_sc_hd__a22o_1 \U$$1597  (.A1(net1749),
    .A2(net618),
    .B1(net1741),
    .B2(net891),
    .X(\t$5221 ));
 sky130_fd_sc_hd__xor2_1 \U$$1598  (.A(\t$5221 ),
    .B(net1484),
    .X(booth_b22_m42));
 sky130_fd_sc_hd__a22o_1 \U$$1599  (.A1(net1741),
    .A2(net615),
    .B1(net1733),
    .B2(net888),
    .X(\t$5222 ));
 sky130_fd_sc_hd__a22o_1 \U$$16  (.A1(net1675),
    .A2(net446),
    .B1(net1565),
    .B2(net688),
    .X(\t$4415 ));
 sky130_fd_sc_hd__xor2_1 \U$$160  (.A(\t$4487 ),
    .B(net1389),
    .X(booth_b2_m8));
 sky130_fd_sc_hd__xor2_1 \U$$1600  (.A(\t$5222 ),
    .B(net1480),
    .X(booth_b22_m43));
 sky130_fd_sc_hd__a22o_1 \U$$1601  (.A1(net1733),
    .A2(net615),
    .B1(net1724),
    .B2(net888),
    .X(\t$5223 ));
 sky130_fd_sc_hd__xor2_1 \U$$1602  (.A(\t$5223 ),
    .B(net1480),
    .X(booth_b22_m44));
 sky130_fd_sc_hd__a22o_1 \U$$1603  (.A1(net1727),
    .A2(net618),
    .B1(net1719),
    .B2(net891),
    .X(\t$5224 ));
 sky130_fd_sc_hd__xor2_1 \U$$1604  (.A(\t$5224 ),
    .B(net1484),
    .X(booth_b22_m45));
 sky130_fd_sc_hd__a22o_1 \U$$1605  (.A1(net1719),
    .A2(net618),
    .B1(net1710),
    .B2(net891),
    .X(\t$5225 ));
 sky130_fd_sc_hd__xor2_1 \U$$1606  (.A(\t$5225 ),
    .B(net1484),
    .X(booth_b22_m46));
 sky130_fd_sc_hd__a22o_1 \U$$1607  (.A1(net1706),
    .A2(net618),
    .B1(net1698),
    .B2(net891),
    .X(\t$5226 ));
 sky130_fd_sc_hd__xor2_1 \U$$1608  (.A(\t$5226 ),
    .B(net1484),
    .X(booth_b22_m47));
 sky130_fd_sc_hd__a22o_1 \U$$1609  (.A1(net1698),
    .A2(net618),
    .B1(net1690),
    .B2(net891),
    .X(\t$5227 ));
 sky130_fd_sc_hd__a22o_1 \U$$161  (.A1(net1508),
    .A2(net624),
    .B1(net1499),
    .B2(net897),
    .X(\t$4488 ));
 sky130_fd_sc_hd__xor2_1 \U$$1610  (.A(\t$5227 ),
    .B(net1484),
    .X(booth_b22_m48));
 sky130_fd_sc_hd__a22o_1 \U$$1611  (.A1(net1687),
    .A2(net616),
    .B1(net1679),
    .B2(net889),
    .X(\t$5228 ));
 sky130_fd_sc_hd__xor2_1 \U$$1612  (.A(\t$5228 ),
    .B(net1483),
    .X(booth_b22_m49));
 sky130_fd_sc_hd__a22o_1 \U$$1613  (.A1(net1681),
    .A2(net616),
    .B1(net1654),
    .B2(net889),
    .X(\t$5229 ));
 sky130_fd_sc_hd__xor2_1 \U$$1614  (.A(\t$5229 ),
    .B(net1483),
    .X(booth_b22_m50));
 sky130_fd_sc_hd__a22o_1 \U$$1615  (.A1(net1654),
    .A2(net616),
    .B1(net1646),
    .B2(net889),
    .X(\t$5230 ));
 sky130_fd_sc_hd__xor2_1 \U$$1616  (.A(\t$5230 ),
    .B(net1483),
    .X(booth_b22_m51));
 sky130_fd_sc_hd__a22o_1 \U$$1617  (.A1(net1646),
    .A2(net616),
    .B1(net1638),
    .B2(net889),
    .X(\t$5231 ));
 sky130_fd_sc_hd__xor2_1 \U$$1618  (.A(\t$5231 ),
    .B(net1483),
    .X(booth_b22_m52));
 sky130_fd_sc_hd__a22o_1 \U$$1619  (.A1(net1638),
    .A2(net616),
    .B1(net1629),
    .B2(net889),
    .X(\t$5232 ));
 sky130_fd_sc_hd__xor2_1 \U$$162  (.A(\t$4488 ),
    .B(net1390),
    .X(booth_b2_m9));
 sky130_fd_sc_hd__xor2_1 \U$$1620  (.A(\t$5232 ),
    .B(net1483),
    .X(booth_b22_m53));
 sky130_fd_sc_hd__a22o_1 \U$$1621  (.A1(net1629),
    .A2(net616),
    .B1(net1621),
    .B2(net889),
    .X(\t$5233 ));
 sky130_fd_sc_hd__xor2_1 \U$$1622  (.A(\t$5233 ),
    .B(net1483),
    .X(booth_b22_m54));
 sky130_fd_sc_hd__a22o_1 \U$$1623  (.A1(net1621),
    .A2(net616),
    .B1(net1614),
    .B2(net889),
    .X(\t$5234 ));
 sky130_fd_sc_hd__xor2_1 \U$$1624  (.A(\t$5234 ),
    .B(net1483),
    .X(booth_b22_m55));
 sky130_fd_sc_hd__a22o_1 \U$$1625  (.A1(net1614),
    .A2(net616),
    .B1(net1606),
    .B2(net889),
    .X(\t$5235 ));
 sky130_fd_sc_hd__xor2_1 \U$$1626  (.A(\t$5235 ),
    .B(net1483),
    .X(booth_b22_m56));
 sky130_fd_sc_hd__a22o_1 \U$$1627  (.A1(net1605),
    .A2(net617),
    .B1(net1597),
    .B2(net890),
    .X(\t$5236 ));
 sky130_fd_sc_hd__xor2_1 \U$$1628  (.A(\t$5236 ),
    .B(net1481),
    .X(booth_b22_m57));
 sky130_fd_sc_hd__a22o_1 \U$$1629  (.A1(net1597),
    .A2(net616),
    .B1(net1588),
    .B2(net889),
    .X(\t$5237 ));
 sky130_fd_sc_hd__a22o_1 \U$$163  (.A1(net1499),
    .A2(net624),
    .B1(net1224),
    .B2(net897),
    .X(\t$4489 ));
 sky130_fd_sc_hd__xor2_1 \U$$1630  (.A(\t$5237 ),
    .B(net1482),
    .X(booth_b22_m58));
 sky130_fd_sc_hd__a22o_1 \U$$1631  (.A1(net1588),
    .A2(net617),
    .B1(net1579),
    .B2(net890),
    .X(\t$5238 ));
 sky130_fd_sc_hd__xor2_1 \U$$1632  (.A(\t$5238 ),
    .B(net1482),
    .X(booth_b22_m59));
 sky130_fd_sc_hd__a22o_1 \U$$1633  (.A1(net1579),
    .A2(net617),
    .B1(net1553),
    .B2(net890),
    .X(\t$5239 ));
 sky130_fd_sc_hd__xor2_1 \U$$1634  (.A(\t$5239 ),
    .B(net1481),
    .X(booth_b22_m60));
 sky130_fd_sc_hd__a22o_1 \U$$1635  (.A1(net1553),
    .A2(net617),
    .B1(net1544),
    .B2(net890),
    .X(\t$5240 ));
 sky130_fd_sc_hd__xor2_1 \U$$1636  (.A(\t$5240 ),
    .B(net1481),
    .X(booth_b22_m61));
 sky130_fd_sc_hd__a22o_1 \U$$1637  (.A1(net1544),
    .A2(net617),
    .B1(net1536),
    .B2(net890),
    .X(\t$5241 ));
 sky130_fd_sc_hd__xor2_1 \U$$1638  (.A(\t$5241 ),
    .B(net1481),
    .X(booth_b22_m62));
 sky130_fd_sc_hd__a22o_1 \U$$1639  (.A1(net1536),
    .A2(net617),
    .B1(net1528),
    .B2(net890),
    .X(\t$5242 ));
 sky130_fd_sc_hd__xor2_1 \U$$164  (.A(\t$4489 ),
    .B(net1390),
    .X(booth_b2_m10));
 sky130_fd_sc_hd__xor2_1 \U$$1640  (.A(\t$5242 ),
    .B(net1481),
    .X(booth_b22_m63));
 sky130_fd_sc_hd__a22o_1 \U$$1641  (.A1(net1528),
    .A2(net617),
    .B1(net1764),
    .B2(net890),
    .X(\t$5243 ));
 sky130_fd_sc_hd__xor2_1 \U$$1642  (.A(\t$5243 ),
    .B(net1481),
    .X(booth_b22_m64));
 sky130_fd_sc_hd__inv_1 \U$$1643  (.A(net1481),
    .Y(\notsign$5244 ));
 sky130_fd_sc_hd__inv_1 \U$$1644  (.A(net1481),
    .Y(\notblock$5245[0] ));
 sky130_fd_sc_hd__inv_1 \U$$1645  (.A(net17),
    .Y(\notblock$5245[1] ));
 sky130_fd_sc_hd__inv_1 \U$$1646  (.A(net1471),
    .Y(\notblock$5245[2] ));
 sky130_fd_sc_hd__and2_1 \U$$1647  (.A(net1471),
    .B(\notblock$5245[1] ),
    .X(\t$5246 ));
 sky130_fd_sc_hd__a32o_4 \U$$1648  (.A1(\notblock$5245[2] ),
    .A2(net17),
    .A3(net1482),
    .B1(\t$5246 ),
    .B2(\notblock$5245[0] ),
    .X(\sel_0$5247 ));
 sky130_fd_sc_hd__xor2_4 \U$$1649  (.A(net17),
    .B(net1482),
    .X(\sel_1$5248 ));
 sky130_fd_sc_hd__a22o_1 \U$$165  (.A1(net1224),
    .A2(net625),
    .B1(net1216),
    .B2(net898),
    .X(\t$4490 ));
 sky130_fd_sc_hd__a22o_1 \U$$1650  (.A1(net1765),
    .A2(net603),
    .B1(net1228),
    .B2(net876),
    .X(\t$5249 ));
 sky130_fd_sc_hd__xor2_1 \U$$1651  (.A(\t$5249 ),
    .B(net1466),
    .X(booth_b24_m0));
 sky130_fd_sc_hd__a22o_1 \U$$1652  (.A1(net1228),
    .A2(net602),
    .B1(net1122),
    .B2(net875),
    .X(\t$5250 ));
 sky130_fd_sc_hd__xor2_1 \U$$1653  (.A(\t$5250 ),
    .B(net1466),
    .X(booth_b24_m1));
 sky130_fd_sc_hd__a22o_1 \U$$1654  (.A1(net1123),
    .A2(net603),
    .B1(net1032),
    .B2(net876),
    .X(\t$5251 ));
 sky130_fd_sc_hd__xor2_1 \U$$1655  (.A(\t$5251 ),
    .B(net1467),
    .X(booth_b24_m2));
 sky130_fd_sc_hd__a22o_1 \U$$1656  (.A1(net1031),
    .A2(net602),
    .B1(net932),
    .B2(net875),
    .X(\t$5252 ));
 sky130_fd_sc_hd__xor2_1 \U$$1657  (.A(\t$5252 ),
    .B(net1466),
    .X(booth_b24_m3));
 sky130_fd_sc_hd__a22o_1 \U$$1658  (.A1(net932),
    .A2(net602),
    .B1(net1671),
    .B2(net875),
    .X(\t$5253 ));
 sky130_fd_sc_hd__xor2_1 \U$$1659  (.A(\t$5253 ),
    .B(net1466),
    .X(booth_b24_m4));
 sky130_fd_sc_hd__xor2_1 \U$$166  (.A(\t$4490 ),
    .B(net1391),
    .X(booth_b2_m11));
 sky130_fd_sc_hd__a22o_1 \U$$1660  (.A1(net1671),
    .A2(net602),
    .B1(net1560),
    .B2(net875),
    .X(\t$5254 ));
 sky130_fd_sc_hd__xor2_1 \U$$1661  (.A(\t$5254 ),
    .B(net1466),
    .X(booth_b24_m5));
 sky130_fd_sc_hd__a22o_1 \U$$1662  (.A1(net1560),
    .A2(net602),
    .B1(net1519),
    .B2(net875),
    .X(\t$5255 ));
 sky130_fd_sc_hd__xor2_1 \U$$1663  (.A(\t$5255 ),
    .B(net1466),
    .X(booth_b24_m6));
 sky130_fd_sc_hd__a22o_1 \U$$1664  (.A1(net1519),
    .A2(net602),
    .B1(net1511),
    .B2(net875),
    .X(\t$5256 ));
 sky130_fd_sc_hd__xor2_1 \U$$1665  (.A(\t$5256 ),
    .B(net1466),
    .X(booth_b24_m7));
 sky130_fd_sc_hd__a22o_1 \U$$1666  (.A1(net1515),
    .A2(net605),
    .B1(net1508),
    .B2(net878),
    .X(\t$5257 ));
 sky130_fd_sc_hd__xor2_1 \U$$1667  (.A(\t$5257 ),
    .B(net1469),
    .X(booth_b24_m8));
 sky130_fd_sc_hd__a22o_1 \U$$1668  (.A1(net1509),
    .A2(net605),
    .B1(net1499),
    .B2(net878),
    .X(\t$5258 ));
 sky130_fd_sc_hd__xor2_1 \U$$1669  (.A(\t$5258 ),
    .B(net1469),
    .X(booth_b24_m9));
 sky130_fd_sc_hd__a22o_1 \U$$167  (.A1(net1211),
    .A2(net623),
    .B1(net1203),
    .B2(net896),
    .X(\t$4491 ));
 sky130_fd_sc_hd__a22o_1 \U$$1670  (.A1(net1500),
    .A2(net605),
    .B1(net1225),
    .B2(net878),
    .X(\t$5259 ));
 sky130_fd_sc_hd__xor2_1 \U$$1671  (.A(\t$5259 ),
    .B(net1469),
    .X(booth_b24_m10));
 sky130_fd_sc_hd__a22o_1 \U$$1672  (.A1(net1225),
    .A2(net605),
    .B1(net1216),
    .B2(net878),
    .X(\t$5260 ));
 sky130_fd_sc_hd__xor2_1 \U$$1673  (.A(\t$5260 ),
    .B(net1469),
    .X(booth_b24_m11));
 sky130_fd_sc_hd__a22o_1 \U$$1674  (.A1(net1216),
    .A2(net606),
    .B1(net1206),
    .B2(net879),
    .X(\t$5261 ));
 sky130_fd_sc_hd__xor2_1 \U$$1675  (.A(\t$5261 ),
    .B(net1469),
    .X(booth_b24_m12));
 sky130_fd_sc_hd__a22o_1 \U$$1676  (.A1(net1206),
    .A2(net605),
    .B1(net1198),
    .B2(net878),
    .X(\t$5262 ));
 sky130_fd_sc_hd__xor2_1 \U$$1677  (.A(\t$5262 ),
    .B(net1469),
    .X(booth_b24_m13));
 sky130_fd_sc_hd__a22o_1 \U$$1678  (.A1(net1194),
    .A2(net605),
    .B1(net1175),
    .B2(net878),
    .X(\t$5263 ));
 sky130_fd_sc_hd__xor2_1 \U$$1679  (.A(\t$5263 ),
    .B(net1469),
    .X(booth_b24_m14));
 sky130_fd_sc_hd__xor2_1 \U$$168  (.A(\t$4491 ),
    .B(net1389),
    .X(booth_b2_m12));
 sky130_fd_sc_hd__a22o_1 \U$$1680  (.A1(net1175),
    .A2(net603),
    .B1(net1166),
    .B2(net876),
    .X(\t$5264 ));
 sky130_fd_sc_hd__xor2_1 \U$$1681  (.A(\t$5264 ),
    .B(net1467),
    .X(booth_b24_m15));
 sky130_fd_sc_hd__a22o_1 \U$$1682  (.A1(net1164),
    .A2(net603),
    .B1(net1155),
    .B2(net876),
    .X(\t$5265 ));
 sky130_fd_sc_hd__xor2_1 \U$$1683  (.A(\t$5265 ),
    .B(net1467),
    .X(booth_b24_m16));
 sky130_fd_sc_hd__a22o_1 \U$$1684  (.A1(net1155),
    .A2(net602),
    .B1(net1146),
    .B2(net875),
    .X(\t$5266 ));
 sky130_fd_sc_hd__xor2_1 \U$$1685  (.A(\t$5266 ),
    .B(net1466),
    .X(booth_b24_m17));
 sky130_fd_sc_hd__a22o_1 \U$$1686  (.A1(net1147),
    .A2(net602),
    .B1(net1138),
    .B2(net875),
    .X(\t$5267 ));
 sky130_fd_sc_hd__xor2_1 \U$$1687  (.A(\t$5267 ),
    .B(net1466),
    .X(booth_b24_m18));
 sky130_fd_sc_hd__a22o_1 \U$$1688  (.A1(net1138),
    .A2(net602),
    .B1(net1130),
    .B2(net875),
    .X(\t$5268 ));
 sky130_fd_sc_hd__xor2_1 \U$$1689  (.A(\t$5268 ),
    .B(net1466),
    .X(booth_b24_m19));
 sky130_fd_sc_hd__a22o_1 \U$$169  (.A1(net1203),
    .A2(net620),
    .B1(net1194),
    .B2(net893),
    .X(\t$4492 ));
 sky130_fd_sc_hd__a22o_1 \U$$1690  (.A1(net1131),
    .A2(net603),
    .B1(net1115),
    .B2(net876),
    .X(\t$5269 ));
 sky130_fd_sc_hd__xor2_1 \U$$1691  (.A(\t$5269 ),
    .B(net1467),
    .X(booth_b24_m20));
 sky130_fd_sc_hd__a22o_1 \U$$1692  (.A1(net1116),
    .A2(net603),
    .B1(net1106),
    .B2(net876),
    .X(\t$5270 ));
 sky130_fd_sc_hd__xor2_1 \U$$1693  (.A(\t$5270 ),
    .B(net1467),
    .X(booth_b24_m21));
 sky130_fd_sc_hd__a22o_1 \U$$1694  (.A1(net1107),
    .A2(net603),
    .B1(net1098),
    .B2(net876),
    .X(\t$5271 ));
 sky130_fd_sc_hd__xor2_1 \U$$1695  (.A(\t$5271 ),
    .B(net1467),
    .X(booth_b24_m22));
 sky130_fd_sc_hd__a22o_1 \U$$1696  (.A1(net1098),
    .A2(net604),
    .B1(net1090),
    .B2(net877),
    .X(\t$5272 ));
 sky130_fd_sc_hd__xor2_1 \U$$1697  (.A(\t$5272 ),
    .B(net1468),
    .X(booth_b24_m23));
 sky130_fd_sc_hd__a22o_1 \U$$1698  (.A1(net1090),
    .A2(net604),
    .B1(net1082),
    .B2(net877),
    .X(\t$5273 ));
 sky130_fd_sc_hd__xor2_1 \U$$1699  (.A(\t$5273 ),
    .B(net1468),
    .X(booth_b24_m24));
 sky130_fd_sc_hd__xor2_1 \U$$17  (.A(\t$4415 ),
    .B(net1573),
    .X(booth_b0_m5));
 sky130_fd_sc_hd__xor2_1 \U$$170  (.A(\t$4492 ),
    .B(net1386),
    .X(booth_b2_m13));
 sky130_fd_sc_hd__a22o_1 \U$$1700  (.A1(net1082),
    .A2(net602),
    .B1(net1073),
    .B2(net875),
    .X(\t$5274 ));
 sky130_fd_sc_hd__xor2_1 \U$$1701  (.A(\t$5274 ),
    .B(net1468),
    .X(booth_b24_m25));
 sky130_fd_sc_hd__a22o_1 \U$$1702  (.A1(net1073),
    .A2(net604),
    .B1(net1064),
    .B2(net877),
    .X(\t$5275 ));
 sky130_fd_sc_hd__xor2_1 \U$$1703  (.A(\t$5275 ),
    .B(net1468),
    .X(booth_b24_m26));
 sky130_fd_sc_hd__a22o_1 \U$$1704  (.A1(net1066),
    .A2(net605),
    .B1(net1057),
    .B2(net878),
    .X(\t$5276 ));
 sky130_fd_sc_hd__xor2_1 \U$$1705  (.A(\t$5276 ),
    .B(net1469),
    .X(booth_b24_m27));
 sky130_fd_sc_hd__a22o_1 \U$$1706  (.A1(net1057),
    .A2(net605),
    .B1(net1049),
    .B2(net878),
    .X(\t$5277 ));
 sky130_fd_sc_hd__xor2_1 \U$$1707  (.A(\t$5277 ),
    .B(net1469),
    .X(booth_b24_m28));
 sky130_fd_sc_hd__a22o_1 \U$$1708  (.A1(net1049),
    .A2(net605),
    .B1(net1041),
    .B2(net878),
    .X(\t$5278 ));
 sky130_fd_sc_hd__xor2_1 \U$$1709  (.A(\t$5278 ),
    .B(net1470),
    .X(booth_b24_m29));
 sky130_fd_sc_hd__a22o_1 \U$$171  (.A1(net1194),
    .A2(net620),
    .B1(net1175),
    .B2(net893),
    .X(\t$4493 ));
 sky130_fd_sc_hd__a22o_1 \U$$1710  (.A1(net1041),
    .A2(net606),
    .B1(net1026),
    .B2(net879),
    .X(\t$5279 ));
 sky130_fd_sc_hd__xor2_1 \U$$1711  (.A(\t$5279 ),
    .B(net1470),
    .X(booth_b24_m30));
 sky130_fd_sc_hd__a22o_1 \U$$1712  (.A1(net1026),
    .A2(net606),
    .B1(net1018),
    .B2(net879),
    .X(\t$5280 ));
 sky130_fd_sc_hd__xor2_1 \U$$1713  (.A(\t$5280 ),
    .B(net1470),
    .X(booth_b24_m31));
 sky130_fd_sc_hd__a22o_1 \U$$1714  (.A1(net1017),
    .A2(net606),
    .B1(net1000),
    .B2(net879),
    .X(\t$5281 ));
 sky130_fd_sc_hd__xor2_1 \U$$1715  (.A(\t$5281 ),
    .B(net1470),
    .X(booth_b24_m32));
 sky130_fd_sc_hd__a22o_1 \U$$1716  (.A1(net1000),
    .A2(net605),
    .B1(net992),
    .B2(net878),
    .X(\t$5282 ));
 sky130_fd_sc_hd__xor2_1 \U$$1717  (.A(\t$5282 ),
    .B(net1469),
    .X(booth_b24_m33));
 sky130_fd_sc_hd__a22o_1 \U$$1718  (.A1(net996),
    .A2(net609),
    .B1(net988),
    .B2(net882),
    .X(\t$5283 ));
 sky130_fd_sc_hd__xor2_1 \U$$1719  (.A(\t$5283 ),
    .B(net1474),
    .X(booth_b24_m34));
 sky130_fd_sc_hd__xor2_1 \U$$172  (.A(\t$4493 ),
    .B(net1386),
    .X(booth_b2_m14));
 sky130_fd_sc_hd__a22o_1 \U$$1720  (.A1(net983),
    .A2(net604),
    .B1(net974),
    .B2(net877),
    .X(\t$5284 ));
 sky130_fd_sc_hd__xor2_1 \U$$1721  (.A(\t$5284 ),
    .B(net1468),
    .X(booth_b24_m35));
 sky130_fd_sc_hd__a22o_1 \U$$1722  (.A1(net974),
    .A2(net606),
    .B1(net965),
    .B2(net879),
    .X(\t$5285 ));
 sky130_fd_sc_hd__xor2_1 \U$$1723  (.A(\t$5285 ),
    .B(net1470),
    .X(booth_b24_m36));
 sky130_fd_sc_hd__a22o_1 \U$$1724  (.A1(net965),
    .A2(net604),
    .B1(net957),
    .B2(net877),
    .X(\t$5286 ));
 sky130_fd_sc_hd__xor2_1 \U$$1725  (.A(\t$5286 ),
    .B(net1468),
    .X(booth_b24_m37));
 sky130_fd_sc_hd__a22o_1 \U$$1726  (.A1(net957),
    .A2(net604),
    .B1(net948),
    .B2(net877),
    .X(\t$5287 ));
 sky130_fd_sc_hd__xor2_1 \U$$1727  (.A(\t$5287 ),
    .B(net1468),
    .X(booth_b24_m38));
 sky130_fd_sc_hd__a22o_1 \U$$1728  (.A1(net949),
    .A2(net607),
    .B1(net941),
    .B2(net880),
    .X(\t$5288 ));
 sky130_fd_sc_hd__xor2_1 \U$$1729  (.A(\t$5288 ),
    .B(net1473),
    .X(booth_b24_m39));
 sky130_fd_sc_hd__a22o_1 \U$$173  (.A1(net1175),
    .A2(net620),
    .B1(net1166),
    .B2(net893),
    .X(\t$4494 ));
 sky130_fd_sc_hd__a22o_1 \U$$1730  (.A1(net944),
    .A2(net606),
    .B1(net928),
    .B2(net879),
    .X(\t$5289 ));
 sky130_fd_sc_hd__xor2_1 \U$$1731  (.A(\t$5289 ),
    .B(net1470),
    .X(booth_b24_m40));
 sky130_fd_sc_hd__a22o_1 \U$$1732  (.A1(net928),
    .A2(net609),
    .B1(net1749),
    .B2(net882),
    .X(\t$5290 ));
 sky130_fd_sc_hd__xor2_1 \U$$1733  (.A(\t$5290 ),
    .B(net1474),
    .X(booth_b24_m41));
 sky130_fd_sc_hd__a22o_1 \U$$1734  (.A1(net1749),
    .A2(net606),
    .B1(net1741),
    .B2(net879),
    .X(\t$5291 ));
 sky130_fd_sc_hd__xor2_1 \U$$1735  (.A(\t$5291 ),
    .B(net1470),
    .X(booth_b24_m42));
 sky130_fd_sc_hd__a22o_1 \U$$1736  (.A1(net1743),
    .A2(net609),
    .B1(net1735),
    .B2(net882),
    .X(\t$5292 ));
 sky130_fd_sc_hd__xor2_1 \U$$1737  (.A(\t$5292 ),
    .B(net1474),
    .X(booth_b24_m43));
 sky130_fd_sc_hd__a22o_1 \U$$1738  (.A1(net1735),
    .A2(net609),
    .B1(net1727),
    .B2(net882),
    .X(\t$5293 ));
 sky130_fd_sc_hd__xor2_1 \U$$1739  (.A(\t$5293 ),
    .B(net1474),
    .X(booth_b24_m44));
 sky130_fd_sc_hd__xor2_1 \U$$174  (.A(\t$4494 ),
    .B(net1386),
    .X(booth_b2_m15));
 sky130_fd_sc_hd__a22o_1 \U$$1740  (.A1(net1724),
    .A2(net609),
    .B1(net1715),
    .B2(net882),
    .X(\t$5294 ));
 sky130_fd_sc_hd__xor2_1 \U$$1741  (.A(\t$5294 ),
    .B(net1474),
    .X(booth_b24_m45));
 sky130_fd_sc_hd__a22o_1 \U$$1742  (.A1(net1715),
    .A2(net609),
    .B1(net1706),
    .B2(net882),
    .X(\t$5295 ));
 sky130_fd_sc_hd__xor2_1 \U$$1743  (.A(\t$5295 ),
    .B(net1474),
    .X(booth_b24_m46));
 sky130_fd_sc_hd__a22o_1 \U$$1744  (.A1(net1705),
    .A2(net607),
    .B1(net1695),
    .B2(net880),
    .X(\t$5296 ));
 sky130_fd_sc_hd__xor2_1 \U$$1745  (.A(\t$5296 ),
    .B(net1473),
    .X(booth_b24_m47));
 sky130_fd_sc_hd__a22o_1 \U$$1746  (.A1(net1697),
    .A2(net607),
    .B1(net1689),
    .B2(net880),
    .X(\t$5297 ));
 sky130_fd_sc_hd__xor2_1 \U$$1747  (.A(\t$5297 ),
    .B(net1473),
    .X(booth_b24_m48));
 sky130_fd_sc_hd__a22o_1 \U$$1748  (.A1(net1687),
    .A2(net607),
    .B1(net1679),
    .B2(net880),
    .X(\t$5298 ));
 sky130_fd_sc_hd__xor2_1 \U$$1749  (.A(\t$5298 ),
    .B(net1473),
    .X(booth_b24_m49));
 sky130_fd_sc_hd__a22o_1 \U$$175  (.A1(net1166),
    .A2(net620),
    .B1(net1157),
    .B2(net893),
    .X(\t$4495 ));
 sky130_fd_sc_hd__a22o_1 \U$$1750  (.A1(net1679),
    .A2(net607),
    .B1(net1654),
    .B2(net880),
    .X(\t$5299 ));
 sky130_fd_sc_hd__xor2_1 \U$$1751  (.A(\t$5299 ),
    .B(net1473),
    .X(booth_b24_m50));
 sky130_fd_sc_hd__a22o_1 \U$$1752  (.A1(net1654),
    .A2(net607),
    .B1(net1646),
    .B2(net880),
    .X(\t$5300 ));
 sky130_fd_sc_hd__xor2_1 \U$$1753  (.A(\t$5300 ),
    .B(net1473),
    .X(booth_b24_m51));
 sky130_fd_sc_hd__a22o_1 \U$$1754  (.A1(net1646),
    .A2(net607),
    .B1(net1638),
    .B2(net880),
    .X(\t$5301 ));
 sky130_fd_sc_hd__xor2_1 \U$$1755  (.A(\t$5301 ),
    .B(net1473),
    .X(booth_b24_m52));
 sky130_fd_sc_hd__a22o_1 \U$$1756  (.A1(net1639),
    .A2(net609),
    .B1(net1631),
    .B2(net882),
    .X(\t$5302 ));
 sky130_fd_sc_hd__xor2_1 \U$$1757  (.A(\t$5302 ),
    .B(net1474),
    .X(booth_b24_m53));
 sky130_fd_sc_hd__a22o_1 \U$$1758  (.A1(net1630),
    .A2(net607),
    .B1(net1621),
    .B2(net880),
    .X(\t$5303 ));
 sky130_fd_sc_hd__xor2_1 \U$$1759  (.A(\t$5303 ),
    .B(net1473),
    .X(booth_b24_m54));
 sky130_fd_sc_hd__xor2_1 \U$$176  (.A(\t$4495 ),
    .B(net1386),
    .X(booth_b2_m16));
 sky130_fd_sc_hd__a22o_1 \U$$1760  (.A1(net1622),
    .A2(net608),
    .B1(net1613),
    .B2(net881),
    .X(\t$5304 ));
 sky130_fd_sc_hd__xor2_1 \U$$1761  (.A(\t$5304 ),
    .B(net1471),
    .X(booth_b24_m55));
 sky130_fd_sc_hd__a22o_1 \U$$1762  (.A1(net1613),
    .A2(net608),
    .B1(net1605),
    .B2(net881),
    .X(\t$5305 ));
 sky130_fd_sc_hd__xor2_1 \U$$1763  (.A(\t$5305 ),
    .B(net1472),
    .X(booth_b24_m56));
 sky130_fd_sc_hd__a22o_1 \U$$1764  (.A1(net1605),
    .A2(net608),
    .B1(net1597),
    .B2(net881),
    .X(\t$5306 ));
 sky130_fd_sc_hd__xor2_1 \U$$1765  (.A(\t$5306 ),
    .B(net1472),
    .X(booth_b24_m57));
 sky130_fd_sc_hd__a22o_1 \U$$1766  (.A1(net1597),
    .A2(net607),
    .B1(net1588),
    .B2(net880),
    .X(\t$5307 ));
 sky130_fd_sc_hd__xor2_1 \U$$1767  (.A(\t$5307 ),
    .B(net1471),
    .X(booth_b24_m58));
 sky130_fd_sc_hd__a22o_1 \U$$1768  (.A1(net1588),
    .A2(net608),
    .B1(net1579),
    .B2(net881),
    .X(\t$5308 ));
 sky130_fd_sc_hd__xor2_1 \U$$1769  (.A(\t$5308 ),
    .B(net1471),
    .X(booth_b24_m59));
 sky130_fd_sc_hd__a22o_1 \U$$177  (.A1(net1157),
    .A2(net623),
    .B1(net1149),
    .B2(net896),
    .X(\t$4496 ));
 sky130_fd_sc_hd__a22o_1 \U$$1770  (.A1(net1579),
    .A2(net608),
    .B1(net1553),
    .B2(net881),
    .X(\t$5309 ));
 sky130_fd_sc_hd__xor2_1 \U$$1771  (.A(\t$5309 ),
    .B(net1471),
    .X(booth_b24_m60));
 sky130_fd_sc_hd__a22o_1 \U$$1772  (.A1(net1553),
    .A2(net607),
    .B1(net1544),
    .B2(net880),
    .X(\t$5310 ));
 sky130_fd_sc_hd__xor2_1 \U$$1773  (.A(\t$5310 ),
    .B(net1471),
    .X(booth_b24_m61));
 sky130_fd_sc_hd__a22o_1 \U$$1774  (.A1(net1544),
    .A2(net608),
    .B1(net1536),
    .B2(net881),
    .X(\t$5311 ));
 sky130_fd_sc_hd__xor2_1 \U$$1775  (.A(\t$5311 ),
    .B(net1471),
    .X(booth_b24_m62));
 sky130_fd_sc_hd__a22o_1 \U$$1776  (.A1(net1536),
    .A2(net608),
    .B1(net1528),
    .B2(net881),
    .X(\t$5312 ));
 sky130_fd_sc_hd__xor2_1 \U$$1777  (.A(\t$5312 ),
    .B(net1471),
    .X(booth_b24_m63));
 sky130_fd_sc_hd__a22o_1 \U$$1778  (.A1(net1529),
    .A2(net609),
    .B1(net1766),
    .B2(net882),
    .X(\t$5313 ));
 sky130_fd_sc_hd__xor2_1 \U$$1779  (.A(\t$5313 ),
    .B(net1474),
    .X(booth_b24_m64));
 sky130_fd_sc_hd__xor2_1 \U$$178  (.A(\t$4496 ),
    .B(net1389),
    .X(booth_b2_m17));
 sky130_fd_sc_hd__inv_1 \U$$1780  (.A(net1474),
    .Y(\notsign$5314 ));
 sky130_fd_sc_hd__inv_1 \U$$1781  (.A(net1471),
    .Y(\notblock$5315[0] ));
 sky130_fd_sc_hd__inv_1 \U$$1782  (.A(net19),
    .Y(\notblock$5315[1] ));
 sky130_fd_sc_hd__inv_1 \U$$1783  (.A(net1463),
    .Y(\notblock$5315[2] ));
 sky130_fd_sc_hd__and2_1 \U$$1784  (.A(net1463),
    .B(\notblock$5315[1] ),
    .X(\t$5316 ));
 sky130_fd_sc_hd__a32o_1 \U$$1785  (.A1(\notblock$5315[2] ),
    .A2(net19),
    .A3(net1472),
    .B1(\t$5316 ),
    .B2(\notblock$5315[0] ),
    .X(\sel_0$5317 ));
 sky130_fd_sc_hd__xor2_1 \U$$1786  (.A(net19),
    .B(net1472),
    .X(\sel_1$5318 ));
 sky130_fd_sc_hd__a22o_1 \U$$1787  (.A1(net1767),
    .A2(net594),
    .B1(net1228),
    .B2(net867),
    .X(\t$5319 ));
 sky130_fd_sc_hd__xor2_1 \U$$1788  (.A(\t$5319 ),
    .B(net1457),
    .X(booth_b26_m0));
 sky130_fd_sc_hd__a22o_1 \U$$1789  (.A1(net1227),
    .A2(net593),
    .B1(net1122),
    .B2(net866),
    .X(\t$5320 ));
 sky130_fd_sc_hd__a22o_1 \U$$179  (.A1(net1149),
    .A2(net623),
    .B1(net1143),
    .B2(net896),
    .X(\t$4497 ));
 sky130_fd_sc_hd__xor2_1 \U$$1790  (.A(\t$5320 ),
    .B(net1457),
    .X(booth_b26_m1));
 sky130_fd_sc_hd__a22o_1 \U$$1791  (.A1(net1122),
    .A2(net593),
    .B1(net1031),
    .B2(net866),
    .X(\t$5321 ));
 sky130_fd_sc_hd__xor2_1 \U$$1792  (.A(\t$5321 ),
    .B(net1457),
    .X(booth_b26_m2));
 sky130_fd_sc_hd__a22o_1 \U$$1793  (.A1(net1031),
    .A2(net593),
    .B1(net932),
    .B2(net866),
    .X(\t$5322 ));
 sky130_fd_sc_hd__xor2_1 \U$$1794  (.A(\t$5322 ),
    .B(net1457),
    .X(booth_b26_m3));
 sky130_fd_sc_hd__a22o_1 \U$$1795  (.A1(net932),
    .A2(net593),
    .B1(net1671),
    .B2(net866),
    .X(\t$5323 ));
 sky130_fd_sc_hd__xor2_1 \U$$1796  (.A(\t$5323 ),
    .B(net1457),
    .X(booth_b26_m4));
 sky130_fd_sc_hd__a22o_1 \U$$1797  (.A1(net1671),
    .A2(net593),
    .B1(net1560),
    .B2(net866),
    .X(\t$5324 ));
 sky130_fd_sc_hd__xor2_1 \U$$1798  (.A(\t$5324 ),
    .B(net1457),
    .X(booth_b26_m5));
 sky130_fd_sc_hd__a22o_1 \U$$1799  (.A1(net1564),
    .A2(net596),
    .B1(net1524),
    .B2(net869),
    .X(\t$5325 ));
 sky130_fd_sc_hd__a22o_1 \U$$18  (.A1(net1565),
    .A2(net447),
    .B1(net1524),
    .B2(net689),
    .X(\t$4416 ));
 sky130_fd_sc_hd__xor2_1 \U$$180  (.A(\t$4497 ),
    .B(net1389),
    .X(booth_b2_m18));
 sky130_fd_sc_hd__xor2_1 \U$$1800  (.A(\t$5325 ),
    .B(net1460),
    .X(booth_b26_m6));
 sky130_fd_sc_hd__a22o_1 \U$$1801  (.A1(net1524),
    .A2(net597),
    .B1(net1516),
    .B2(net870),
    .X(\t$5326 ));
 sky130_fd_sc_hd__xor2_1 \U$$1802  (.A(\t$5326 ),
    .B(net1460),
    .X(booth_b26_m7));
 sky130_fd_sc_hd__a22o_1 \U$$1803  (.A1(net1516),
    .A2(net596),
    .B1(net1509),
    .B2(net869),
    .X(\t$5327 ));
 sky130_fd_sc_hd__xor2_1 \U$$1804  (.A(\t$5327 ),
    .B(net1460),
    .X(booth_b26_m8));
 sky130_fd_sc_hd__a22o_1 \U$$1805  (.A1(net1509),
    .A2(net597),
    .B1(net1500),
    .B2(net870),
    .X(\t$5328 ));
 sky130_fd_sc_hd__xor2_1 \U$$1806  (.A(\t$5328 ),
    .B(net1460),
    .X(booth_b26_m9));
 sky130_fd_sc_hd__a22o_1 \U$$1807  (.A1(net1499),
    .A2(net596),
    .B1(net1224),
    .B2(net869),
    .X(\t$5329 ));
 sky130_fd_sc_hd__xor2_1 \U$$1808  (.A(\t$5329 ),
    .B(net1460),
    .X(booth_b26_m10));
 sky130_fd_sc_hd__a22o_1 \U$$1809  (.A1(net1224),
    .A2(net596),
    .B1(net1216),
    .B2(net869),
    .X(\t$5330 ));
 sky130_fd_sc_hd__a22o_1 \U$$181  (.A1(net1143),
    .A2(net623),
    .B1(net1133),
    .B2(net896),
    .X(\t$4498 ));
 sky130_fd_sc_hd__xor2_1 \U$$1810  (.A(\t$5330 ),
    .B(net1460),
    .X(booth_b26_m11));
 sky130_fd_sc_hd__a22o_1 \U$$1811  (.A1(net1211),
    .A2(net596),
    .B1(net1203),
    .B2(net869),
    .X(\t$5331 ));
 sky130_fd_sc_hd__xor2_1 \U$$1812  (.A(\t$5331 ),
    .B(net1460),
    .X(booth_b26_m12));
 sky130_fd_sc_hd__a22o_1 \U$$1813  (.A1(net1203),
    .A2(net594),
    .B1(net1194),
    .B2(net867),
    .X(\t$5332 ));
 sky130_fd_sc_hd__xor2_1 \U$$1814  (.A(\t$5332 ),
    .B(net1457),
    .X(booth_b26_m13));
 sky130_fd_sc_hd__a22o_1 \U$$1815  (.A1(net1192),
    .A2(net594),
    .B1(net1173),
    .B2(net867),
    .X(\t$5333 ));
 sky130_fd_sc_hd__xor2_1 \U$$1816  (.A(\t$5333 ),
    .B(net1458),
    .X(booth_b26_m14));
 sky130_fd_sc_hd__a22o_1 \U$$1817  (.A1(net1173),
    .A2(net593),
    .B1(net1164),
    .B2(net866),
    .X(\t$5334 ));
 sky130_fd_sc_hd__xor2_1 \U$$1818  (.A(\t$5334 ),
    .B(net1457),
    .X(booth_b26_m15));
 sky130_fd_sc_hd__a22o_1 \U$$1819  (.A1(net1165),
    .A2(net593),
    .B1(net1155),
    .B2(net866),
    .X(\t$5335 ));
 sky130_fd_sc_hd__xor2_1 \U$$182  (.A(\t$4498 ),
    .B(net1389),
    .X(booth_b2_m19));
 sky130_fd_sc_hd__xor2_1 \U$$1820  (.A(\t$5335 ),
    .B(net1457),
    .X(booth_b26_m16));
 sky130_fd_sc_hd__a22o_1 \U$$1821  (.A1(net1156),
    .A2(net593),
    .B1(net1147),
    .B2(net866),
    .X(\t$5336 ));
 sky130_fd_sc_hd__xor2_1 \U$$1822  (.A(\t$5336 ),
    .B(net1457),
    .X(booth_b26_m17));
 sky130_fd_sc_hd__a22o_1 \U$$1823  (.A1(net1147),
    .A2(net594),
    .B1(net1139),
    .B2(net867),
    .X(\t$5337 ));
 sky130_fd_sc_hd__xor2_1 \U$$1824  (.A(\t$5337 ),
    .B(net1458),
    .X(booth_b26_m18));
 sky130_fd_sc_hd__a22o_1 \U$$1825  (.A1(net1139),
    .A2(net593),
    .B1(net1132),
    .B2(net866),
    .X(\t$5338 ));
 sky130_fd_sc_hd__xor2_1 \U$$1826  (.A(\t$5338 ),
    .B(net1458),
    .X(booth_b26_m19));
 sky130_fd_sc_hd__a22o_1 \U$$1827  (.A1(net1132),
    .A2(net594),
    .B1(net1116),
    .B2(net867),
    .X(\t$5339 ));
 sky130_fd_sc_hd__xor2_1 \U$$1828  (.A(\t$5339 ),
    .B(net1458),
    .X(booth_b26_m20));
 sky130_fd_sc_hd__a22o_1 \U$$1829  (.A1(net1116),
    .A2(net595),
    .B1(net1107),
    .B2(net868),
    .X(\t$5340 ));
 sky130_fd_sc_hd__a22o_1 \U$$183  (.A1(net1133),
    .A2(net623),
    .B1(net1117),
    .B2(net896),
    .X(\t$4499 ));
 sky130_fd_sc_hd__xor2_1 \U$$1830  (.A(\t$5340 ),
    .B(net1459),
    .X(booth_b26_m21));
 sky130_fd_sc_hd__a22o_1 \U$$1831  (.A1(net1107),
    .A2(net595),
    .B1(net1098),
    .B2(net868),
    .X(\t$5341 ));
 sky130_fd_sc_hd__xor2_1 \U$$1832  (.A(\t$5341 ),
    .B(net1459),
    .X(booth_b26_m22));
 sky130_fd_sc_hd__a22o_1 \U$$1833  (.A1(net1098),
    .A2(net593),
    .B1(net1090),
    .B2(net866),
    .X(\t$5342 ));
 sky130_fd_sc_hd__xor2_1 \U$$1834  (.A(\t$5342 ),
    .B(net1458),
    .X(booth_b26_m23));
 sky130_fd_sc_hd__a22o_1 \U$$1835  (.A1(net1090),
    .A2(net596),
    .B1(net1084),
    .B2(net869),
    .X(\t$5343 ));
 sky130_fd_sc_hd__xor2_1 \U$$1836  (.A(\t$5343 ),
    .B(net1460),
    .X(booth_b26_m24));
 sky130_fd_sc_hd__a22o_1 \U$$1837  (.A1(net1083),
    .A2(net596),
    .B1(net1074),
    .B2(net869),
    .X(\t$5344 ));
 sky130_fd_sc_hd__xor2_1 \U$$1838  (.A(\t$5344 ),
    .B(net1461),
    .X(booth_b26_m25));
 sky130_fd_sc_hd__a22o_1 \U$$1839  (.A1(net1074),
    .A2(net596),
    .B1(net1066),
    .B2(net869),
    .X(\t$5345 ));
 sky130_fd_sc_hd__xor2_1 \U$$184  (.A(\t$4499 ),
    .B(net1389),
    .X(booth_b2_m20));
 sky130_fd_sc_hd__xor2_1 \U$$1840  (.A(\t$5345 ),
    .B(net1461),
    .X(booth_b26_m26));
 sky130_fd_sc_hd__a22o_1 \U$$1841  (.A1(net1066),
    .A2(net596),
    .B1(net1057),
    .B2(net869),
    .X(\t$5346 ));
 sky130_fd_sc_hd__xor2_1 \U$$1842  (.A(\t$5346 ),
    .B(net1461),
    .X(booth_b26_m27));
 sky130_fd_sc_hd__a22o_1 \U$$1843  (.A1(net1057),
    .A2(net597),
    .B1(net1049),
    .B2(net870),
    .X(\t$5347 ));
 sky130_fd_sc_hd__xor2_1 \U$$1844  (.A(\t$5347 ),
    .B(net1461),
    .X(booth_b26_m28));
 sky130_fd_sc_hd__a22o_1 \U$$1845  (.A1(net1049),
    .A2(net597),
    .B1(net1042),
    .B2(net870),
    .X(\t$5348 ));
 sky130_fd_sc_hd__xor2_1 \U$$1846  (.A(\t$5348 ),
    .B(net1461),
    .X(booth_b26_m29));
 sky130_fd_sc_hd__a22o_1 \U$$1847  (.A1(net1041),
    .A2(net601),
    .B1(net1025),
    .B2(net874),
    .X(\t$5349 ));
 sky130_fd_sc_hd__xor2_1 \U$$1848  (.A(\t$5349 ),
    .B(net1460),
    .X(booth_b26_m30));
 sky130_fd_sc_hd__a22o_1 \U$$1849  (.A1(net1025),
    .A2(net596),
    .B1(net1017),
    .B2(net869),
    .X(\t$5350 ));
 sky130_fd_sc_hd__a22o_1 \U$$185  (.A1(net1117),
    .A2(net623),
    .B1(net1108),
    .B2(net896),
    .X(\t$4500 ));
 sky130_fd_sc_hd__xor2_1 \U$$1850  (.A(\t$5350 ),
    .B(net1460),
    .X(booth_b26_m31));
 sky130_fd_sc_hd__a22o_1 \U$$1851  (.A1(net1018),
    .A2(net597),
    .B1(net1001),
    .B2(net870),
    .X(\t$5351 ));
 sky130_fd_sc_hd__xor2_1 \U$$1852  (.A(\t$5351 ),
    .B(net1462),
    .X(booth_b26_m32));
 sky130_fd_sc_hd__a22o_1 \U$$1853  (.A1(net999),
    .A2(net597),
    .B1(net991),
    .B2(net870),
    .X(\t$5352 ));
 sky130_fd_sc_hd__xor2_1 \U$$1854  (.A(\t$5352 ),
    .B(net1462),
    .X(booth_b26_m33));
 sky130_fd_sc_hd__a22o_1 \U$$1855  (.A1(net991),
    .A2(net597),
    .B1(net983),
    .B2(net870),
    .X(\t$5353 ));
 sky130_fd_sc_hd__xor2_1 \U$$1856  (.A(\t$5353 ),
    .B(net1462),
    .X(booth_b26_m34));
 sky130_fd_sc_hd__a22o_1 \U$$1857  (.A1(net982),
    .A2(net595),
    .B1(net973),
    .B2(net868),
    .X(\t$5354 ));
 sky130_fd_sc_hd__xor2_1 \U$$1858  (.A(\t$5354 ),
    .B(net1459),
    .X(booth_b26_m35));
 sky130_fd_sc_hd__a22o_1 \U$$1859  (.A1(net974),
    .A2(net595),
    .B1(net965),
    .B2(net868),
    .X(\t$5355 ));
 sky130_fd_sc_hd__xor2_1 \U$$186  (.A(\t$4500 ),
    .B(net1389),
    .X(booth_b2_m21));
 sky130_fd_sc_hd__xor2_1 \U$$1860  (.A(\t$5355 ),
    .B(net1459),
    .X(booth_b26_m36));
 sky130_fd_sc_hd__a22o_1 \U$$1861  (.A1(net965),
    .A2(net598),
    .B1(net957),
    .B2(net871),
    .X(\t$5356 ));
 sky130_fd_sc_hd__xor2_1 \U$$1862  (.A(\t$5356 ),
    .B(net1459),
    .X(booth_b26_m37));
 sky130_fd_sc_hd__a22o_1 \U$$1863  (.A1(net961),
    .A2(net597),
    .B1(net955),
    .B2(net870),
    .X(\t$5357 ));
 sky130_fd_sc_hd__xor2_1 \U$$1864  (.A(\t$5357 ),
    .B(net1462),
    .X(booth_b26_m38));
 sky130_fd_sc_hd__a22o_1 \U$$1865  (.A1(net955),
    .A2(net601),
    .B1(net944),
    .B2(net874),
    .X(\t$5358 ));
 sky130_fd_sc_hd__xor2_1 \U$$1866  (.A(\t$5358 ),
    .B(net1462),
    .X(booth_b26_m39));
 sky130_fd_sc_hd__a22o_1 \U$$1867  (.A1(net944),
    .A2(net597),
    .B1(net928),
    .B2(net870),
    .X(\t$5359 ));
 sky130_fd_sc_hd__xor2_1 \U$$1868  (.A(\t$5359 ),
    .B(net1462),
    .X(booth_b26_m40));
 sky130_fd_sc_hd__a22o_1 \U$$1869  (.A1(net930),
    .A2(net600),
    .B1(net1751),
    .B2(net873),
    .X(\t$5360 ));
 sky130_fd_sc_hd__a22o_1 \U$$187  (.A1(net1106),
    .A2(net620),
    .B1(net1099),
    .B2(net893),
    .X(\t$4501 ));
 sky130_fd_sc_hd__xor2_1 \U$$1870  (.A(\t$5360 ),
    .B(net1465),
    .X(booth_b26_m41));
 sky130_fd_sc_hd__a22o_1 \U$$1871  (.A1(net1747),
    .A2(net600),
    .B1(net1739),
    .B2(net873),
    .X(\t$5361 ));
 sky130_fd_sc_hd__xor2_1 \U$$1872  (.A(\t$5361 ),
    .B(net1465),
    .X(booth_b26_m42));
 sky130_fd_sc_hd__a22o_1 \U$$1873  (.A1(net1741),
    .A2(net600),
    .B1(net1733),
    .B2(net873),
    .X(\t$5362 ));
 sky130_fd_sc_hd__xor2_1 \U$$1874  (.A(\t$5362 ),
    .B(net1465),
    .X(booth_b26_m43));
 sky130_fd_sc_hd__a22o_1 \U$$1875  (.A1(net1733),
    .A2(net600),
    .B1(net1724),
    .B2(net873),
    .X(\t$5363 ));
 sky130_fd_sc_hd__xor2_1 \U$$1876  (.A(\t$5363 ),
    .B(net1465),
    .X(booth_b26_m44));
 sky130_fd_sc_hd__a22o_1 \U$$1877  (.A1(net1721),
    .A2(net598),
    .B1(net1712),
    .B2(net871),
    .X(\t$5364 ));
 sky130_fd_sc_hd__xor2_1 \U$$1878  (.A(\t$5364 ),
    .B(net1464),
    .X(booth_b26_m45));
 sky130_fd_sc_hd__a22o_1 \U$$1879  (.A1(net1712),
    .A2(net598),
    .B1(net1705),
    .B2(net871),
    .X(\t$5365 ));
 sky130_fd_sc_hd__xor2_1 \U$$188  (.A(\t$4501 ),
    .B(net1386),
    .X(booth_b2_m22));
 sky130_fd_sc_hd__xor2_1 \U$$1880  (.A(\t$5365 ),
    .B(net1464),
    .X(booth_b26_m46));
 sky130_fd_sc_hd__a22o_1 \U$$1881  (.A1(net1703),
    .A2(net598),
    .B1(net1695),
    .B2(net871),
    .X(\t$5366 ));
 sky130_fd_sc_hd__xor2_1 \U$$1882  (.A(\t$5366 ),
    .B(net1464),
    .X(booth_b26_m47));
 sky130_fd_sc_hd__a22o_1 \U$$1883  (.A1(net1695),
    .A2(net598),
    .B1(net1687),
    .B2(net871),
    .X(\t$5367 ));
 sky130_fd_sc_hd__xor2_1 \U$$1884  (.A(\t$5367 ),
    .B(net1459),
    .X(booth_b26_m48));
 sky130_fd_sc_hd__a22o_1 \U$$1885  (.A1(net1687),
    .A2(net598),
    .B1(net1679),
    .B2(net871),
    .X(\t$5368 ));
 sky130_fd_sc_hd__xor2_1 \U$$1886  (.A(\t$5368 ),
    .B(net1464),
    .X(booth_b26_m49));
 sky130_fd_sc_hd__a22o_1 \U$$1887  (.A1(net1679),
    .A2(net598),
    .B1(net1654),
    .B2(net871),
    .X(\t$5369 ));
 sky130_fd_sc_hd__xor2_1 \U$$1888  (.A(\t$5369 ),
    .B(net1464),
    .X(booth_b26_m50));
 sky130_fd_sc_hd__a22o_1 \U$$1889  (.A1(net1659),
    .A2(net600),
    .B1(net1647),
    .B2(net873),
    .X(\t$5370 ));
 sky130_fd_sc_hd__a22o_1 \U$$189  (.A1(net1097),
    .A2(net620),
    .B1(net1088),
    .B2(net893),
    .X(\t$4502 ));
 sky130_fd_sc_hd__xor2_1 \U$$1890  (.A(\t$5370 ),
    .B(net1465),
    .X(booth_b26_m51));
 sky130_fd_sc_hd__a22o_1 \U$$1891  (.A1(net1647),
    .A2(net598),
    .B1(net1638),
    .B2(net871),
    .X(\t$5371 ));
 sky130_fd_sc_hd__xor2_1 \U$$1892  (.A(\t$5371 ),
    .B(net1464),
    .X(booth_b26_m52));
 sky130_fd_sc_hd__a22o_1 \U$$1893  (.A1(net1639),
    .A2(net598),
    .B1(net1631),
    .B2(net871),
    .X(\t$5372 ));
 sky130_fd_sc_hd__xor2_1 \U$$1894  (.A(\t$5372 ),
    .B(net1464),
    .X(booth_b26_m53));
 sky130_fd_sc_hd__a22o_1 \U$$1895  (.A1(net1631),
    .A2(net598),
    .B1(net1622),
    .B2(net871),
    .X(\t$5373 ));
 sky130_fd_sc_hd__xor2_1 \U$$1896  (.A(\t$5373 ),
    .B(net1463),
    .X(booth_b26_m54));
 sky130_fd_sc_hd__a22o_1 \U$$1897  (.A1(net1622),
    .A2(net599),
    .B1(net1613),
    .B2(net872),
    .X(\t$5374 ));
 sky130_fd_sc_hd__xor2_1 \U$$1898  (.A(\t$5374 ),
    .B(net1464),
    .X(booth_b26_m55));
 sky130_fd_sc_hd__a22o_1 \U$$1899  (.A1(net1613),
    .A2(net599),
    .B1(net1605),
    .B2(net872),
    .X(\t$5375 ));
 sky130_fd_sc_hd__xor2_1 \U$$19  (.A(\t$4416 ),
    .B(net1574),
    .X(booth_b0_m6));
 sky130_fd_sc_hd__xor2_1 \U$$190  (.A(\t$4502 ),
    .B(net1386),
    .X(booth_b2_m23));
 sky130_fd_sc_hd__xor2_1 \U$$1900  (.A(\t$5375 ),
    .B(net1463),
    .X(booth_b26_m56));
 sky130_fd_sc_hd__a22o_1 \U$$1901  (.A1(net1605),
    .A2(net599),
    .B1(net1597),
    .B2(net872),
    .X(\t$5376 ));
 sky130_fd_sc_hd__xor2_1 \U$$1902  (.A(\t$5376 ),
    .B(net1464),
    .X(booth_b26_m57));
 sky130_fd_sc_hd__a22o_1 \U$$1903  (.A1(net1597),
    .A2(net599),
    .B1(net1588),
    .B2(net872),
    .X(\t$5377 ));
 sky130_fd_sc_hd__xor2_1 \U$$1904  (.A(\t$5377 ),
    .B(net1463),
    .X(booth_b26_m58));
 sky130_fd_sc_hd__a22o_1 \U$$1905  (.A1(net1588),
    .A2(net599),
    .B1(net1579),
    .B2(net872),
    .X(\t$5378 ));
 sky130_fd_sc_hd__xor2_1 \U$$1906  (.A(\t$5378 ),
    .B(net1463),
    .X(booth_b26_m59));
 sky130_fd_sc_hd__a22o_1 \U$$1907  (.A1(net1579),
    .A2(net599),
    .B1(net1553),
    .B2(net872),
    .X(\t$5379 ));
 sky130_fd_sc_hd__xor2_1 \U$$1908  (.A(\t$5379 ),
    .B(net1463),
    .X(booth_b26_m60));
 sky130_fd_sc_hd__a22o_1 \U$$1909  (.A1(net1553),
    .A2(net599),
    .B1(net1544),
    .B2(net872),
    .X(\t$5380 ));
 sky130_fd_sc_hd__a22o_1 \U$$191  (.A1(net1088),
    .A2(net619),
    .B1(net1080),
    .B2(net892),
    .X(\t$4503 ));
 sky130_fd_sc_hd__xor2_1 \U$$1910  (.A(\t$5380 ),
    .B(net1463),
    .X(booth_b26_m61));
 sky130_fd_sc_hd__a22o_1 \U$$1911  (.A1(net1545),
    .A2(net600),
    .B1(net1537),
    .B2(net873),
    .X(\t$5381 ));
 sky130_fd_sc_hd__xor2_1 \U$$1912  (.A(\t$5381 ),
    .B(net1465),
    .X(booth_b26_m62));
 sky130_fd_sc_hd__a22o_1 \U$$1913  (.A1(net1540),
    .A2(net600),
    .B1(net1532),
    .B2(net873),
    .X(\t$5382 ));
 sky130_fd_sc_hd__xor2_1 \U$$1914  (.A(\t$5382 ),
    .B(net1465),
    .X(booth_b26_m63));
 sky130_fd_sc_hd__a22o_1 \U$$1915  (.A1(net1532),
    .A2(net600),
    .B1(net1768),
    .B2(net873),
    .X(\t$5383 ));
 sky130_fd_sc_hd__xor2_1 \U$$1916  (.A(\t$5383 ),
    .B(net1465),
    .X(booth_b26_m64));
 sky130_fd_sc_hd__inv_1 \U$$1917  (.A(net20),
    .Y(\notsign$5384 ));
 sky130_fd_sc_hd__inv_1 \U$$1918  (.A(net1463),
    .Y(\notblock$5385[0] ));
 sky130_fd_sc_hd__inv_1 \U$$1919  (.A(net21),
    .Y(\notblock$5385[1] ));
 sky130_fd_sc_hd__xor2_1 \U$$192  (.A(\t$4503 ),
    .B(net1385),
    .X(booth_b2_m24));
 sky130_fd_sc_hd__inv_1 \U$$1920  (.A(net1453),
    .Y(\notblock$5385[2] ));
 sky130_fd_sc_hd__and2_1 \U$$1921  (.A(net1453),
    .B(\notblock$5385[1] ),
    .X(\t$5386 ));
 sky130_fd_sc_hd__a32o_1 \U$$1922  (.A1(\notblock$5385[2] ),
    .A2(net21),
    .A3(net1463),
    .B1(\t$5386 ),
    .B2(\notblock$5385[0] ),
    .X(\sel_0$5387 ));
 sky130_fd_sc_hd__xor2_2 \U$$1923  (.A(net21),
    .B(net1464),
    .X(\sel_1$5388 ));
 sky130_fd_sc_hd__a22o_1 \U$$1924  (.A1(net1769),
    .A2(net584),
    .B1(net1227),
    .B2(net857),
    .X(\t$5389 ));
 sky130_fd_sc_hd__xor2_1 \U$$1925  (.A(\t$5389 ),
    .B(net1448),
    .X(booth_b28_m0));
 sky130_fd_sc_hd__a22o_1 \U$$1926  (.A1(net1227),
    .A2(net584),
    .B1(net1122),
    .B2(net857),
    .X(\t$5390 ));
 sky130_fd_sc_hd__xor2_1 \U$$1927  (.A(\t$5390 ),
    .B(net1448),
    .X(booth_b28_m1));
 sky130_fd_sc_hd__a22o_1 \U$$1928  (.A1(net1122),
    .A2(net584),
    .B1(net1031),
    .B2(net857),
    .X(\t$5391 ));
 sky130_fd_sc_hd__xor2_1 \U$$1929  (.A(\t$5391 ),
    .B(net1448),
    .X(booth_b28_m2));
 sky130_fd_sc_hd__a22o_1 \U$$193  (.A1(net1080),
    .A2(net619),
    .B1(net1071),
    .B2(net892),
    .X(\t$4504 ));
 sky130_fd_sc_hd__a22o_1 \U$$1930  (.A1(net1031),
    .A2(net584),
    .B1(net932),
    .B2(net857),
    .X(\t$5392 ));
 sky130_fd_sc_hd__xor2_1 \U$$1931  (.A(\t$5392 ),
    .B(net1448),
    .X(booth_b28_m3));
 sky130_fd_sc_hd__a22o_1 \U$$1932  (.A1(net936),
    .A2(net587),
    .B1(net1676),
    .B2(net860),
    .X(\t$5393 ));
 sky130_fd_sc_hd__xor2_1 \U$$1933  (.A(\t$5393 ),
    .B(net1451),
    .X(booth_b28_m4));
 sky130_fd_sc_hd__a22o_1 \U$$1934  (.A1(net1675),
    .A2(net588),
    .B1(net1565),
    .B2(net861),
    .X(\t$5394 ));
 sky130_fd_sc_hd__xor2_1 \U$$1935  (.A(\t$5394 ),
    .B(net1451),
    .X(booth_b28_m5));
 sky130_fd_sc_hd__a22o_1 \U$$1936  (.A1(net1565),
    .A2(net587),
    .B1(net1524),
    .B2(net860),
    .X(\t$5395 ));
 sky130_fd_sc_hd__xor2_1 \U$$1937  (.A(\t$5395 ),
    .B(net1451),
    .X(booth_b28_m6));
 sky130_fd_sc_hd__a22o_1 \U$$1938  (.A1(net1524),
    .A2(net587),
    .B1(net1516),
    .B2(net860),
    .X(\t$5396 ));
 sky130_fd_sc_hd__xor2_1 \U$$1939  (.A(\t$5396 ),
    .B(net1451),
    .X(booth_b28_m7));
 sky130_fd_sc_hd__xor2_1 \U$$194  (.A(\t$4504 ),
    .B(net1385),
    .X(booth_b2_m25));
 sky130_fd_sc_hd__a22o_1 \U$$1940  (.A1(net1516),
    .A2(net588),
    .B1(net1508),
    .B2(net861),
    .X(\t$5397 ));
 sky130_fd_sc_hd__xor2_1 \U$$1941  (.A(\t$5397 ),
    .B(net1451),
    .X(booth_b28_m8));
 sky130_fd_sc_hd__a22o_1 \U$$1942  (.A1(net1508),
    .A2(net587),
    .B1(net1499),
    .B2(net860),
    .X(\t$5398 ));
 sky130_fd_sc_hd__xor2_1 \U$$1943  (.A(\t$5398 ),
    .B(net1451),
    .X(booth_b28_m9));
 sky130_fd_sc_hd__a22o_1 \U$$1944  (.A1(net1494),
    .A2(net584),
    .B1(net1219),
    .B2(net857),
    .X(\t$5399 ));
 sky130_fd_sc_hd__xor2_1 \U$$1945  (.A(\t$5399 ),
    .B(net1448),
    .X(booth_b28_m10));
 sky130_fd_sc_hd__a22o_1 \U$$1946  (.A1(net1221),
    .A2(net585),
    .B1(net1211),
    .B2(net858),
    .X(\t$5400 ));
 sky130_fd_sc_hd__xor2_1 \U$$1947  (.A(\t$5400 ),
    .B(net1449),
    .X(booth_b28_m11));
 sky130_fd_sc_hd__a22o_1 \U$$1948  (.A1(net1211),
    .A2(net585),
    .B1(net1201),
    .B2(net858),
    .X(\t$5401 ));
 sky130_fd_sc_hd__xor2_1 \U$$1949  (.A(\t$5401 ),
    .B(net1449),
    .X(booth_b28_m12));
 sky130_fd_sc_hd__a22o_1 \U$$195  (.A1(net1071),
    .A2(net619),
    .B1(net1063),
    .B2(net892),
    .X(\t$4505 ));
 sky130_fd_sc_hd__a22o_1 \U$$1950  (.A1(net1201),
    .A2(net584),
    .B1(net1192),
    .B2(net857),
    .X(\t$5402 ));
 sky130_fd_sc_hd__xor2_1 \U$$1951  (.A(\t$5402 ),
    .B(net1448),
    .X(booth_b28_m13));
 sky130_fd_sc_hd__a22o_1 \U$$1952  (.A1(net1192),
    .A2(net584),
    .B1(net1173),
    .B2(net857),
    .X(\t$5403 ));
 sky130_fd_sc_hd__xor2_1 \U$$1953  (.A(\t$5403 ),
    .B(net1448),
    .X(booth_b28_m14));
 sky130_fd_sc_hd__a22o_1 \U$$1954  (.A1(net1173),
    .A2(net584),
    .B1(net1164),
    .B2(net857),
    .X(\t$5404 ));
 sky130_fd_sc_hd__xor2_1 \U$$1955  (.A(\t$5404 ),
    .B(net1448),
    .X(booth_b28_m15));
 sky130_fd_sc_hd__a22o_1 \U$$1956  (.A1(net1166),
    .A2(net585),
    .B1(net1157),
    .B2(net858),
    .X(\t$5405 ));
 sky130_fd_sc_hd__xor2_1 \U$$1957  (.A(\t$5405 ),
    .B(net1449),
    .X(booth_b28_m16));
 sky130_fd_sc_hd__a22o_1 \U$$1958  (.A1(net1158),
    .A2(net585),
    .B1(net1147),
    .B2(net858),
    .X(\t$5406 ));
 sky130_fd_sc_hd__xor2_1 \U$$1959  (.A(\t$5406 ),
    .B(net1449),
    .X(booth_b28_m17));
 sky130_fd_sc_hd__xor2_1 \U$$196  (.A(\t$4505 ),
    .B(net1385),
    .X(booth_b2_m26));
 sky130_fd_sc_hd__a22o_1 \U$$1960  (.A1(net1148),
    .A2(net585),
    .B1(net1138),
    .B2(net858),
    .X(\t$5407 ));
 sky130_fd_sc_hd__xor2_1 \U$$1961  (.A(\t$5407 ),
    .B(net1449),
    .X(booth_b28_m18));
 sky130_fd_sc_hd__a22o_1 \U$$1962  (.A1(net1140),
    .A2(net586),
    .B1(net1132),
    .B2(net859),
    .X(\t$5408 ));
 sky130_fd_sc_hd__xor2_1 \U$$1963  (.A(\t$5408 ),
    .B(net1450),
    .X(booth_b28_m19));
 sky130_fd_sc_hd__a22o_1 \U$$1964  (.A1(net1132),
    .A2(net584),
    .B1(net1116),
    .B2(net857),
    .X(\t$5409 ));
 sky130_fd_sc_hd__xor2_1 \U$$1965  (.A(\t$5409 ),
    .B(net1448),
    .X(booth_b28_m20));
 sky130_fd_sc_hd__a22o_1 \U$$1966  (.A1(net1116),
    .A2(net584),
    .B1(net1107),
    .B2(net857),
    .X(\t$5410 ));
 sky130_fd_sc_hd__xor2_1 \U$$1967  (.A(\t$5410 ),
    .B(net1449),
    .X(booth_b28_m21));
 sky130_fd_sc_hd__a22o_1 \U$$1968  (.A1(net1107),
    .A2(net585),
    .B1(net1098),
    .B2(net858),
    .X(\t$5411 ));
 sky130_fd_sc_hd__xor2_1 \U$$1969  (.A(\t$5411 ),
    .B(net1449),
    .X(booth_b28_m22));
 sky130_fd_sc_hd__a22o_1 \U$$197  (.A1(net1063),
    .A2(net619),
    .B1(net1055),
    .B2(net892),
    .X(\t$4506 ));
 sky130_fd_sc_hd__a22o_1 \U$$1970  (.A1(net1101),
    .A2(net587),
    .B1(net1091),
    .B2(net860),
    .X(\t$5412 ));
 sky130_fd_sc_hd__xor2_1 \U$$1971  (.A(\t$5412 ),
    .B(net1451),
    .X(booth_b28_m23));
 sky130_fd_sc_hd__a22o_1 \U$$1972  (.A1(net1091),
    .A2(net587),
    .B1(net1083),
    .B2(net860),
    .X(\t$5413 ));
 sky130_fd_sc_hd__xor2_1 \U$$1973  (.A(\t$5413 ),
    .B(net1451),
    .X(booth_b28_m24));
 sky130_fd_sc_hd__a22o_1 \U$$1974  (.A1(net1083),
    .A2(net587),
    .B1(net1074),
    .B2(net860),
    .X(\t$5414 ));
 sky130_fd_sc_hd__xor2_1 \U$$1975  (.A(\t$5414 ),
    .B(net1451),
    .X(booth_b28_m25));
 sky130_fd_sc_hd__a22o_1 \U$$1976  (.A1(net1074),
    .A2(net587),
    .B1(net1066),
    .B2(net860),
    .X(\t$5415 ));
 sky130_fd_sc_hd__xor2_1 \U$$1977  (.A(\t$5415 ),
    .B(net1452),
    .X(booth_b28_m26));
 sky130_fd_sc_hd__a22o_1 \U$$1978  (.A1(net1067),
    .A2(net587),
    .B1(net1057),
    .B2(net860),
    .X(\t$5416 ));
 sky130_fd_sc_hd__xor2_1 \U$$1979  (.A(\t$5416 ),
    .B(net1452),
    .X(booth_b28_m27));
 sky130_fd_sc_hd__xor2_1 \U$$198  (.A(\t$4506 ),
    .B(net1385),
    .X(booth_b2_m27));
 sky130_fd_sc_hd__a22o_1 \U$$1980  (.A1(net1058),
    .A2(net588),
    .B1(net1050),
    .B2(net861),
    .X(\t$5417 ));
 sky130_fd_sc_hd__xor2_1 \U$$1981  (.A(\t$5417 ),
    .B(net1452),
    .X(booth_b28_m28));
 sky130_fd_sc_hd__a22o_1 \U$$1982  (.A1(net1049),
    .A2(net587),
    .B1(net1041),
    .B2(net860),
    .X(\t$5418 ));
 sky130_fd_sc_hd__xor2_1 \U$$1983  (.A(\t$5418 ),
    .B(net1451),
    .X(booth_b28_m29));
 sky130_fd_sc_hd__a22o_1 \U$$1984  (.A1(net1042),
    .A2(net588),
    .B1(net1026),
    .B2(net861),
    .X(\t$5419 ));
 sky130_fd_sc_hd__xor2_1 \U$$1985  (.A(\t$5419 ),
    .B(net1452),
    .X(booth_b28_m30));
 sky130_fd_sc_hd__a22o_1 \U$$1986  (.A1(net1026),
    .A2(net588),
    .B1(net1018),
    .B2(net861),
    .X(\t$5420 ));
 sky130_fd_sc_hd__xor2_1 \U$$1987  (.A(\t$5420 ),
    .B(net1452),
    .X(booth_b28_m31));
 sky130_fd_sc_hd__a22o_1 \U$$1988  (.A1(net1016),
    .A2(net586),
    .B1(net999),
    .B2(net859),
    .X(\t$5421 ));
 sky130_fd_sc_hd__xor2_1 \U$$1989  (.A(\t$5421 ),
    .B(net1450),
    .X(booth_b28_m32));
 sky130_fd_sc_hd__a22o_1 \U$$199  (.A1(net1055),
    .A2(net619),
    .B1(net1047),
    .B2(net892),
    .X(\t$4507 ));
 sky130_fd_sc_hd__a22o_1 \U$$1990  (.A1(net1001),
    .A2(net591),
    .B1(net996),
    .B2(net864),
    .X(\t$5422 ));
 sky130_fd_sc_hd__xor2_1 \U$$1991  (.A(\t$5422 ),
    .B(net1452),
    .X(booth_b28_m33));
 sky130_fd_sc_hd__a22o_1 \U$$1992  (.A1(net991),
    .A2(net586),
    .B1(net982),
    .B2(net859),
    .X(\t$5423 ));
 sky130_fd_sc_hd__xor2_1 \U$$1993  (.A(\t$5423 ),
    .B(net1450),
    .X(booth_b28_m34));
 sky130_fd_sc_hd__a22o_1 \U$$1994  (.A1(net983),
    .A2(net586),
    .B1(net974),
    .B2(net859),
    .X(\t$5424 ));
 sky130_fd_sc_hd__xor2_1 \U$$1995  (.A(\t$5424 ),
    .B(net1450),
    .X(booth_b28_m35));
 sky130_fd_sc_hd__a22o_1 \U$$1996  (.A1(net977),
    .A2(net588),
    .B1(net969),
    .B2(net861),
    .X(\t$5425 ));
 sky130_fd_sc_hd__xor2_1 \U$$1997  (.A(\t$5425 ),
    .B(net1452),
    .X(booth_b28_m36));
 sky130_fd_sc_hd__a22o_1 \U$$1998  (.A1(net969),
    .A2(net588),
    .B1(net961),
    .B2(net861),
    .X(\t$5426 ));
 sky130_fd_sc_hd__xor2_1 \U$$1999  (.A(\t$5426 ),
    .B(net1452),
    .X(booth_b28_m37));
 sky130_fd_sc_hd__inv_1 \U$$2  (.A(net1571),
    .Y(\notblock[2] ));
 sky130_fd_sc_hd__a22o_1 \U$$20  (.A1(net1524),
    .A2(net446),
    .B1(net1516),
    .B2(net688),
    .X(\t$4417 ));
 sky130_fd_sc_hd__xor2_1 \U$$200  (.A(\t$4507 ),
    .B(net1385),
    .X(booth_b2_m28));
 sky130_fd_sc_hd__a22o_1 \U$$2000  (.A1(net961),
    .A2(net588),
    .B1(net955),
    .B2(net861),
    .X(\t$5427 ));
 sky130_fd_sc_hd__xor2_1 \U$$2001  (.A(\t$5427 ),
    .B(net1452),
    .X(booth_b28_m38));
 sky130_fd_sc_hd__a22o_1 \U$$2002  (.A1(net954),
    .A2(net591),
    .B1(net946),
    .B2(net864),
    .X(\t$5428 ));
 sky130_fd_sc_hd__xor2_1 \U$$2003  (.A(\t$5428 ),
    .B(net1455),
    .X(booth_b28_m39));
 sky130_fd_sc_hd__a22o_1 \U$$2004  (.A1(net942),
    .A2(net591),
    .B1(net926),
    .B2(net864),
    .X(\t$5429 ));
 sky130_fd_sc_hd__xor2_1 \U$$2005  (.A(\t$5429 ),
    .B(net1455),
    .X(booth_b28_m40));
 sky130_fd_sc_hd__a22o_1 \U$$2006  (.A1(net930),
    .A2(net591),
    .B1(net1751),
    .B2(net864),
    .X(\t$5430 ));
 sky130_fd_sc_hd__xor2_1 \U$$2007  (.A(\t$5430 ),
    .B(net1455),
    .X(booth_b28_m41));
 sky130_fd_sc_hd__a22o_1 \U$$2008  (.A1(net1751),
    .A2(net591),
    .B1(net1743),
    .B2(net864),
    .X(\t$5431 ));
 sky130_fd_sc_hd__xor2_1 \U$$2009  (.A(\t$5431 ),
    .B(net1455),
    .X(booth_b28_m42));
 sky130_fd_sc_hd__a22o_1 \U$$201  (.A1(net1047),
    .A2(net619),
    .B1(net1039),
    .B2(net892),
    .X(\t$4508 ));
 sky130_fd_sc_hd__a22o_1 \U$$2010  (.A1(net1738),
    .A2(net589),
    .B1(net1730),
    .B2(net862),
    .X(\t$5432 ));
 sky130_fd_sc_hd__xor2_1 \U$$2011  (.A(\t$5432 ),
    .B(net1454),
    .X(booth_b28_m43));
 sky130_fd_sc_hd__a22o_1 \U$$2012  (.A1(net1730),
    .A2(net589),
    .B1(net1721),
    .B2(net862),
    .X(\t$5433 ));
 sky130_fd_sc_hd__xor2_1 \U$$2013  (.A(\t$5433 ),
    .B(net1454),
    .X(booth_b28_m44));
 sky130_fd_sc_hd__a22o_1 \U$$2014  (.A1(net1720),
    .A2(net589),
    .B1(net1711),
    .B2(net862),
    .X(\t$5434 ));
 sky130_fd_sc_hd__xor2_1 \U$$2015  (.A(\t$5434 ),
    .B(net1450),
    .X(booth_b28_m45));
 sky130_fd_sc_hd__a22o_1 \U$$2016  (.A1(net1711),
    .A2(net586),
    .B1(net1703),
    .B2(net859),
    .X(\t$5435 ));
 sky130_fd_sc_hd__xor2_1 \U$$2017  (.A(\t$5435 ),
    .B(net1450),
    .X(booth_b28_m46));
 sky130_fd_sc_hd__a22o_1 \U$$2018  (.A1(net1704),
    .A2(net589),
    .B1(net1696),
    .B2(net862),
    .X(\t$5436 ));
 sky130_fd_sc_hd__xor2_1 \U$$2019  (.A(\t$5436 ),
    .B(net1454),
    .X(booth_b28_m47));
 sky130_fd_sc_hd__xor2_1 \U$$202  (.A(\t$4508 ),
    .B(net1385),
    .X(booth_b2_m29));
 sky130_fd_sc_hd__a22o_1 \U$$2020  (.A1(net1695),
    .A2(net589),
    .B1(net1687),
    .B2(net862),
    .X(\t$5437 ));
 sky130_fd_sc_hd__xor2_1 \U$$2021  (.A(\t$5437 ),
    .B(net1454),
    .X(booth_b28_m48));
 sky130_fd_sc_hd__a22o_1 \U$$2022  (.A1(net1692),
    .A2(net591),
    .B1(net1685),
    .B2(net864),
    .X(\t$5438 ));
 sky130_fd_sc_hd__xor2_1 \U$$2023  (.A(\t$5438 ),
    .B(net1455),
    .X(booth_b28_m49));
 sky130_fd_sc_hd__a22o_1 \U$$2024  (.A1(net1680),
    .A2(net590),
    .B1(net1655),
    .B2(net863),
    .X(\t$5439 ));
 sky130_fd_sc_hd__xor2_1 \U$$2025  (.A(\t$5439 ),
    .B(net1453),
    .X(booth_b28_m50));
 sky130_fd_sc_hd__a22o_1 \U$$2026  (.A1(net1655),
    .A2(net589),
    .B1(net1647),
    .B2(net862),
    .X(\t$5440 ));
 sky130_fd_sc_hd__xor2_1 \U$$2027  (.A(\t$5440 ),
    .B(net1454),
    .X(booth_b28_m51));
 sky130_fd_sc_hd__a22o_1 \U$$2028  (.A1(net1647),
    .A2(net589),
    .B1(net1639),
    .B2(net862),
    .X(\t$5441 ));
 sky130_fd_sc_hd__xor2_1 \U$$2029  (.A(\t$5441 ),
    .B(net1453),
    .X(booth_b28_m52));
 sky130_fd_sc_hd__a22o_1 \U$$203  (.A1(net1039),
    .A2(net620),
    .B1(net1024),
    .B2(net893),
    .X(\t$4509 ));
 sky130_fd_sc_hd__a22o_1 \U$$2030  (.A1(net1639),
    .A2(net590),
    .B1(net1631),
    .B2(net863),
    .X(\t$5442 ));
 sky130_fd_sc_hd__xor2_1 \U$$2031  (.A(\t$5442 ),
    .B(net1453),
    .X(booth_b28_m53));
 sky130_fd_sc_hd__a22o_1 \U$$2032  (.A1(net1631),
    .A2(net590),
    .B1(net1622),
    .B2(net863),
    .X(\t$5443 ));
 sky130_fd_sc_hd__xor2_1 \U$$2033  (.A(\t$5443 ),
    .B(net1454),
    .X(booth_b28_m54));
 sky130_fd_sc_hd__a22o_1 \U$$2034  (.A1(net1622),
    .A2(net589),
    .B1(net1613),
    .B2(net862),
    .X(\t$5444 ));
 sky130_fd_sc_hd__xor2_1 \U$$2035  (.A(\t$5444 ),
    .B(net1454),
    .X(booth_b28_m55));
 sky130_fd_sc_hd__a22o_1 \U$$2036  (.A1(net1613),
    .A2(net589),
    .B1(net1605),
    .B2(net862),
    .X(\t$5445 ));
 sky130_fd_sc_hd__xor2_1 \U$$2037  (.A(\t$5445 ),
    .B(net1453),
    .X(booth_b28_m56));
 sky130_fd_sc_hd__a22o_1 \U$$2038  (.A1(net1605),
    .A2(net590),
    .B1(net1597),
    .B2(net863),
    .X(\t$5446 ));
 sky130_fd_sc_hd__xor2_1 \U$$2039  (.A(\t$5446 ),
    .B(net1453),
    .X(booth_b28_m57));
 sky130_fd_sc_hd__xor2_1 \U$$204  (.A(\t$4509 ),
    .B(net1386),
    .X(booth_b2_m30));
 sky130_fd_sc_hd__a22o_1 \U$$2040  (.A1(net1597),
    .A2(net590),
    .B1(net1588),
    .B2(net863),
    .X(\t$5447 ));
 sky130_fd_sc_hd__xor2_1 \U$$2041  (.A(\t$5447 ),
    .B(net1453),
    .X(booth_b28_m58));
 sky130_fd_sc_hd__a22o_1 \U$$2042  (.A1(net1588),
    .A2(net589),
    .B1(net1579),
    .B2(net862),
    .X(\t$5448 ));
 sky130_fd_sc_hd__xor2_1 \U$$2043  (.A(\t$5448 ),
    .B(net1453),
    .X(booth_b28_m59));
 sky130_fd_sc_hd__a22o_1 \U$$2044  (.A1(net1580),
    .A2(net591),
    .B1(net1553),
    .B2(net864),
    .X(\t$5449 ));
 sky130_fd_sc_hd__xor2_1 \U$$2045  (.A(\t$5449 ),
    .B(net1455),
    .X(booth_b28_m60));
 sky130_fd_sc_hd__a22o_1 \U$$2046  (.A1(net1556),
    .A2(net591),
    .B1(net1548),
    .B2(net864),
    .X(\t$5450 ));
 sky130_fd_sc_hd__xor2_1 \U$$2047  (.A(\t$5450 ),
    .B(net1455),
    .X(booth_b28_m61));
 sky130_fd_sc_hd__a22o_1 \U$$2048  (.A1(net1548),
    .A2(net592),
    .B1(net1540),
    .B2(net865),
    .X(\t$5451 ));
 sky130_fd_sc_hd__xor2_1 \U$$2049  (.A(\t$5451 ),
    .B(net1456),
    .X(booth_b28_m62));
 sky130_fd_sc_hd__a22o_1 \U$$205  (.A1(net1025),
    .A2(net623),
    .B1(net1017),
    .B2(net896),
    .X(\t$4510 ));
 sky130_fd_sc_hd__a22o_1 \U$$2050  (.A1(net1539),
    .A2(net591),
    .B1(net1531),
    .B2(net864),
    .X(\t$5452 ));
 sky130_fd_sc_hd__xor2_1 \U$$2051  (.A(\t$5452 ),
    .B(net1455),
    .X(booth_b28_m63));
 sky130_fd_sc_hd__a22o_1 \U$$2052  (.A1(net1532),
    .A2(net591),
    .B1(net1770),
    .B2(net864),
    .X(\t$5453 ));
 sky130_fd_sc_hd__xor2_1 \U$$2053  (.A(\t$5453 ),
    .B(net1455),
    .X(booth_b28_m64));
 sky130_fd_sc_hd__inv_1 \U$$2054  (.A(net1455),
    .Y(\notsign$5454 ));
 sky130_fd_sc_hd__inv_1 \U$$2055  (.A(net1454),
    .Y(\notblock$5455[0] ));
 sky130_fd_sc_hd__inv_1 \U$$2056  (.A(net24),
    .Y(\notblock$5455[1] ));
 sky130_fd_sc_hd__inv_1 \U$$2057  (.A(net1444),
    .Y(\notblock$5455[2] ));
 sky130_fd_sc_hd__and2_1 \U$$2058  (.A(net1444),
    .B(\notblock$5455[1] ),
    .X(\t$5456 ));
 sky130_fd_sc_hd__a32o_1 \U$$2059  (.A1(\notblock$5455[2] ),
    .A2(net24),
    .A3(net1454),
    .B1(\t$5456 ),
    .B2(\notblock$5455[0] ),
    .X(\sel_0$5457 ));
 sky130_fd_sc_hd__xor2_1 \U$$206  (.A(\t$4510 ),
    .B(net1389),
    .X(booth_b2_m31));
 sky130_fd_sc_hd__xor2_1 \U$$2060  (.A(net24),
    .B(net1453),
    .X(\sel_1$5458 ));
 sky130_fd_sc_hd__a22o_1 \U$$2061  (.A1(net1771),
    .A2(net576),
    .B1(net1227),
    .B2(net849),
    .X(\t$5459 ));
 sky130_fd_sc_hd__xor2_1 \U$$2062  (.A(\t$5459 ),
    .B(net1439),
    .X(booth_b30_m0));
 sky130_fd_sc_hd__a22o_1 \U$$2063  (.A1(net1227),
    .A2(net576),
    .B1(net1122),
    .B2(net849),
    .X(\t$5460 ));
 sky130_fd_sc_hd__xor2_1 \U$$2064  (.A(\t$5460 ),
    .B(net1439),
    .X(booth_b30_m1));
 sky130_fd_sc_hd__a22o_1 \U$$2065  (.A1(net1126),
    .A2(net581),
    .B1(net1032),
    .B2(net854),
    .X(\t$5461 ));
 sky130_fd_sc_hd__xor2_1 \U$$2066  (.A(\t$5461 ),
    .B(net1441),
    .X(booth_b30_m2));
 sky130_fd_sc_hd__a22o_1 \U$$2067  (.A1(net1036),
    .A2(net581),
    .B1(net936),
    .B2(net854),
    .X(\t$5462 ));
 sky130_fd_sc_hd__xor2_1 \U$$2068  (.A(\t$5462 ),
    .B(net1441),
    .X(booth_b30_m3));
 sky130_fd_sc_hd__a22o_1 \U$$2069  (.A1(net937),
    .A2(net580),
    .B1(net1675),
    .B2(net853),
    .X(\t$5463 ));
 sky130_fd_sc_hd__a22o_1 \U$$207  (.A1(net1017),
    .A2(net623),
    .B1(net1000),
    .B2(net896),
    .X(\t$4511 ));
 sky130_fd_sc_hd__xor2_1 \U$$2070  (.A(\t$5463 ),
    .B(net1441),
    .X(booth_b30_m4));
 sky130_fd_sc_hd__a22o_1 \U$$2071  (.A1(net1675),
    .A2(net580),
    .B1(net1565),
    .B2(net853),
    .X(\t$5464 ));
 sky130_fd_sc_hd__xor2_1 \U$$2072  (.A(\t$5464 ),
    .B(net1441),
    .X(booth_b30_m5));
 sky130_fd_sc_hd__a22o_1 \U$$2073  (.A1(net1565),
    .A2(net581),
    .B1(net1524),
    .B2(net854),
    .X(\t$5465 ));
 sky130_fd_sc_hd__xor2_1 \U$$2074  (.A(\t$5465 ),
    .B(net1441),
    .X(booth_b30_m6));
 sky130_fd_sc_hd__a22o_1 \U$$2075  (.A1(net1521),
    .A2(net581),
    .B1(net1515),
    .B2(net854),
    .X(\t$5466 ));
 sky130_fd_sc_hd__xor2_1 \U$$2076  (.A(\t$5466 ),
    .B(net1441),
    .X(booth_b30_m7));
 sky130_fd_sc_hd__a22o_1 \U$$2077  (.A1(net1511),
    .A2(net576),
    .B1(net1503),
    .B2(net849),
    .X(\t$5467 ));
 sky130_fd_sc_hd__xor2_1 \U$$2078  (.A(\t$5467 ),
    .B(net1439),
    .X(booth_b30_m8));
 sky130_fd_sc_hd__a22o_1 \U$$2079  (.A1(net1505),
    .A2(net577),
    .B1(net1496),
    .B2(net850),
    .X(\t$5468 ));
 sky130_fd_sc_hd__xor2_1 \U$$208  (.A(\t$4511 ),
    .B(net1389),
    .X(booth_b2_m32));
 sky130_fd_sc_hd__xor2_1 \U$$2080  (.A(\t$5468 ),
    .B(net1439),
    .X(booth_b30_m9));
 sky130_fd_sc_hd__a22o_1 \U$$2081  (.A1(net1494),
    .A2(net577),
    .B1(net1219),
    .B2(net850),
    .X(\t$5469 ));
 sky130_fd_sc_hd__xor2_1 \U$$2082  (.A(\t$5469 ),
    .B(net1439),
    .X(booth_b30_m10));
 sky130_fd_sc_hd__a22o_1 \U$$2083  (.A1(net1220),
    .A2(net576),
    .B1(net1210),
    .B2(net849),
    .X(\t$5470 ));
 sky130_fd_sc_hd__xor2_1 \U$$2084  (.A(\t$5470 ),
    .B(net1439),
    .X(booth_b30_m11));
 sky130_fd_sc_hd__a22o_1 \U$$2085  (.A1(net1210),
    .A2(net576),
    .B1(net1201),
    .B2(net849),
    .X(\t$5471 ));
 sky130_fd_sc_hd__xor2_1 \U$$2086  (.A(\t$5471 ),
    .B(net1439),
    .X(booth_b30_m12));
 sky130_fd_sc_hd__a22o_1 \U$$2087  (.A1(net1201),
    .A2(net576),
    .B1(net1192),
    .B2(net849),
    .X(\t$5472 ));
 sky130_fd_sc_hd__xor2_1 \U$$2088  (.A(\t$5472 ),
    .B(net1439),
    .X(booth_b30_m13));
 sky130_fd_sc_hd__a22o_1 \U$$2089  (.A1(net1195),
    .A2(net577),
    .B1(net1175),
    .B2(net850),
    .X(\t$5473 ));
 sky130_fd_sc_hd__a22o_1 \U$$209  (.A1(net1000),
    .A2(net623),
    .B1(net992),
    .B2(net896),
    .X(\t$4512 ));
 sky130_fd_sc_hd__xor2_1 \U$$2090  (.A(\t$5473 ),
    .B(net1440),
    .X(booth_b30_m14));
 sky130_fd_sc_hd__a22o_1 \U$$2091  (.A1(net1176),
    .A2(net577),
    .B1(net1167),
    .B2(net850),
    .X(\t$5474 ));
 sky130_fd_sc_hd__xor2_1 \U$$2092  (.A(\t$5474 ),
    .B(net1440),
    .X(booth_b30_m15));
 sky130_fd_sc_hd__a22o_1 \U$$2093  (.A1(net1165),
    .A2(net577),
    .B1(net1156),
    .B2(net850),
    .X(\t$5475 ));
 sky130_fd_sc_hd__xor2_1 \U$$2094  (.A(\t$5475 ),
    .B(net1440),
    .X(booth_b30_m16));
 sky130_fd_sc_hd__a22o_1 \U$$2095  (.A1(net1156),
    .A2(net576),
    .B1(net1148),
    .B2(net849),
    .X(\t$5476 ));
 sky130_fd_sc_hd__xor2_1 \U$$2096  (.A(\t$5476 ),
    .B(net1440),
    .X(booth_b30_m17));
 sky130_fd_sc_hd__a22o_1 \U$$2097  (.A1(net1148),
    .A2(net576),
    .B1(net1140),
    .B2(net849),
    .X(\t$5477 ));
 sky130_fd_sc_hd__xor2_1 \U$$2098  (.A(\t$5477 ),
    .B(net1439),
    .X(booth_b30_m18));
 sky130_fd_sc_hd__a22o_1 \U$$2099  (.A1(net1139),
    .A2(net577),
    .B1(net1132),
    .B2(net850),
    .X(\t$5478 ));
 sky130_fd_sc_hd__xor2_1 \U$$21  (.A(\t$4417 ),
    .B(net1573),
    .X(booth_b0_m7));
 sky130_fd_sc_hd__xor2_1 \U$$210  (.A(\t$4512 ),
    .B(net1389),
    .X(booth_b2_m33));
 sky130_fd_sc_hd__xor2_1 \U$$2100  (.A(\t$5478 ),
    .B(net1440),
    .X(booth_b30_m19));
 sky130_fd_sc_hd__a22o_1 \U$$2101  (.A1(net1134),
    .A2(net580),
    .B1(net1117),
    .B2(net853),
    .X(\t$5479 ));
 sky130_fd_sc_hd__xor2_1 \U$$2102  (.A(\t$5479 ),
    .B(net1441),
    .X(booth_b30_m20));
 sky130_fd_sc_hd__a22o_1 \U$$2103  (.A1(net1118),
    .A2(net580),
    .B1(net1109),
    .B2(net853),
    .X(\t$5480 ));
 sky130_fd_sc_hd__xor2_1 \U$$2104  (.A(\t$5480 ),
    .B(net1441),
    .X(booth_b30_m21));
 sky130_fd_sc_hd__a22o_1 \U$$2105  (.A1(net1108),
    .A2(net580),
    .B1(net1100),
    .B2(net853),
    .X(\t$5481 ));
 sky130_fd_sc_hd__xor2_1 \U$$2106  (.A(\t$5481 ),
    .B(net1441),
    .X(booth_b30_m22));
 sky130_fd_sc_hd__a22o_1 \U$$2107  (.A1(net1100),
    .A2(net580),
    .B1(net1091),
    .B2(net853),
    .X(\t$5482 ));
 sky130_fd_sc_hd__xor2_1 \U$$2108  (.A(\t$5482 ),
    .B(net1442),
    .X(booth_b30_m23));
 sky130_fd_sc_hd__a22o_1 \U$$2109  (.A1(net1092),
    .A2(net580),
    .B1(net1083),
    .B2(net853),
    .X(\t$5483 ));
 sky130_fd_sc_hd__a22o_1 \U$$211  (.A1(net992),
    .A2(net625),
    .B1(net987),
    .B2(net898),
    .X(\t$4513 ));
 sky130_fd_sc_hd__xor2_1 \U$$2110  (.A(\t$5483 ),
    .B(net1442),
    .X(booth_b30_m24));
 sky130_fd_sc_hd__a22o_1 \U$$2111  (.A1(net1084),
    .A2(net580),
    .B1(net1074),
    .B2(net853),
    .X(\t$5484 ));
 sky130_fd_sc_hd__xor2_1 \U$$2112  (.A(\t$5484 ),
    .B(net1442),
    .X(booth_b30_m25));
 sky130_fd_sc_hd__a22o_1 \U$$2113  (.A1(net1075),
    .A2(net581),
    .B1(net1067),
    .B2(net854),
    .X(\t$5485 ));
 sky130_fd_sc_hd__xor2_1 \U$$2114  (.A(\t$5485 ),
    .B(net1442),
    .X(booth_b30_m26));
 sky130_fd_sc_hd__a22o_1 \U$$2115  (.A1(net1066),
    .A2(net581),
    .B1(net1057),
    .B2(net854),
    .X(\t$5486 ));
 sky130_fd_sc_hd__xor2_1 \U$$2116  (.A(\t$5486 ),
    .B(net1441),
    .X(booth_b30_m27));
 sky130_fd_sc_hd__a22o_1 \U$$2117  (.A1(net1058),
    .A2(net581),
    .B1(net1050),
    .B2(net854),
    .X(\t$5487 ));
 sky130_fd_sc_hd__xor2_1 \U$$2118  (.A(\t$5487 ),
    .B(net1442),
    .X(booth_b30_m28));
 sky130_fd_sc_hd__a22o_1 \U$$2119  (.A1(net1050),
    .A2(net581),
    .B1(net1042),
    .B2(net854),
    .X(\t$5488 ));
 sky130_fd_sc_hd__xor2_1 \U$$212  (.A(\t$4513 ),
    .B(net1391),
    .X(booth_b2_m34));
 sky130_fd_sc_hd__xor2_1 \U$$2120  (.A(\t$5488 ),
    .B(net1442),
    .X(booth_b30_m29));
 sky130_fd_sc_hd__a22o_1 \U$$2121  (.A1(net1040),
    .A2(net577),
    .B1(net1024),
    .B2(net850),
    .X(\t$5489 ));
 sky130_fd_sc_hd__xor2_1 \U$$2122  (.A(\t$5489 ),
    .B(net1440),
    .X(booth_b30_m30));
 sky130_fd_sc_hd__a22o_1 \U$$2123  (.A1(net1026),
    .A2(net582),
    .B1(net1018),
    .B2(net855),
    .X(\t$5490 ));
 sky130_fd_sc_hd__xor2_1 \U$$2124  (.A(\t$5490 ),
    .B(net1442),
    .X(booth_b30_m31));
 sky130_fd_sc_hd__a22o_1 \U$$2125  (.A1(net1016),
    .A2(net576),
    .B1(net999),
    .B2(net849),
    .X(\t$5491 ));
 sky130_fd_sc_hd__xor2_1 \U$$2126  (.A(\t$5491 ),
    .B(net1440),
    .X(booth_b30_m32));
 sky130_fd_sc_hd__a22o_1 \U$$2127  (.A1(net999),
    .A2(net579),
    .B1(net991),
    .B2(net852),
    .X(\t$5492 ));
 sky130_fd_sc_hd__xor2_1 \U$$2128  (.A(\t$5492 ),
    .B(net1440),
    .X(booth_b30_m33));
 sky130_fd_sc_hd__a22o_1 \U$$2129  (.A1(net991),
    .A2(net581),
    .B1(net983),
    .B2(net854),
    .X(\t$5493 ));
 sky130_fd_sc_hd__a22o_1 \U$$213  (.A1(net982),
    .A2(net619),
    .B1(net973),
    .B2(net892),
    .X(\t$4514 ));
 sky130_fd_sc_hd__xor2_1 \U$$2130  (.A(\t$5493 ),
    .B(net1442),
    .X(booth_b30_m34));
 sky130_fd_sc_hd__a22o_1 \U$$2131  (.A1(net989),
    .A2(net580),
    .B1(net978),
    .B2(net853),
    .X(\t$5494 ));
 sky130_fd_sc_hd__xor2_1 \U$$2132  (.A(\t$5494 ),
    .B(net1442),
    .X(booth_b30_m35));
 sky130_fd_sc_hd__a22o_1 \U$$2133  (.A1(net978),
    .A2(net580),
    .B1(net972),
    .B2(net853),
    .X(\t$5495 ));
 sky130_fd_sc_hd__xor2_1 \U$$2134  (.A(\t$5495 ),
    .B(net1443),
    .X(booth_b30_m36));
 sky130_fd_sc_hd__a22o_1 \U$$2135  (.A1(net972),
    .A2(net582),
    .B1(net963),
    .B2(net855),
    .X(\t$5496 ));
 sky130_fd_sc_hd__xor2_1 \U$$2136  (.A(\t$5496 ),
    .B(net1443),
    .X(booth_b30_m37));
 sky130_fd_sc_hd__a22o_1 \U$$2137  (.A1(net958),
    .A2(net582),
    .B1(net950),
    .B2(net855),
    .X(\t$5497 ));
 sky130_fd_sc_hd__xor2_1 \U$$2138  (.A(\t$5497 ),
    .B(net1446),
    .X(booth_b30_m38));
 sky130_fd_sc_hd__a22o_1 \U$$2139  (.A1(net954),
    .A2(net583),
    .B1(net946),
    .B2(net856),
    .X(\t$5498 ));
 sky130_fd_sc_hd__xor2_1 \U$$214  (.A(\t$4514 ),
    .B(net1385),
    .X(booth_b2_m35));
 sky130_fd_sc_hd__xor2_1 \U$$2140  (.A(\t$5498 ),
    .B(net1446),
    .X(booth_b30_m39));
 sky130_fd_sc_hd__a22o_1 \U$$2141  (.A1(net946),
    .A2(net582),
    .B1(net930),
    .B2(net855),
    .X(\t$5499 ));
 sky130_fd_sc_hd__xor2_1 \U$$2142  (.A(\t$5499 ),
    .B(net1446),
    .X(booth_b30_m40));
 sky130_fd_sc_hd__a22o_1 \U$$2143  (.A1(net926),
    .A2(net579),
    .B1(net1748),
    .B2(net852),
    .X(\t$5500 ));
 sky130_fd_sc_hd__xor2_1 \U$$2144  (.A(\t$5500 ),
    .B(net1445),
    .X(booth_b30_m41));
 sky130_fd_sc_hd__a22o_1 \U$$2145  (.A1(net1746),
    .A2(net579),
    .B1(net1738),
    .B2(net852),
    .X(\t$5501 ));
 sky130_fd_sc_hd__xor2_1 \U$$2146  (.A(\t$5501 ),
    .B(net1445),
    .X(booth_b30_m42));
 sky130_fd_sc_hd__a22o_1 \U$$2147  (.A1(net1737),
    .A2(net578),
    .B1(net1729),
    .B2(net851),
    .X(\t$5502 ));
 sky130_fd_sc_hd__xor2_1 \U$$2148  (.A(\t$5502 ),
    .B(net1440),
    .X(booth_b30_m43));
 sky130_fd_sc_hd__a22o_1 \U$$2149  (.A1(net1729),
    .A2(net576),
    .B1(net1720),
    .B2(net849),
    .X(\t$5503 ));
 sky130_fd_sc_hd__a22o_1 \U$$215  (.A1(net974),
    .A2(net625),
    .B1(net965),
    .B2(net898),
    .X(\t$4515 ));
 sky130_fd_sc_hd__xor2_1 \U$$2150  (.A(\t$5503 ),
    .B(net1443),
    .X(booth_b30_m44));
 sky130_fd_sc_hd__a22o_1 \U$$2151  (.A1(net1722),
    .A2(net578),
    .B1(net1713),
    .B2(net851),
    .X(\t$5504 ));
 sky130_fd_sc_hd__xor2_1 \U$$2152  (.A(\t$5504 ),
    .B(net1445),
    .X(booth_b30_m45));
 sky130_fd_sc_hd__a22o_1 \U$$2153  (.A1(net1713),
    .A2(net578),
    .B1(net1704),
    .B2(net851),
    .X(\t$5505 ));
 sky130_fd_sc_hd__xor2_1 \U$$2154  (.A(\t$5505 ),
    .B(net1445),
    .X(booth_b30_m46));
 sky130_fd_sc_hd__a22o_1 \U$$2155  (.A1(net1705),
    .A2(net579),
    .B1(net1697),
    .B2(net852),
    .X(\t$5506 ));
 sky130_fd_sc_hd__xor2_1 \U$$2156  (.A(\t$5506 ),
    .B(net1445),
    .X(booth_b30_m47));
 sky130_fd_sc_hd__a22o_1 \U$$2157  (.A1(net1696),
    .A2(net579),
    .B1(net1688),
    .B2(net852),
    .X(\t$5507 ));
 sky130_fd_sc_hd__xor2_1 \U$$2158  (.A(\t$5507 ),
    .B(net1446),
    .X(booth_b30_m48));
 sky130_fd_sc_hd__a22o_1 \U$$2159  (.A1(net1688),
    .A2(net579),
    .B1(net1680),
    .B2(net852),
    .X(\t$5508 ));
 sky130_fd_sc_hd__xor2_1 \U$$216  (.A(\t$4515 ),
    .B(net1386),
    .X(booth_b2_m36));
 sky130_fd_sc_hd__xor2_1 \U$$2160  (.A(\t$5508 ),
    .B(net1445),
    .X(booth_b30_m49));
 sky130_fd_sc_hd__a22o_1 \U$$2161  (.A1(net1680),
    .A2(net578),
    .B1(net1655),
    .B2(net851),
    .X(\t$5509 ));
 sky130_fd_sc_hd__xor2_1 \U$$2162  (.A(\t$5509 ),
    .B(net1444),
    .X(booth_b30_m50));
 sky130_fd_sc_hd__a22o_1 \U$$2163  (.A1(net1655),
    .A2(net579),
    .B1(net1647),
    .B2(net852),
    .X(\t$5510 ));
 sky130_fd_sc_hd__xor2_1 \U$$2164  (.A(\t$5510 ),
    .B(net1446),
    .X(booth_b30_m51));
 sky130_fd_sc_hd__a22o_1 \U$$2165  (.A1(net1647),
    .A2(net578),
    .B1(net1639),
    .B2(net851),
    .X(\t$5511 ));
 sky130_fd_sc_hd__xor2_1 \U$$2166  (.A(\t$5511 ),
    .B(net1445),
    .X(booth_b30_m52));
 sky130_fd_sc_hd__a22o_1 \U$$2167  (.A1(net1639),
    .A2(net578),
    .B1(net1631),
    .B2(net851),
    .X(\t$5512 ));
 sky130_fd_sc_hd__xor2_1 \U$$2168  (.A(\t$5512 ),
    .B(net1445),
    .X(booth_b30_m53));
 sky130_fd_sc_hd__a22o_1 \U$$2169  (.A1(net1631),
    .A2(net578),
    .B1(net1622),
    .B2(net851),
    .X(\t$5513 ));
 sky130_fd_sc_hd__a22o_1 \U$$217  (.A1(net968),
    .A2(net625),
    .B1(net957),
    .B2(net898),
    .X(\t$4516 ));
 sky130_fd_sc_hd__xor2_1 \U$$2170  (.A(\t$5513 ),
    .B(net1444),
    .X(booth_b30_m54));
 sky130_fd_sc_hd__a22o_1 \U$$2171  (.A1(net1622),
    .A2(net578),
    .B1(net1613),
    .B2(net851),
    .X(\t$5514 ));
 sky130_fd_sc_hd__xor2_1 \U$$2172  (.A(\t$5514 ),
    .B(net1444),
    .X(booth_b30_m55));
 sky130_fd_sc_hd__a22o_1 \U$$2173  (.A1(net1613),
    .A2(net578),
    .B1(net1605),
    .B2(net851),
    .X(\t$5515 ));
 sky130_fd_sc_hd__xor2_1 \U$$2174  (.A(\t$5515 ),
    .B(net1444),
    .X(booth_b30_m56));
 sky130_fd_sc_hd__a22o_1 \U$$2175  (.A1(net1605),
    .A2(net578),
    .B1(net1597),
    .B2(net851),
    .X(\t$5516 ));
 sky130_fd_sc_hd__xor2_1 \U$$2176  (.A(\t$5516 ),
    .B(net1444),
    .X(booth_b30_m57));
 sky130_fd_sc_hd__a22o_1 \U$$2177  (.A1(net1598),
    .A2(net582),
    .B1(net1589),
    .B2(net855),
    .X(\t$5517 ));
 sky130_fd_sc_hd__xor2_1 \U$$2178  (.A(\t$5517 ),
    .B(net1446),
    .X(booth_b30_m58));
 sky130_fd_sc_hd__a22o_1 \U$$2179  (.A1(net1589),
    .A2(net579),
    .B1(net1580),
    .B2(net852),
    .X(\t$5518 ));
 sky130_fd_sc_hd__xor2_1 \U$$218  (.A(\t$4516 ),
    .B(net1391),
    .X(booth_b2_m37));
 sky130_fd_sc_hd__xor2_1 \U$$2180  (.A(\t$5518 ),
    .B(net1445),
    .X(booth_b30_m59));
 sky130_fd_sc_hd__a22o_1 \U$$2181  (.A1(net1580),
    .A2(net579),
    .B1(net1554),
    .B2(net852),
    .X(\t$5519 ));
 sky130_fd_sc_hd__xor2_1 \U$$2182  (.A(\t$5519 ),
    .B(net1446),
    .X(booth_b30_m60));
 sky130_fd_sc_hd__a22o_1 \U$$2183  (.A1(net1555),
    .A2(net582),
    .B1(net1547),
    .B2(net855),
    .X(\t$5520 ));
 sky130_fd_sc_hd__xor2_1 \U$$2184  (.A(\t$5520 ),
    .B(net1446),
    .X(booth_b30_m61));
 sky130_fd_sc_hd__a22o_1 \U$$2185  (.A1(net1548),
    .A2(net582),
    .B1(net1540),
    .B2(net855),
    .X(\t$5521 ));
 sky130_fd_sc_hd__xor2_1 \U$$2186  (.A(\t$5521 ),
    .B(net1446),
    .X(booth_b30_m62));
 sky130_fd_sc_hd__a22o_1 \U$$2187  (.A1(net1539),
    .A2(net582),
    .B1(net1531),
    .B2(net855),
    .X(\t$5522 ));
 sky130_fd_sc_hd__xor2_1 \U$$2188  (.A(\t$5522 ),
    .B(net1447),
    .X(booth_b30_m63));
 sky130_fd_sc_hd__a22o_1 \U$$2189  (.A1(net1531),
    .A2(net582),
    .B1(net1772),
    .B2(net855),
    .X(\t$5523 ));
 sky130_fd_sc_hd__a22o_1 \U$$219  (.A1(net956),
    .A2(net619),
    .B1(net948),
    .B2(net892),
    .X(\t$4517 ));
 sky130_fd_sc_hd__xor2_1 \U$$2190  (.A(\t$5523 ),
    .B(net1447),
    .X(booth_b30_m64));
 sky130_fd_sc_hd__inv_1 \U$$2191  (.A(net1447),
    .Y(\notsign$5524 ));
 sky130_fd_sc_hd__inv_1 \U$$2192  (.A(net1444),
    .Y(\notblock$5525[0] ));
 sky130_fd_sc_hd__inv_1 \U$$2193  (.A(net26),
    .Y(\notblock$5525[1] ));
 sky130_fd_sc_hd__inv_1 \U$$2194  (.A(net1435),
    .Y(\notblock$5525[2] ));
 sky130_fd_sc_hd__and2_1 \U$$2195  (.A(net1435),
    .B(\notblock$5525[1] ),
    .X(\t$5526 ));
 sky130_fd_sc_hd__a32o_4 \U$$2196  (.A1(\notblock$5525[2] ),
    .A2(net26),
    .A3(net1444),
    .B1(\t$5526 ),
    .B2(\notblock$5525[0] ),
    .X(\sel_0$5527 ));
 sky130_fd_sc_hd__xor2_4 \U$$2197  (.A(net26),
    .B(net1444),
    .X(\sel_1$5528 ));
 sky130_fd_sc_hd__a22o_1 \U$$2198  (.A1(net1773),
    .A2(net571),
    .B1(net1230),
    .B2(net844),
    .X(\t$5529 ));
 sky130_fd_sc_hd__xor2_1 \U$$2199  (.A(\t$5529 ),
    .B(net1432),
    .X(booth_b32_m0));
 sky130_fd_sc_hd__a22o_1 \U$$22  (.A1(net1515),
    .A2(net446),
    .B1(net1508),
    .B2(net688),
    .X(\t$4418 ));
 sky130_fd_sc_hd__xor2_1 \U$$220  (.A(\t$4517 ),
    .B(net1385),
    .X(booth_b2_m38));
 sky130_fd_sc_hd__a22o_1 \U$$2200  (.A1(net1230),
    .A2(net571),
    .B1(net1126),
    .B2(net844),
    .X(\t$5530 ));
 sky130_fd_sc_hd__xor2_1 \U$$2201  (.A(\t$5530 ),
    .B(net1432),
    .X(booth_b32_m1));
 sky130_fd_sc_hd__a22o_1 \U$$2202  (.A1(net1128),
    .A2(net572),
    .B1(net1035),
    .B2(net845),
    .X(\t$5531 ));
 sky130_fd_sc_hd__xor2_1 \U$$2203  (.A(\t$5531 ),
    .B(net1432),
    .X(booth_b32_m2));
 sky130_fd_sc_hd__a22o_1 \U$$2204  (.A1(net1038),
    .A2(net572),
    .B1(net937),
    .B2(net845),
    .X(\t$5532 ));
 sky130_fd_sc_hd__xor2_1 \U$$2205  (.A(\t$5532 ),
    .B(net1432),
    .X(booth_b32_m3));
 sky130_fd_sc_hd__a22o_1 \U$$2206  (.A1(net936),
    .A2(net571),
    .B1(net1676),
    .B2(net844),
    .X(\t$5533 ));
 sky130_fd_sc_hd__xor2_1 \U$$2207  (.A(\t$5533 ),
    .B(net1432),
    .X(booth_b32_m4));
 sky130_fd_sc_hd__a22o_1 \U$$2208  (.A1(net1676),
    .A2(net571),
    .B1(net1561),
    .B2(net844),
    .X(\t$5534 ));
 sky130_fd_sc_hd__xor2_1 \U$$2209  (.A(\t$5534 ),
    .B(net1432),
    .X(booth_b32_m5));
 sky130_fd_sc_hd__a22o_1 \U$$221  (.A1(net948),
    .A2(net619),
    .B1(net940),
    .B2(net892),
    .X(\t$4518 ));
 sky130_fd_sc_hd__a22o_1 \U$$2210  (.A1(net1560),
    .A2(net569),
    .B1(net1519),
    .B2(net842),
    .X(\t$5535 ));
 sky130_fd_sc_hd__xor2_1 \U$$2211  (.A(\t$5535 ),
    .B(net1430),
    .X(booth_b32_m6));
 sky130_fd_sc_hd__a22o_1 \U$$2212  (.A1(net1521),
    .A2(net569),
    .B1(net1513),
    .B2(net842),
    .X(\t$5536 ));
 sky130_fd_sc_hd__xor2_1 \U$$2213  (.A(\t$5536 ),
    .B(net1430),
    .X(booth_b32_m7));
 sky130_fd_sc_hd__a22o_1 \U$$2214  (.A1(net1511),
    .A2(net569),
    .B1(net1503),
    .B2(net842),
    .X(\t$5537 ));
 sky130_fd_sc_hd__xor2_1 \U$$2215  (.A(\t$5537 ),
    .B(net1430),
    .X(booth_b32_m8));
 sky130_fd_sc_hd__a22o_1 \U$$2216  (.A1(net1503),
    .A2(net569),
    .B1(net1495),
    .B2(net842),
    .X(\t$5538 ));
 sky130_fd_sc_hd__xor2_1 \U$$2217  (.A(\t$5538 ),
    .B(net1430),
    .X(booth_b32_m9));
 sky130_fd_sc_hd__a22o_1 \U$$2218  (.A1(net1494),
    .A2(net569),
    .B1(net1219),
    .B2(net842),
    .X(\t$5539 ));
 sky130_fd_sc_hd__xor2_1 \U$$2219  (.A(\t$5539 ),
    .B(net1430),
    .X(booth_b32_m10));
 sky130_fd_sc_hd__xor2_1 \U$$222  (.A(\t$4518 ),
    .B(net1385),
    .X(booth_b2_m39));
 sky130_fd_sc_hd__a22o_1 \U$$2220  (.A1(net1220),
    .A2(net569),
    .B1(net1210),
    .B2(net842),
    .X(\t$5540 ));
 sky130_fd_sc_hd__xor2_1 \U$$2221  (.A(\t$5540 ),
    .B(net1430),
    .X(booth_b32_m11));
 sky130_fd_sc_hd__a22o_1 \U$$2222  (.A1(net1212),
    .A2(net569),
    .B1(net1204),
    .B2(net842),
    .X(\t$5541 ));
 sky130_fd_sc_hd__xor2_1 \U$$2223  (.A(\t$5541 ),
    .B(net1430),
    .X(booth_b32_m12));
 sky130_fd_sc_hd__a22o_1 \U$$2224  (.A1(net1203),
    .A2(net570),
    .B1(net1194),
    .B2(net843),
    .X(\t$5542 ));
 sky130_fd_sc_hd__xor2_1 \U$$2225  (.A(\t$5542 ),
    .B(net1431),
    .X(booth_b32_m13));
 sky130_fd_sc_hd__a22o_1 \U$$2226  (.A1(net1193),
    .A2(net569),
    .B1(net1174),
    .B2(net842),
    .X(\t$5543 ));
 sky130_fd_sc_hd__xor2_1 \U$$2227  (.A(\t$5543 ),
    .B(net1430),
    .X(booth_b32_m14));
 sky130_fd_sc_hd__a22o_1 \U$$2228  (.A1(net1174),
    .A2(net570),
    .B1(net1165),
    .B2(net843),
    .X(\t$5544 ));
 sky130_fd_sc_hd__xor2_1 \U$$2229  (.A(\t$5544 ),
    .B(net1431),
    .X(booth_b32_m15));
 sky130_fd_sc_hd__a22o_1 \U$$223  (.A1(net940),
    .A2(net619),
    .B1(net924),
    .B2(net892),
    .X(\t$4519 ));
 sky130_fd_sc_hd__a22o_1 \U$$2230  (.A1(net1165),
    .A2(net569),
    .B1(net1156),
    .B2(net842),
    .X(\t$5545 ));
 sky130_fd_sc_hd__xor2_1 \U$$2231  (.A(\t$5545 ),
    .B(net1430),
    .X(booth_b32_m16));
 sky130_fd_sc_hd__a22o_1 \U$$2232  (.A1(net1158),
    .A2(net569),
    .B1(net1148),
    .B2(net842),
    .X(\t$5546 ));
 sky130_fd_sc_hd__xor2_1 \U$$2233  (.A(\t$5546 ),
    .B(net1431),
    .X(booth_b32_m17));
 sky130_fd_sc_hd__a22o_1 \U$$2234  (.A1(net1150),
    .A2(net571),
    .B1(net1144),
    .B2(net844),
    .X(\t$5547 ));
 sky130_fd_sc_hd__xor2_1 \U$$2235  (.A(\t$5547 ),
    .B(net1432),
    .X(booth_b32_m18));
 sky130_fd_sc_hd__a22o_1 \U$$2236  (.A1(net1144),
    .A2(net571),
    .B1(net1134),
    .B2(net844),
    .X(\t$5548 ));
 sky130_fd_sc_hd__xor2_1 \U$$2237  (.A(\t$5548 ),
    .B(net1432),
    .X(booth_b32_m19));
 sky130_fd_sc_hd__a22o_1 \U$$2238  (.A1(net1133),
    .A2(net571),
    .B1(net1117),
    .B2(net844),
    .X(\t$5549 ));
 sky130_fd_sc_hd__xor2_1 \U$$2239  (.A(\t$5549 ),
    .B(net1432),
    .X(booth_b32_m20));
 sky130_fd_sc_hd__xor2_1 \U$$224  (.A(\t$4519 ),
    .B(net1385),
    .X(booth_b2_m40));
 sky130_fd_sc_hd__a22o_1 \U$$2240  (.A1(net1118),
    .A2(net571),
    .B1(net1108),
    .B2(net844),
    .X(\t$5550 ));
 sky130_fd_sc_hd__xor2_1 \U$$2241  (.A(\t$5550 ),
    .B(net1433),
    .X(booth_b32_m21));
 sky130_fd_sc_hd__a22o_1 \U$$2242  (.A1(net1108),
    .A2(net571),
    .B1(net1101),
    .B2(net844),
    .X(\t$5551 ));
 sky130_fd_sc_hd__xor2_1 \U$$2243  (.A(\t$5551 ),
    .B(net1433),
    .X(booth_b32_m22));
 sky130_fd_sc_hd__a22o_1 \U$$2244  (.A1(net1101),
    .A2(net571),
    .B1(net1092),
    .B2(net844),
    .X(\t$5552 ));
 sky130_fd_sc_hd__xor2_1 \U$$2245  (.A(\t$5552 ),
    .B(net1433),
    .X(booth_b32_m23));
 sky130_fd_sc_hd__a22o_1 \U$$2246  (.A1(net1092),
    .A2(net572),
    .B1(net1084),
    .B2(net845),
    .X(\t$5553 ));
 sky130_fd_sc_hd__xor2_1 \U$$2247  (.A(\t$5553 ),
    .B(net1433),
    .X(booth_b32_m24));
 sky130_fd_sc_hd__a22o_1 \U$$2248  (.A1(net1083),
    .A2(net570),
    .B1(net1074),
    .B2(net843),
    .X(\t$5554 ));
 sky130_fd_sc_hd__xor2_1 \U$$2249  (.A(\t$5554 ),
    .B(net1432),
    .X(booth_b32_m25));
 sky130_fd_sc_hd__a22o_1 \U$$225  (.A1(net924),
    .A2(net621),
    .B1(net1745),
    .B2(net894),
    .X(\t$4520 ));
 sky130_fd_sc_hd__a22o_1 \U$$2250  (.A1(net1075),
    .A2(net572),
    .B1(net1067),
    .B2(net845),
    .X(\t$5555 ));
 sky130_fd_sc_hd__xor2_1 \U$$2251  (.A(\t$5555 ),
    .B(net1433),
    .X(booth_b32_m26));
 sky130_fd_sc_hd__a22o_1 \U$$2252  (.A1(net1067),
    .A2(net572),
    .B1(net1058),
    .B2(net845),
    .X(\t$5556 ));
 sky130_fd_sc_hd__xor2_1 \U$$2253  (.A(\t$5556 ),
    .B(net1433),
    .X(booth_b32_m27));
 sky130_fd_sc_hd__a22o_1 \U$$2254  (.A1(net1056),
    .A2(net570),
    .B1(net1048),
    .B2(net843),
    .X(\t$5557 ));
 sky130_fd_sc_hd__xor2_1 \U$$2255  (.A(\t$5557 ),
    .B(net1431),
    .X(booth_b32_m28));
 sky130_fd_sc_hd__a22o_1 \U$$2256  (.A1(net1050),
    .A2(net572),
    .B1(net1042),
    .B2(net845),
    .X(\t$5558 ));
 sky130_fd_sc_hd__xor2_1 \U$$2257  (.A(\t$5558 ),
    .B(net1433),
    .X(booth_b32_m29));
 sky130_fd_sc_hd__a22o_1 \U$$2258  (.A1(net1040),
    .A2(net570),
    .B1(net1024),
    .B2(net843),
    .X(\t$5559 ));
 sky130_fd_sc_hd__xor2_1 \U$$2259  (.A(\t$5559 ),
    .B(net1431),
    .X(booth_b32_m30));
 sky130_fd_sc_hd__xor2_1 \U$$226  (.A(\t$4520 ),
    .B(net1387),
    .X(booth_b2_m41));
 sky130_fd_sc_hd__a22o_1 \U$$2260  (.A1(net1024),
    .A2(\sel_0$5527 ),
    .B1(net1016),
    .B2(\sel_1$5528 ),
    .X(\t$5560 ));
 sky130_fd_sc_hd__xor2_1 \U$$2261  (.A(\t$5560 ),
    .B(net1431),
    .X(booth_b32_m31));
 sky130_fd_sc_hd__a22o_1 \U$$2262  (.A1(net1018),
    .A2(net570),
    .B1(net1001),
    .B2(net843),
    .X(\t$5561 ));
 sky130_fd_sc_hd__xor2_1 \U$$2263  (.A(\t$5561 ),
    .B(net1431),
    .X(booth_b32_m32));
 sky130_fd_sc_hd__a22o_1 \U$$2264  (.A1(net1001),
    .A2(net572),
    .B1(net993),
    .B2(net845),
    .X(\t$5562 ));
 sky130_fd_sc_hd__xor2_1 \U$$2265  (.A(\t$5562 ),
    .B(net1433),
    .X(booth_b32_m33));
 sky130_fd_sc_hd__a22o_1 \U$$2266  (.A1(net993),
    .A2(net572),
    .B1(net989),
    .B2(net845),
    .X(\t$5563 ));
 sky130_fd_sc_hd__xor2_1 \U$$2267  (.A(\t$5563 ),
    .B(net1433),
    .X(booth_b32_m34));
 sky130_fd_sc_hd__a22o_1 \U$$2268  (.A1(net989),
    .A2(net572),
    .B1(net978),
    .B2(net845),
    .X(\t$5564 ));
 sky130_fd_sc_hd__xor2_1 \U$$2269  (.A(\t$5564 ),
    .B(net1438),
    .X(booth_b32_m35));
 sky130_fd_sc_hd__a22o_1 \U$$227  (.A1(net1745),
    .A2(net622),
    .B1(net1737),
    .B2(net895),
    .X(\t$4521 ));
 sky130_fd_sc_hd__a22o_1 \U$$2270  (.A1(net979),
    .A2(net575),
    .B1(net970),
    .B2(net848),
    .X(\t$5565 ));
 sky130_fd_sc_hd__xor2_1 \U$$2271  (.A(\t$5565 ),
    .B(net1437),
    .X(booth_b32_m36));
 sky130_fd_sc_hd__a22o_1 \U$$2272  (.A1(net970),
    .A2(net575),
    .B1(net962),
    .B2(net848),
    .X(\t$5566 ));
 sky130_fd_sc_hd__xor2_1 \U$$2273  (.A(\t$5566 ),
    .B(net1437),
    .X(booth_b32_m37));
 sky130_fd_sc_hd__a22o_1 \U$$2274  (.A1(net958),
    .A2(net573),
    .B1(net950),
    .B2(net846),
    .X(\t$5567 ));
 sky130_fd_sc_hd__xor2_1 \U$$2275  (.A(\t$5567 ),
    .B(net1434),
    .X(booth_b32_m38));
 sky130_fd_sc_hd__a22o_1 \U$$2276  (.A1(net951),
    .A2(net573),
    .B1(net942),
    .B2(net846),
    .X(\t$5568 ));
 sky130_fd_sc_hd__xor2_1 \U$$2277  (.A(\t$5568 ),
    .B(net1434),
    .X(booth_b32_m39));
 sky130_fd_sc_hd__a22o_1 \U$$2278  (.A1(net941),
    .A2(net570),
    .B1(net925),
    .B2(net843),
    .X(\t$5569 ));
 sky130_fd_sc_hd__xor2_1 \U$$2279  (.A(\t$5569 ),
    .B(net1431),
    .X(booth_b32_m40));
 sky130_fd_sc_hd__xor2_1 \U$$228  (.A(\t$4521 ),
    .B(net1388),
    .X(booth_b2_m42));
 sky130_fd_sc_hd__a22o_1 \U$$2280  (.A1(net925),
    .A2(net570),
    .B1(net1746),
    .B2(net843),
    .X(\t$5570 ));
 sky130_fd_sc_hd__xor2_1 \U$$2281  (.A(\t$5570 ),
    .B(net1431),
    .X(booth_b32_m41));
 sky130_fd_sc_hd__a22o_1 \U$$2282  (.A1(net1746),
    .A2(net570),
    .B1(net1738),
    .B2(net843),
    .X(\t$5571 ));
 sky130_fd_sc_hd__xor2_1 \U$$2283  (.A(\t$5571 ),
    .B(net1438),
    .X(booth_b32_m42));
 sky130_fd_sc_hd__a22o_1 \U$$2284  (.A1(net1739),
    .A2(net573),
    .B1(net1731),
    .B2(net846),
    .X(\t$5572 ));
 sky130_fd_sc_hd__xor2_1 \U$$2285  (.A(\t$5572 ),
    .B(net1434),
    .X(booth_b32_m43));
 sky130_fd_sc_hd__a22o_1 \U$$2286  (.A1(net1731),
    .A2(net573),
    .B1(net1722),
    .B2(net846),
    .X(\t$5573 ));
 sky130_fd_sc_hd__xor2_1 \U$$2287  (.A(\t$5573 ),
    .B(net1434),
    .X(booth_b32_m44));
 sky130_fd_sc_hd__a22o_1 \U$$2288  (.A1(net1721),
    .A2(net573),
    .B1(net1712),
    .B2(net846),
    .X(\t$5574 ));
 sky130_fd_sc_hd__xor2_1 \U$$2289  (.A(\t$5574 ),
    .B(net1434),
    .X(booth_b32_m45));
 sky130_fd_sc_hd__a22o_1 \U$$229  (.A1(net1738),
    .A2(net622),
    .B1(net1730),
    .B2(net895),
    .X(\t$4522 ));
 sky130_fd_sc_hd__a22o_1 \U$$2290  (.A1(net1713),
    .A2(net574),
    .B1(net1704),
    .B2(net847),
    .X(\t$5575 ));
 sky130_fd_sc_hd__xor2_1 \U$$2291  (.A(\t$5575 ),
    .B(net1435),
    .X(booth_b32_m46));
 sky130_fd_sc_hd__a22o_1 \U$$2292  (.A1(net1704),
    .A2(net573),
    .B1(net1696),
    .B2(net846),
    .X(\t$5576 ));
 sky130_fd_sc_hd__xor2_1 \U$$2293  (.A(\t$5576 ),
    .B(net1434),
    .X(booth_b32_m47));
 sky130_fd_sc_hd__a22o_1 \U$$2294  (.A1(net1696),
    .A2(net573),
    .B1(net1688),
    .B2(net846),
    .X(\t$5577 ));
 sky130_fd_sc_hd__xor2_1 \U$$2295  (.A(\t$5577 ),
    .B(net1434),
    .X(booth_b32_m48));
 sky130_fd_sc_hd__a22o_1 \U$$2296  (.A1(net1688),
    .A2(net574),
    .B1(net1681),
    .B2(net847),
    .X(\t$5578 ));
 sky130_fd_sc_hd__xor2_1 \U$$2297  (.A(\t$5578 ),
    .B(net1435),
    .X(booth_b32_m49));
 sky130_fd_sc_hd__a22o_1 \U$$2298  (.A1(net1680),
    .A2(net573),
    .B1(net1655),
    .B2(net846),
    .X(\t$5579 ));
 sky130_fd_sc_hd__xor2_1 \U$$2299  (.A(\t$5579 ),
    .B(net1434),
    .X(booth_b32_m50));
 sky130_fd_sc_hd__xor2_1 \U$$23  (.A(\t$4418 ),
    .B(net1573),
    .X(booth_b0_m8));
 sky130_fd_sc_hd__xor2_1 \U$$230  (.A(\t$4522 ),
    .B(net1388),
    .X(booth_b2_m43));
 sky130_fd_sc_hd__a22o_1 \U$$2300  (.A1(net1655),
    .A2(net573),
    .B1(net1647),
    .B2(net846),
    .X(\t$5580 ));
 sky130_fd_sc_hd__xor2_1 \U$$2301  (.A(\t$5580 ),
    .B(net1434),
    .X(booth_b32_m51));
 sky130_fd_sc_hd__a22o_1 \U$$2302  (.A1(net1647),
    .A2(net574),
    .B1(net1639),
    .B2(net847),
    .X(\t$5581 ));
 sky130_fd_sc_hd__xor2_1 \U$$2303  (.A(\t$5581 ),
    .B(net1435),
    .X(booth_b32_m52));
 sky130_fd_sc_hd__a22o_1 \U$$2304  (.A1(net1639),
    .A2(net574),
    .B1(net1631),
    .B2(net847),
    .X(\t$5582 ));
 sky130_fd_sc_hd__xor2_1 \U$$2305  (.A(\t$5582 ),
    .B(net1436),
    .X(booth_b32_m53));
 sky130_fd_sc_hd__a22o_1 \U$$2306  (.A1(net1631),
    .A2(net574),
    .B1(net1622),
    .B2(net847),
    .X(\t$5583 ));
 sky130_fd_sc_hd__xor2_1 \U$$2307  (.A(\t$5583 ),
    .B(net1435),
    .X(booth_b32_m54));
 sky130_fd_sc_hd__a22o_1 \U$$2308  (.A1(net1622),
    .A2(net574),
    .B1(net1613),
    .B2(net847),
    .X(\t$5584 ));
 sky130_fd_sc_hd__xor2_1 \U$$2309  (.A(\t$5584 ),
    .B(net1435),
    .X(booth_b32_m55));
 sky130_fd_sc_hd__a22o_1 \U$$231  (.A1(net1729),
    .A2(net621),
    .B1(net1720),
    .B2(net894),
    .X(\t$4523 ));
 sky130_fd_sc_hd__a22o_1 \U$$2310  (.A1(net1613),
    .A2(net574),
    .B1(net1606),
    .B2(net847),
    .X(\t$5585 ));
 sky130_fd_sc_hd__xor2_1 \U$$2311  (.A(\t$5585 ),
    .B(net1434),
    .X(booth_b32_m56));
 sky130_fd_sc_hd__a22o_1 \U$$2312  (.A1(net1606),
    .A2(net574),
    .B1(net1598),
    .B2(net847),
    .X(\t$5586 ));
 sky130_fd_sc_hd__xor2_1 \U$$2313  (.A(\t$5586 ),
    .B(net1436),
    .X(booth_b32_m57));
 sky130_fd_sc_hd__a22o_1 \U$$2314  (.A1(net1596),
    .A2(net573),
    .B1(net1587),
    .B2(net846),
    .X(\t$5587 ));
 sky130_fd_sc_hd__xor2_1 \U$$2315  (.A(\t$5587 ),
    .B(net1436),
    .X(booth_b32_m58));
 sky130_fd_sc_hd__a22o_1 \U$$2316  (.A1(net1590),
    .A2(net575),
    .B1(net1582),
    .B2(net848),
    .X(\t$5588 ));
 sky130_fd_sc_hd__xor2_1 \U$$2317  (.A(\t$5588 ),
    .B(net1437),
    .X(booth_b32_m59));
 sky130_fd_sc_hd__a22o_1 \U$$2318  (.A1(net1584),
    .A2(net575),
    .B1(net1557),
    .B2(net848),
    .X(\t$5589 ));
 sky130_fd_sc_hd__xor2_1 \U$$2319  (.A(\t$5589 ),
    .B(net1437),
    .X(booth_b32_m60));
 sky130_fd_sc_hd__xor2_1 \U$$232  (.A(\t$4523 ),
    .B(net1386),
    .X(booth_b2_m44));
 sky130_fd_sc_hd__a22o_1 \U$$2320  (.A1(net1555),
    .A2(net575),
    .B1(net1547),
    .B2(net848),
    .X(\t$5590 ));
 sky130_fd_sc_hd__xor2_1 \U$$2321  (.A(\t$5590 ),
    .B(net1437),
    .X(booth_b32_m61));
 sky130_fd_sc_hd__a22o_1 \U$$2322  (.A1(net1547),
    .A2(net575),
    .B1(net1539),
    .B2(net848),
    .X(\t$5591 ));
 sky130_fd_sc_hd__xor2_1 \U$$2323  (.A(\t$5591 ),
    .B(net1437),
    .X(booth_b32_m62));
 sky130_fd_sc_hd__a22o_1 \U$$2324  (.A1(net1542),
    .A2(net575),
    .B1(net1534),
    .B2(net848),
    .X(\t$5592 ));
 sky130_fd_sc_hd__xor2_1 \U$$2325  (.A(\t$5592 ),
    .B(net1437),
    .X(booth_b32_m63));
 sky130_fd_sc_hd__a22o_1 \U$$2326  (.A1(net124),
    .A2(net575),
    .B1(net1774),
    .B2(net848),
    .X(\t$5593 ));
 sky130_fd_sc_hd__xor2_1 \U$$2327  (.A(\t$5593 ),
    .B(net1437),
    .X(booth_b32_m64));
 sky130_fd_sc_hd__inv_1 \U$$2328  (.A(net1437),
    .Y(\notsign$5594 ));
 sky130_fd_sc_hd__inv_1 \U$$2329  (.A(net1435),
    .Y(\notblock$5595[0] ));
 sky130_fd_sc_hd__a22o_1 \U$$233  (.A1(net1720),
    .A2(net621),
    .B1(net1711),
    .B2(net894),
    .X(\t$4524 ));
 sky130_fd_sc_hd__inv_1 \U$$2330  (.A(net28),
    .Y(\notblock$5595[1] ));
 sky130_fd_sc_hd__inv_1 \U$$2331  (.A(net1426),
    .Y(\notblock$5595[2] ));
 sky130_fd_sc_hd__and2_1 \U$$2332  (.A(net1426),
    .B(\notblock$5595[1] ),
    .X(\t$5596 ));
 sky130_fd_sc_hd__a32o_1 \U$$2333  (.A1(\notblock$5595[2] ),
    .A2(net28),
    .A3(net1435),
    .B1(\t$5596 ),
    .B2(\notblock$5595[0] ),
    .X(\sel_0$5597 ));
 sky130_fd_sc_hd__xor2_2 \U$$2334  (.A(net28),
    .B(net1435),
    .X(\sel_1$5598 ));
 sky130_fd_sc_hd__a22o_1 \U$$2335  (.A1(net1775),
    .A2(net563),
    .B1(net1230),
    .B2(net836),
    .X(\t$5599 ));
 sky130_fd_sc_hd__xor2_1 \U$$2336  (.A(\t$5599 ),
    .B(net1423),
    .X(booth_b34_m0));
 sky130_fd_sc_hd__a22o_1 \U$$2337  (.A1(net1232),
    .A2(net563),
    .B1(net1126),
    .B2(net836),
    .X(\t$5600 ));
 sky130_fd_sc_hd__xor2_1 \U$$2338  (.A(\t$5600 ),
    .B(net1423),
    .X(booth_b34_m1));
 sky130_fd_sc_hd__a22o_1 \U$$2339  (.A1(net1126),
    .A2(net563),
    .B1(net1036),
    .B2(net836),
    .X(\t$5601 ));
 sky130_fd_sc_hd__xor2_1 \U$$234  (.A(\t$4524 ),
    .B(net1387),
    .X(booth_b2_m45));
 sky130_fd_sc_hd__xor2_1 \U$$2340  (.A(\t$5601 ),
    .B(net1423),
    .X(booth_b34_m2));
 sky130_fd_sc_hd__a22o_1 \U$$2341  (.A1(net1036),
    .A2(net563),
    .B1(net936),
    .B2(net836),
    .X(\t$5602 ));
 sky130_fd_sc_hd__xor2_1 \U$$2342  (.A(\t$5602 ),
    .B(net1423),
    .X(booth_b34_m3));
 sky130_fd_sc_hd__a22o_1 \U$$2343  (.A1(net932),
    .A2(net560),
    .B1(net1671),
    .B2(net833),
    .X(\t$5603 ));
 sky130_fd_sc_hd__xor2_1 \U$$2344  (.A(\t$5603 ),
    .B(net1420),
    .X(booth_b34_m4));
 sky130_fd_sc_hd__a22o_1 \U$$2345  (.A1(net1672),
    .A2(net561),
    .B1(net1561),
    .B2(net834),
    .X(\t$5604 ));
 sky130_fd_sc_hd__xor2_1 \U$$2346  (.A(\t$5604 ),
    .B(net1420),
    .X(booth_b34_m5));
 sky130_fd_sc_hd__a22o_1 \U$$2347  (.A1(net1561),
    .A2(net561),
    .B1(net1521),
    .B2(net834),
    .X(\t$5605 ));
 sky130_fd_sc_hd__xor2_1 \U$$2348  (.A(\t$5605 ),
    .B(net1421),
    .X(booth_b34_m6));
 sky130_fd_sc_hd__a22o_1 \U$$2349  (.A1(net1519),
    .A2(net560),
    .B1(net1511),
    .B2(net833),
    .X(\t$5606 ));
 sky130_fd_sc_hd__a22o_1 \U$$235  (.A1(net1711),
    .A2(net621),
    .B1(net1703),
    .B2(net894),
    .X(\t$4525 ));
 sky130_fd_sc_hd__xor2_1 \U$$2350  (.A(\t$5606 ),
    .B(net1420),
    .X(booth_b34_m7));
 sky130_fd_sc_hd__a22o_1 \U$$2351  (.A1(net1512),
    .A2(net560),
    .B1(net1504),
    .B2(net833),
    .X(\t$5607 ));
 sky130_fd_sc_hd__xor2_1 \U$$2352  (.A(\t$5607 ),
    .B(net1420),
    .X(booth_b34_m8));
 sky130_fd_sc_hd__a22o_1 \U$$2353  (.A1(net1504),
    .A2(net560),
    .B1(net1495),
    .B2(net833),
    .X(\t$5608 ));
 sky130_fd_sc_hd__xor2_1 \U$$2354  (.A(\t$5608 ),
    .B(net1420),
    .X(booth_b34_m9));
 sky130_fd_sc_hd__a22o_1 \U$$2355  (.A1(net1494),
    .A2(net560),
    .B1(net1219),
    .B2(net833),
    .X(\t$5609 ));
 sky130_fd_sc_hd__xor2_1 \U$$2356  (.A(\t$5609 ),
    .B(net1420),
    .X(booth_b34_m10));
 sky130_fd_sc_hd__a22o_1 \U$$2357  (.A1(net1220),
    .A2(net560),
    .B1(net1213),
    .B2(net833),
    .X(\t$5610 ));
 sky130_fd_sc_hd__xor2_1 \U$$2358  (.A(\t$5610 ),
    .B(net1420),
    .X(booth_b34_m11));
 sky130_fd_sc_hd__a22o_1 \U$$2359  (.A1(net1213),
    .A2(net560),
    .B1(net1202),
    .B2(net833),
    .X(\t$5611 ));
 sky130_fd_sc_hd__xor2_1 \U$$236  (.A(\t$4525 ),
    .B(net1387),
    .X(booth_b2_m46));
 sky130_fd_sc_hd__xor2_1 \U$$2360  (.A(\t$5611 ),
    .B(net1420),
    .X(booth_b34_m12));
 sky130_fd_sc_hd__a22o_1 \U$$2361  (.A1(net1202),
    .A2(net560),
    .B1(net1193),
    .B2(net833),
    .X(\t$5612 ));
 sky130_fd_sc_hd__xor2_1 \U$$2362  (.A(\t$5612 ),
    .B(net1420),
    .X(booth_b34_m13));
 sky130_fd_sc_hd__a22o_1 \U$$2363  (.A1(net1193),
    .A2(net560),
    .B1(net1174),
    .B2(net833),
    .X(\t$5613 ));
 sky130_fd_sc_hd__xor2_1 \U$$2364  (.A(\t$5613 ),
    .B(net1420),
    .X(booth_b34_m14));
 sky130_fd_sc_hd__a22o_1 \U$$2365  (.A1(net1176),
    .A2(net561),
    .B1(net1167),
    .B2(net834),
    .X(\t$5614 ));
 sky130_fd_sc_hd__xor2_1 \U$$2366  (.A(\t$5614 ),
    .B(net1421),
    .X(booth_b34_m15));
 sky130_fd_sc_hd__a22o_1 \U$$2367  (.A1(net1170),
    .A2(net563),
    .B1(net1161),
    .B2(net836),
    .X(\t$5615 ));
 sky130_fd_sc_hd__xor2_1 \U$$2368  (.A(\t$5615 ),
    .B(net1423),
    .X(booth_b34_m16));
 sky130_fd_sc_hd__a22o_1 \U$$2369  (.A1(net1162),
    .A2(net563),
    .B1(net1150),
    .B2(net836),
    .X(\t$5616 ));
 sky130_fd_sc_hd__a22o_1 \U$$237  (.A1(net1706),
    .A2(net626),
    .B1(net1698),
    .B2(net899),
    .X(\t$4526 ));
 sky130_fd_sc_hd__xor2_1 \U$$2370  (.A(\t$5616 ),
    .B(net1423),
    .X(booth_b34_m17));
 sky130_fd_sc_hd__a22o_1 \U$$2371  (.A1(net1150),
    .A2(net563),
    .B1(net1144),
    .B2(net836),
    .X(\t$5617 ));
 sky130_fd_sc_hd__xor2_1 \U$$2372  (.A(\t$5617 ),
    .B(net1423),
    .X(booth_b34_m18));
 sky130_fd_sc_hd__a22o_1 \U$$2373  (.A1(net1144),
    .A2(net563),
    .B1(net1134),
    .B2(net836),
    .X(\t$5618 ));
 sky130_fd_sc_hd__xor2_1 \U$$2374  (.A(\t$5618 ),
    .B(net1423),
    .X(booth_b34_m19));
 sky130_fd_sc_hd__a22o_1 \U$$2375  (.A1(net1134),
    .A2(net564),
    .B1(net1118),
    .B2(net837),
    .X(\t$5619 ));
 sky130_fd_sc_hd__xor2_1 \U$$2376  (.A(\t$5619 ),
    .B(net1423),
    .X(booth_b34_m20));
 sky130_fd_sc_hd__a22o_1 \U$$2377  (.A1(net1118),
    .A2(net563),
    .B1(net1109),
    .B2(net836),
    .X(\t$5620 ));
 sky130_fd_sc_hd__xor2_1 \U$$2378  (.A(\t$5620 ),
    .B(net1424),
    .X(booth_b34_m21));
 sky130_fd_sc_hd__a22o_1 \U$$2379  (.A1(net1109),
    .A2(net564),
    .B1(net1101),
    .B2(net837),
    .X(\t$5621 ));
 sky130_fd_sc_hd__xor2_1 \U$$238  (.A(\t$4526 ),
    .B(net1392),
    .X(booth_b2_m47));
 sky130_fd_sc_hd__xor2_1 \U$$2380  (.A(\t$5621 ),
    .B(net1424),
    .X(booth_b34_m22));
 sky130_fd_sc_hd__a22o_1 \U$$2381  (.A1(net1100),
    .A2(net560),
    .B1(net1091),
    .B2(net833),
    .X(\t$5622 ));
 sky130_fd_sc_hd__xor2_1 \U$$2382  (.A(\t$5622 ),
    .B(net1421),
    .X(booth_b34_m23));
 sky130_fd_sc_hd__a22o_1 \U$$2383  (.A1(net1092),
    .A2(net563),
    .B1(net1084),
    .B2(net836),
    .X(\t$5623 ));
 sky130_fd_sc_hd__xor2_1 \U$$2384  (.A(\t$5623 ),
    .B(net1421),
    .X(booth_b34_m24));
 sky130_fd_sc_hd__a22o_1 \U$$2385  (.A1(net1082),
    .A2(net561),
    .B1(net1073),
    .B2(net834),
    .X(\t$5624 ));
 sky130_fd_sc_hd__xor2_1 \U$$2386  (.A(\t$5624 ),
    .B(net1421),
    .X(booth_b34_m25));
 sky130_fd_sc_hd__a22o_1 \U$$2387  (.A1(net1073),
    .A2(net561),
    .B1(net1065),
    .B2(net834),
    .X(\t$5625 ));
 sky130_fd_sc_hd__xor2_1 \U$$2388  (.A(\t$5625 ),
    .B(net1421),
    .X(booth_b34_m26));
 sky130_fd_sc_hd__a22o_1 \U$$2389  (.A1(net1065),
    .A2(net562),
    .B1(net1059),
    .B2(net835),
    .X(\t$5626 ));
 sky130_fd_sc_hd__a22o_1 \U$$239  (.A1(net1695),
    .A2(net621),
    .B1(net1687),
    .B2(net894),
    .X(\t$4527 ));
 sky130_fd_sc_hd__xor2_1 \U$$2390  (.A(\t$5626 ),
    .B(net1422),
    .X(booth_b34_m27));
 sky130_fd_sc_hd__a22o_1 \U$$2391  (.A1(net1062),
    .A2(net565),
    .B1(net1053),
    .B2(net838),
    .X(\t$5627 ));
 sky130_fd_sc_hd__xor2_1 \U$$2392  (.A(\t$5627 ),
    .B(net1425),
    .X(booth_b34_m28));
 sky130_fd_sc_hd__a22o_1 \U$$2393  (.A1(net1051),
    .A2(net562),
    .B1(net1043),
    .B2(net835),
    .X(\t$5628 ));
 sky130_fd_sc_hd__xor2_1 \U$$2394  (.A(\t$5628 ),
    .B(net1422),
    .X(booth_b34_m29));
 sky130_fd_sc_hd__a22o_1 \U$$2395  (.A1(net1042),
    .A2(net562),
    .B1(net1026),
    .B2(net835),
    .X(\t$5629 ));
 sky130_fd_sc_hd__xor2_1 \U$$2396  (.A(\t$5629 ),
    .B(net1422),
    .X(booth_b34_m30));
 sky130_fd_sc_hd__a22o_1 \U$$2397  (.A1(net1026),
    .A2(net564),
    .B1(net1018),
    .B2(net837),
    .X(\t$5630 ));
 sky130_fd_sc_hd__xor2_1 \U$$2398  (.A(\t$5630 ),
    .B(net1424),
    .X(booth_b34_m31));
 sky130_fd_sc_hd__a22o_1 \U$$2399  (.A1(net1018),
    .A2(net564),
    .B1(net1001),
    .B2(net837),
    .X(\t$5631 ));
 sky130_fd_sc_hd__a22o_1 \U$$24  (.A1(net1508),
    .A2(net446),
    .B1(net1499),
    .B2(net688),
    .X(\t$4419 ));
 sky130_fd_sc_hd__xor2_1 \U$$240  (.A(\t$4527 ),
    .B(net1387),
    .X(booth_b2_m48));
 sky130_fd_sc_hd__xor2_1 \U$$2400  (.A(\t$5631 ),
    .B(net1424),
    .X(booth_b34_m32));
 sky130_fd_sc_hd__a22o_1 \U$$2401  (.A1(net1001),
    .A2(net564),
    .B1(net993),
    .B2(net837),
    .X(\t$5632 ));
 sky130_fd_sc_hd__xor2_1 \U$$2402  (.A(\t$5632 ),
    .B(net1424),
    .X(booth_b34_m33));
 sky130_fd_sc_hd__a22o_1 \U$$2403  (.A1(net996),
    .A2(net567),
    .B1(net988),
    .B2(net840),
    .X(\t$5633 ));
 sky130_fd_sc_hd__xor2_1 \U$$2404  (.A(\t$5633 ),
    .B(net1428),
    .X(booth_b34_m34));
 sky130_fd_sc_hd__a22o_1 \U$$2405  (.A1(net988),
    .A2(net567),
    .B1(net979),
    .B2(net840),
    .X(\t$5634 ));
 sky130_fd_sc_hd__xor2_1 \U$$2406  (.A(\t$5634 ),
    .B(net1428),
    .X(booth_b34_m35));
 sky130_fd_sc_hd__a22o_1 \U$$2407  (.A1(net975),
    .A2(net565),
    .B1(net966),
    .B2(net838),
    .X(\t$5635 ));
 sky130_fd_sc_hd__xor2_1 \U$$2408  (.A(\t$5635 ),
    .B(net1425),
    .X(booth_b34_m36));
 sky130_fd_sc_hd__a22o_1 \U$$2409  (.A1(net967),
    .A2(net565),
    .B1(net958),
    .B2(net838),
    .X(\t$5636 ));
 sky130_fd_sc_hd__a22o_1 \U$$241  (.A1(net1691),
    .A2(net626),
    .B1(net1683),
    .B2(net899),
    .X(\t$4528 ));
 sky130_fd_sc_hd__xor2_1 \U$$2410  (.A(\t$5636 ),
    .B(net1425),
    .X(booth_b34_m37));
 sky130_fd_sc_hd__a22o_1 \U$$2411  (.A1(net958),
    .A2(net562),
    .B1(net949),
    .B2(net835),
    .X(\t$5637 ));
 sky130_fd_sc_hd__xor2_1 \U$$2412  (.A(\t$5637 ),
    .B(net1422),
    .X(booth_b34_m38));
 sky130_fd_sc_hd__a22o_1 \U$$2413  (.A1(net949),
    .A2(net562),
    .B1(net941),
    .B2(net835),
    .X(\t$5638 ));
 sky130_fd_sc_hd__xor2_1 \U$$2414  (.A(\t$5638 ),
    .B(net1422),
    .X(booth_b34_m39));
 sky130_fd_sc_hd__a22o_1 \U$$2415  (.A1(net941),
    .A2(net562),
    .B1(net925),
    .B2(net835),
    .X(\t$5639 ));
 sky130_fd_sc_hd__xor2_1 \U$$2416  (.A(\t$5639 ),
    .B(net1422),
    .X(booth_b34_m40));
 sky130_fd_sc_hd__a22o_1 \U$$2417  (.A1(net926),
    .A2(net565),
    .B1(net1747),
    .B2(net838),
    .X(\t$5640 ));
 sky130_fd_sc_hd__xor2_1 \U$$2418  (.A(\t$5640 ),
    .B(net1425),
    .X(booth_b34_m41));
 sky130_fd_sc_hd__a22o_1 \U$$2419  (.A1(net1747),
    .A2(net565),
    .B1(net1739),
    .B2(net838),
    .X(\t$5641 ));
 sky130_fd_sc_hd__xor2_1 \U$$242  (.A(\t$4528 ),
    .B(net1392),
    .X(booth_b2_m49));
 sky130_fd_sc_hd__xor2_1 \U$$2420  (.A(\t$5641 ),
    .B(net1425),
    .X(booth_b34_m42));
 sky130_fd_sc_hd__a22o_1 \U$$2421  (.A1(net1738),
    .A2(net565),
    .B1(net1730),
    .B2(net838),
    .X(\t$5642 ));
 sky130_fd_sc_hd__xor2_1 \U$$2422  (.A(\t$5642 ),
    .B(net1425),
    .X(booth_b34_m43));
 sky130_fd_sc_hd__a22o_1 \U$$2423  (.A1(net1731),
    .A2(net566),
    .B1(net1722),
    .B2(net839),
    .X(\t$5643 ));
 sky130_fd_sc_hd__xor2_1 \U$$2424  (.A(\t$5643 ),
    .B(net1426),
    .X(booth_b34_m44));
 sky130_fd_sc_hd__a22o_1 \U$$2425  (.A1(net1722),
    .A2(net565),
    .B1(net1713),
    .B2(net838),
    .X(\t$5644 ));
 sky130_fd_sc_hd__xor2_1 \U$$2426  (.A(\t$5644 ),
    .B(net1425),
    .X(booth_b34_m45));
 sky130_fd_sc_hd__a22o_1 \U$$2427  (.A1(net1713),
    .A2(net565),
    .B1(net1704),
    .B2(net838),
    .X(\t$5645 ));
 sky130_fd_sc_hd__xor2_1 \U$$2428  (.A(\t$5645 ),
    .B(net1425),
    .X(booth_b34_m46));
 sky130_fd_sc_hd__a22o_1 \U$$2429  (.A1(net1705),
    .A2(net566),
    .B1(net1697),
    .B2(net839),
    .X(\t$5646 ));
 sky130_fd_sc_hd__a22o_1 \U$$243  (.A1(net1683),
    .A2(net626),
    .B1(net1658),
    .B2(net899),
    .X(\t$4529 ));
 sky130_fd_sc_hd__xor2_1 \U$$2430  (.A(\t$5646 ),
    .B(net1426),
    .X(booth_b34_m47));
 sky130_fd_sc_hd__a22o_1 \U$$2431  (.A1(net1696),
    .A2(net566),
    .B1(net1688),
    .B2(net839),
    .X(\t$5647 ));
 sky130_fd_sc_hd__xor2_1 \U$$2432  (.A(\t$5647 ),
    .B(net1426),
    .X(booth_b34_m48));
 sky130_fd_sc_hd__a22o_1 \U$$2433  (.A1(net1688),
    .A2(net565),
    .B1(net1680),
    .B2(net838),
    .X(\t$5648 ));
 sky130_fd_sc_hd__xor2_1 \U$$2434  (.A(\t$5648 ),
    .B(net1425),
    .X(booth_b34_m49));
 sky130_fd_sc_hd__a22o_1 \U$$2435  (.A1(net1680),
    .A2(net566),
    .B1(net1655),
    .B2(net839),
    .X(\t$5649 ));
 sky130_fd_sc_hd__xor2_1 \U$$2436  (.A(\t$5649 ),
    .B(net1426),
    .X(booth_b34_m50));
 sky130_fd_sc_hd__a22o_1 \U$$2437  (.A1(net1656),
    .A2(net566),
    .B1(net1648),
    .B2(net839),
    .X(\t$5650 ));
 sky130_fd_sc_hd__xor2_1 \U$$2438  (.A(\t$5650 ),
    .B(net1427),
    .X(booth_b34_m51));
 sky130_fd_sc_hd__a22o_1 \U$$2439  (.A1(net1647),
    .A2(net566),
    .B1(net1639),
    .B2(net839),
    .X(\t$5651 ));
 sky130_fd_sc_hd__xor2_1 \U$$244  (.A(\t$4529 ),
    .B(net1392),
    .X(booth_b2_m50));
 sky130_fd_sc_hd__xor2_1 \U$$2440  (.A(\t$5651 ),
    .B(net1426),
    .X(booth_b34_m52));
 sky130_fd_sc_hd__a22o_1 \U$$2441  (.A1(net1639),
    .A2(net566),
    .B1(net1631),
    .B2(net839),
    .X(\t$5652 ));
 sky130_fd_sc_hd__xor2_1 \U$$2442  (.A(\t$5652 ),
    .B(net1426),
    .X(booth_b34_m53));
 sky130_fd_sc_hd__a22o_1 \U$$2443  (.A1(net1632),
    .A2(net566),
    .B1(net1622),
    .B2(net839),
    .X(\t$5653 ));
 sky130_fd_sc_hd__xor2_1 \U$$2444  (.A(\t$5653 ),
    .B(net1427),
    .X(booth_b34_m54));
 sky130_fd_sc_hd__a22o_1 \U$$2445  (.A1(net1628),
    .A2(net565),
    .B1(net1614),
    .B2(net838),
    .X(\t$5654 ));
 sky130_fd_sc_hd__xor2_1 \U$$2446  (.A(\t$5654 ),
    .B(net1425),
    .X(booth_b34_m55));
 sky130_fd_sc_hd__a22o_1 \U$$2447  (.A1(net1615),
    .A2(net567),
    .B1(net1607),
    .B2(net840),
    .X(\t$5655 ));
 sky130_fd_sc_hd__xor2_1 \U$$2448  (.A(\t$5655 ),
    .B(net1427),
    .X(booth_b34_m56));
 sky130_fd_sc_hd__a22o_1 \U$$2449  (.A1(net1608),
    .A2(net567),
    .B1(net1600),
    .B2(net840),
    .X(\t$5656 ));
 sky130_fd_sc_hd__a22o_1 \U$$245  (.A1(net1658),
    .A2(net626),
    .B1(net1650),
    .B2(net899),
    .X(\t$4530 ));
 sky130_fd_sc_hd__xor2_1 \U$$2450  (.A(\t$5656 ),
    .B(net1428),
    .X(booth_b34_m57));
 sky130_fd_sc_hd__a22o_1 \U$$2451  (.A1(net1602),
    .A2(net567),
    .B1(net1592),
    .B2(net840),
    .X(\t$5657 ));
 sky130_fd_sc_hd__xor2_1 \U$$2452  (.A(\t$5657 ),
    .B(net1428),
    .X(booth_b34_m58));
 sky130_fd_sc_hd__a22o_1 \U$$2453  (.A1(net1590),
    .A2(net567),
    .B1(net1582),
    .B2(net840),
    .X(\t$5658 ));
 sky130_fd_sc_hd__xor2_1 \U$$2454  (.A(\t$5658 ),
    .B(net1428),
    .X(booth_b34_m59));
 sky130_fd_sc_hd__a22o_1 \U$$2455  (.A1(net1582),
    .A2(net567),
    .B1(net1555),
    .B2(net840),
    .X(\t$5659 ));
 sky130_fd_sc_hd__xor2_1 \U$$2456  (.A(\t$5659 ),
    .B(net1428),
    .X(booth_b34_m60));
 sky130_fd_sc_hd__a22o_1 \U$$2457  (.A1(net1557),
    .A2(net568),
    .B1(net1550),
    .B2(net841),
    .X(\t$5660 ));
 sky130_fd_sc_hd__xor2_1 \U$$2458  (.A(\t$5660 ),
    .B(net1428),
    .X(booth_b34_m61));
 sky130_fd_sc_hd__a22o_1 \U$$2459  (.A1(net1547),
    .A2(net567),
    .B1(net123),
    .B2(net840),
    .X(\t$5661 ));
 sky130_fd_sc_hd__xor2_1 \U$$246  (.A(\t$4530 ),
    .B(net1392),
    .X(booth_b2_m51));
 sky130_fd_sc_hd__xor2_1 \U$$2460  (.A(\t$5661 ),
    .B(net1428),
    .X(booth_b34_m62));
 sky130_fd_sc_hd__a22o_1 \U$$2461  (.A1(net1542),
    .A2(net567),
    .B1(net1534),
    .B2(net840),
    .X(\t$5662 ));
 sky130_fd_sc_hd__xor2_1 \U$$2462  (.A(\t$5662 ),
    .B(net1428),
    .X(booth_b34_m63));
 sky130_fd_sc_hd__a22o_1 \U$$2463  (.A1(net1534),
    .A2(net567),
    .B1(net1776),
    .B2(net840),
    .X(\t$5663 ));
 sky130_fd_sc_hd__xor2_1 \U$$2464  (.A(\t$5663 ),
    .B(net1428),
    .X(booth_b34_m64));
 sky130_fd_sc_hd__inv_1 \U$$2465  (.A(net1429),
    .Y(\notsign$5664 ));
 sky130_fd_sc_hd__inv_1 \U$$2466  (.A(net1426),
    .Y(\notblock$5665[0] ));
 sky130_fd_sc_hd__inv_1 \U$$2467  (.A(net30),
    .Y(\notblock$5665[1] ));
 sky130_fd_sc_hd__inv_1 \U$$2468  (.A(net1408),
    .Y(\notblock$5665[2] ));
 sky130_fd_sc_hd__and2_1 \U$$2469  (.A(net1408),
    .B(\notblock$5665[1] ),
    .X(\t$5666 ));
 sky130_fd_sc_hd__a22o_1 \U$$247  (.A1(net1650),
    .A2(net626),
    .B1(net1642),
    .B2(net899),
    .X(\t$4531 ));
 sky130_fd_sc_hd__a32o_1 \U$$2470  (.A1(\notblock$5665[2] ),
    .A2(net30),
    .A3(net1426),
    .B1(\t$5666 ),
    .B2(\notblock$5665[0] ),
    .X(\sel_0$5667 ));
 sky130_fd_sc_hd__xor2_1 \U$$2471  (.A(net30),
    .B(net1427),
    .X(\sel_1$5668 ));
 sky130_fd_sc_hd__a22o_1 \U$$2472  (.A1(net1777),
    .A2(net554),
    .B1(net1232),
    .B2(net827),
    .X(\t$5669 ));
 sky130_fd_sc_hd__xor2_1 \U$$2473  (.A(\t$5669 ),
    .B(net1406),
    .X(booth_b36_m0));
 sky130_fd_sc_hd__a22o_1 \U$$2474  (.A1(net1232),
    .A2(net552),
    .B1(net1128),
    .B2(net825),
    .X(\t$5670 ));
 sky130_fd_sc_hd__xor2_1 \U$$2475  (.A(\t$5670 ),
    .B(net1403),
    .X(booth_b36_m1));
 sky130_fd_sc_hd__a22o_1 \U$$2476  (.A1(net1122),
    .A2(net551),
    .B1(net1031),
    .B2(net824),
    .X(\t$5671 ));
 sky130_fd_sc_hd__xor2_1 \U$$2477  (.A(\t$5671 ),
    .B(net1403),
    .X(booth_b36_m2));
 sky130_fd_sc_hd__a22o_1 \U$$2478  (.A1(net1032),
    .A2(net551),
    .B1(net933),
    .B2(net824),
    .X(\t$5672 ));
 sky130_fd_sc_hd__xor2_1 \U$$2479  (.A(\t$5672 ),
    .B(net1404),
    .X(booth_b36_m3));
 sky130_fd_sc_hd__xor2_1 \U$$248  (.A(\t$4531 ),
    .B(net1392),
    .X(booth_b2_m52));
 sky130_fd_sc_hd__a22o_1 \U$$2480  (.A1(net933),
    .A2(net552),
    .B1(net1672),
    .B2(net825),
    .X(\t$5673 ));
 sky130_fd_sc_hd__xor2_1 \U$$2481  (.A(\t$5673 ),
    .B(net1404),
    .X(booth_b36_m4));
 sky130_fd_sc_hd__a22o_1 \U$$2482  (.A1(net1671),
    .A2(net551),
    .B1(net1560),
    .B2(net824),
    .X(\t$5674 ));
 sky130_fd_sc_hd__xor2_1 \U$$2483  (.A(\t$5674 ),
    .B(net1403),
    .X(booth_b36_m5));
 sky130_fd_sc_hd__a22o_1 \U$$2484  (.A1(net1560),
    .A2(net551),
    .B1(net1520),
    .B2(net824),
    .X(\t$5675 ));
 sky130_fd_sc_hd__xor2_1 \U$$2485  (.A(\t$5675 ),
    .B(net1403),
    .X(booth_b36_m6));
 sky130_fd_sc_hd__a22o_1 \U$$2486  (.A1(net1520),
    .A2(net551),
    .B1(net1512),
    .B2(net824),
    .X(\t$5676 ));
 sky130_fd_sc_hd__xor2_1 \U$$2487  (.A(\t$5676 ),
    .B(net1403),
    .X(booth_b36_m7));
 sky130_fd_sc_hd__a22o_1 \U$$2488  (.A1(net1511),
    .A2(net551),
    .B1(net1503),
    .B2(net824),
    .X(\t$5677 ));
 sky130_fd_sc_hd__xor2_1 \U$$2489  (.A(\t$5677 ),
    .B(net1403),
    .X(booth_b36_m8));
 sky130_fd_sc_hd__a22o_1 \U$$249  (.A1(net1642),
    .A2(net626),
    .B1(net1637),
    .B2(net899),
    .X(\t$4532 ));
 sky130_fd_sc_hd__a22o_1 \U$$2490  (.A1(net1504),
    .A2(net551),
    .B1(net1497),
    .B2(net824),
    .X(\t$5678 ));
 sky130_fd_sc_hd__xor2_1 \U$$2491  (.A(\t$5678 ),
    .B(net1403),
    .X(booth_b36_m9));
 sky130_fd_sc_hd__a22o_1 \U$$2492  (.A1(net1497),
    .A2(net551),
    .B1(net1223),
    .B2(net824),
    .X(\t$5679 ));
 sky130_fd_sc_hd__xor2_1 \U$$2493  (.A(\t$5679 ),
    .B(net1403),
    .X(booth_b36_m10));
 sky130_fd_sc_hd__a22o_1 \U$$2494  (.A1(net1220),
    .A2(net551),
    .B1(net1213),
    .B2(net824),
    .X(\t$5680 ));
 sky130_fd_sc_hd__xor2_1 \U$$2495  (.A(\t$5680 ),
    .B(net1403),
    .X(booth_b36_m11));
 sky130_fd_sc_hd__a22o_1 \U$$2496  (.A1(net1213),
    .A2(net551),
    .B1(net1202),
    .B2(net824),
    .X(\t$5681 ));
 sky130_fd_sc_hd__xor2_1 \U$$2497  (.A(\t$5681 ),
    .B(net1403),
    .X(booth_b36_m12));
 sky130_fd_sc_hd__a22o_1 \U$$2498  (.A1(net1204),
    .A2(net552),
    .B1(net1195),
    .B2(net825),
    .X(\t$5682 ));
 sky130_fd_sc_hd__xor2_1 \U$$2499  (.A(\t$5682 ),
    .B(net1404),
    .X(booth_b36_m13));
 sky130_fd_sc_hd__xor2_1 \U$$25  (.A(\t$4419 ),
    .B(net1573),
    .X(booth_b0_m9));
 sky130_fd_sc_hd__xor2_1 \U$$250  (.A(\t$4532 ),
    .B(net1392),
    .X(booth_b2_m53));
 sky130_fd_sc_hd__a22o_1 \U$$2500  (.A1(net1198),
    .A2(net554),
    .B1(net1180),
    .B2(net827),
    .X(\t$5683 ));
 sky130_fd_sc_hd__xor2_1 \U$$2501  (.A(\t$5683 ),
    .B(net1406),
    .X(booth_b36_m14));
 sky130_fd_sc_hd__a22o_1 \U$$2502  (.A1(net1180),
    .A2(net554),
    .B1(net1171),
    .B2(net827),
    .X(\t$5684 ));
 sky130_fd_sc_hd__xor2_1 \U$$2503  (.A(\t$5684 ),
    .B(net1406),
    .X(booth_b36_m15));
 sky130_fd_sc_hd__a22o_1 \U$$2504  (.A1(net1171),
    .A2(net554),
    .B1(net1162),
    .B2(net827),
    .X(\t$5685 ));
 sky130_fd_sc_hd__xor2_1 \U$$2505  (.A(\t$5685 ),
    .B(net1406),
    .X(booth_b36_m16));
 sky130_fd_sc_hd__a22o_1 \U$$2506  (.A1(net1162),
    .A2(net554),
    .B1(net1150),
    .B2(net827),
    .X(\t$5686 ));
 sky130_fd_sc_hd__xor2_1 \U$$2507  (.A(\t$5686 ),
    .B(net1406),
    .X(booth_b36_m17));
 sky130_fd_sc_hd__a22o_1 \U$$2508  (.A1(net1149),
    .A2(net554),
    .B1(net1144),
    .B2(net827),
    .X(\t$5687 ));
 sky130_fd_sc_hd__xor2_1 \U$$2509  (.A(\t$5687 ),
    .B(net1406),
    .X(booth_b36_m18));
 sky130_fd_sc_hd__a22o_1 \U$$251  (.A1(net1633),
    .A2(\sel_0$4477 ),
    .B1(net1623),
    .B2(\sel_1$4478 ),
    .X(\t$4533 ));
 sky130_fd_sc_hd__a22o_1 \U$$2510  (.A1(net1144),
    .A2(net554),
    .B1(net1134),
    .B2(net827),
    .X(\t$5688 ));
 sky130_fd_sc_hd__xor2_1 \U$$2511  (.A(\t$5688 ),
    .B(net1406),
    .X(booth_b36_m19));
 sky130_fd_sc_hd__a22o_1 \U$$2512  (.A1(net1134),
    .A2(net554),
    .B1(net1118),
    .B2(net827),
    .X(\t$5689 ));
 sky130_fd_sc_hd__xor2_1 \U$$2513  (.A(\t$5689 ),
    .B(net1406),
    .X(booth_b36_m20));
 sky130_fd_sc_hd__a22o_1 \U$$2514  (.A1(net1118),
    .A2(net552),
    .B1(net1109),
    .B2(net825),
    .X(\t$5690 ));
 sky130_fd_sc_hd__xor2_1 \U$$2515  (.A(\t$5690 ),
    .B(net1404),
    .X(booth_b36_m21));
 sky130_fd_sc_hd__a22o_1 \U$$2516  (.A1(net1109),
    .A2(net552),
    .B1(net1101),
    .B2(net825),
    .X(\t$5691 ));
 sky130_fd_sc_hd__xor2_1 \U$$2517  (.A(\t$5691 ),
    .B(net1404),
    .X(booth_b36_m22));
 sky130_fd_sc_hd__a22o_1 \U$$2518  (.A1(net1098),
    .A2(net552),
    .B1(net1090),
    .B2(net825),
    .X(\t$5692 ));
 sky130_fd_sc_hd__xor2_1 \U$$2519  (.A(\t$5692 ),
    .B(net1404),
    .X(booth_b36_m23));
 sky130_fd_sc_hd__xor2_1 \U$$252  (.A(\t$4533 ),
    .B(net1393),
    .X(booth_b2_m54));
 sky130_fd_sc_hd__a22o_1 \U$$2520  (.A1(net1090),
    .A2(net553),
    .B1(net1082),
    .B2(net826),
    .X(\t$5693 ));
 sky130_fd_sc_hd__xor2_1 \U$$2521  (.A(\t$5693 ),
    .B(net1405),
    .X(booth_b36_m24));
 sky130_fd_sc_hd__a22o_1 \U$$2522  (.A1(net1082),
    .A2(net553),
    .B1(net1079),
    .B2(net826),
    .X(\t$5694 ));
 sky130_fd_sc_hd__xor2_1 \U$$2523  (.A(\t$5694 ),
    .B(net1405),
    .X(booth_b36_m25));
 sky130_fd_sc_hd__a22o_1 \U$$2524  (.A1(net1078),
    .A2(net555),
    .B1(net1070),
    .B2(net828),
    .X(\t$5695 ));
 sky130_fd_sc_hd__xor2_1 \U$$2525  (.A(\t$5695 ),
    .B(net1405),
    .X(booth_b36_m26));
 sky130_fd_sc_hd__a22o_1 \U$$2526  (.A1(net1068),
    .A2(net553),
    .B1(net1060),
    .B2(net826),
    .X(\t$5696 ));
 sky130_fd_sc_hd__xor2_1 \U$$2527  (.A(\t$5696 ),
    .B(net1405),
    .X(booth_b36_m27));
 sky130_fd_sc_hd__a22o_1 \U$$2528  (.A1(net1058),
    .A2(net554),
    .B1(net1050),
    .B2(net827),
    .X(\t$5697 ));
 sky130_fd_sc_hd__xor2_1 \U$$2529  (.A(\t$5697 ),
    .B(net1406),
    .X(booth_b36_m28));
 sky130_fd_sc_hd__a22o_1 \U$$253  (.A1(net1623),
    .A2(net626),
    .B1(net1615),
    .B2(net899),
    .X(\t$4534 ));
 sky130_fd_sc_hd__a22o_1 \U$$2530  (.A1(net1050),
    .A2(net554),
    .B1(net1042),
    .B2(net827),
    .X(\t$5698 ));
 sky130_fd_sc_hd__xor2_1 \U$$2531  (.A(\t$5698 ),
    .B(net1407),
    .X(booth_b36_m29));
 sky130_fd_sc_hd__a22o_1 \U$$2532  (.A1(net1046),
    .A2(net559),
    .B1(net1030),
    .B2(net832),
    .X(\t$5699 ));
 sky130_fd_sc_hd__xor2_1 \U$$2533  (.A(\t$5699 ),
    .B(net1407),
    .X(booth_b36_m30));
 sky130_fd_sc_hd__a22o_1 \U$$2534  (.A1(net1029),
    .A2(net559),
    .B1(net1021),
    .B2(net832),
    .X(\t$5700 ));
 sky130_fd_sc_hd__xor2_1 \U$$2535  (.A(\t$5700 ),
    .B(net1407),
    .X(booth_b36_m31));
 sky130_fd_sc_hd__a22o_1 \U$$2536  (.A1(net1021),
    .A2(net557),
    .B1(net1004),
    .B2(net830),
    .X(\t$5701 ));
 sky130_fd_sc_hd__xor2_1 \U$$2537  (.A(\t$5701 ),
    .B(net1410),
    .X(booth_b36_m32));
 sky130_fd_sc_hd__a22o_1 \U$$2538  (.A1(net1004),
    .A2(net557),
    .B1(net996),
    .B2(net830),
    .X(\t$5702 ));
 sky130_fd_sc_hd__xor2_1 \U$$2539  (.A(\t$5702 ),
    .B(net1410),
    .X(booth_b36_m33));
 sky130_fd_sc_hd__xor2_1 \U$$254  (.A(\t$4534 ),
    .B(net1392),
    .X(booth_b2_m55));
 sky130_fd_sc_hd__a22o_1 \U$$2540  (.A1(net994),
    .A2(net555),
    .B1(net984),
    .B2(net828),
    .X(\t$5703 ));
 sky130_fd_sc_hd__xor2_1 \U$$2541  (.A(\t$5703 ),
    .B(net1409),
    .X(booth_b36_m34));
 sky130_fd_sc_hd__a22o_1 \U$$2542  (.A1(net984),
    .A2(net555),
    .B1(net975),
    .B2(net828),
    .X(\t$5704 ));
 sky130_fd_sc_hd__xor2_1 \U$$2543  (.A(\t$5704 ),
    .B(net1409),
    .X(booth_b36_m35));
 sky130_fd_sc_hd__a22o_1 \U$$2544  (.A1(net976),
    .A2(net556),
    .B1(net967),
    .B2(net829),
    .X(\t$5705 ));
 sky130_fd_sc_hd__xor2_1 \U$$2545  (.A(\t$5705 ),
    .B(net1409),
    .X(booth_b36_m36));
 sky130_fd_sc_hd__a22o_1 \U$$2546  (.A1(net965),
    .A2(net553),
    .B1(net957),
    .B2(net826),
    .X(\t$5706 ));
 sky130_fd_sc_hd__xor2_1 \U$$2547  (.A(\t$5706 ),
    .B(net1405),
    .X(booth_b36_m37));
 sky130_fd_sc_hd__a22o_1 \U$$2548  (.A1(net957),
    .A2(net553),
    .B1(net949),
    .B2(net826),
    .X(\t$5707 ));
 sky130_fd_sc_hd__xor2_1 \U$$2549  (.A(\t$5707 ),
    .B(net1405),
    .X(booth_b36_m38));
 sky130_fd_sc_hd__a22o_1 \U$$255  (.A1(net1615),
    .A2(net626),
    .B1(net1607),
    .B2(net899),
    .X(\t$4535 ));
 sky130_fd_sc_hd__a22o_1 \U$$2550  (.A1(net950),
    .A2(net555),
    .B1(net942),
    .B2(net828),
    .X(\t$5708 ));
 sky130_fd_sc_hd__xor2_1 \U$$2551  (.A(\t$5708 ),
    .B(net1409),
    .X(booth_b36_m39));
 sky130_fd_sc_hd__a22o_1 \U$$2552  (.A1(net942),
    .A2(net555),
    .B1(net926),
    .B2(net828),
    .X(\t$5709 ));
 sky130_fd_sc_hd__xor2_1 \U$$2553  (.A(\t$5709 ),
    .B(net1409),
    .X(booth_b36_m40));
 sky130_fd_sc_hd__a22o_1 \U$$2554  (.A1(net927),
    .A2(net555),
    .B1(net1746),
    .B2(net828),
    .X(\t$5710 ));
 sky130_fd_sc_hd__xor2_1 \U$$2555  (.A(\t$5710 ),
    .B(net1409),
    .X(booth_b36_m41));
 sky130_fd_sc_hd__a22o_1 \U$$2556  (.A1(net1748),
    .A2(net556),
    .B1(net1739),
    .B2(net829),
    .X(\t$5711 ));
 sky130_fd_sc_hd__xor2_1 \U$$2557  (.A(\t$5711 ),
    .B(net1408),
    .X(booth_b36_m42));
 sky130_fd_sc_hd__a22o_1 \U$$2558  (.A1(net1739),
    .A2(net555),
    .B1(net1731),
    .B2(net828),
    .X(\t$5712 ));
 sky130_fd_sc_hd__xor2_1 \U$$2559  (.A(\t$5712 ),
    .B(net1409),
    .X(booth_b36_m43));
 sky130_fd_sc_hd__xor2_1 \U$$256  (.A(\t$4535 ),
    .B(net1392),
    .X(booth_b2_m56));
 sky130_fd_sc_hd__a22o_1 \U$$2560  (.A1(net1731),
    .A2(net555),
    .B1(net1722),
    .B2(net828),
    .X(\t$5713 ));
 sky130_fd_sc_hd__xor2_1 \U$$2561  (.A(\t$5713 ),
    .B(net1409),
    .X(booth_b36_m44));
 sky130_fd_sc_hd__a22o_1 \U$$2562  (.A1(net1723),
    .A2(net556),
    .B1(net1713),
    .B2(net829),
    .X(\t$5714 ));
 sky130_fd_sc_hd__xor2_1 \U$$2563  (.A(\t$5714 ),
    .B(net1408),
    .X(booth_b36_m45));
 sky130_fd_sc_hd__a22o_1 \U$$2564  (.A1(net1713),
    .A2(net556),
    .B1(net1704),
    .B2(net829),
    .X(\t$5715 ));
 sky130_fd_sc_hd__xor2_1 \U$$2565  (.A(\t$5715 ),
    .B(net1408),
    .X(booth_b36_m46));
 sky130_fd_sc_hd__a22o_1 \U$$2566  (.A1(net1704),
    .A2(net555),
    .B1(net1696),
    .B2(net828),
    .X(\t$5716 ));
 sky130_fd_sc_hd__xor2_1 \U$$2567  (.A(\t$5716 ),
    .B(net1409),
    .X(booth_b36_m47));
 sky130_fd_sc_hd__a22o_1 \U$$2568  (.A1(net1696),
    .A2(net556),
    .B1(net1688),
    .B2(net829),
    .X(\t$5717 ));
 sky130_fd_sc_hd__xor2_1 \U$$2569  (.A(\t$5717 ),
    .B(net1408),
    .X(booth_b36_m48));
 sky130_fd_sc_hd__a22o_1 \U$$257  (.A1(net1604),
    .A2(net621),
    .B1(net1595),
    .B2(net894),
    .X(\t$4536 ));
 sky130_fd_sc_hd__a22o_1 \U$$2570  (.A1(net1689),
    .A2(net556),
    .B1(net1681),
    .B2(net829),
    .X(\t$5718 ));
 sky130_fd_sc_hd__xor2_1 \U$$2571  (.A(\t$5718 ),
    .B(net1411),
    .X(booth_b36_m49));
 sky130_fd_sc_hd__a22o_1 \U$$2572  (.A1(net1680),
    .A2(net556),
    .B1(net1655),
    .B2(net829),
    .X(\t$5719 ));
 sky130_fd_sc_hd__xor2_1 \U$$2573  (.A(\t$5719 ),
    .B(net1408),
    .X(booth_b36_m50));
 sky130_fd_sc_hd__a22o_1 \U$$2574  (.A1(net1655),
    .A2(net556),
    .B1(net1647),
    .B2(net829),
    .X(\t$5720 ));
 sky130_fd_sc_hd__xor2_1 \U$$2575  (.A(\t$5720 ),
    .B(net1408),
    .X(booth_b36_m51));
 sky130_fd_sc_hd__a22o_1 \U$$2576  (.A1(net1648),
    .A2(net556),
    .B1(net1640),
    .B2(net829),
    .X(\t$5721 ));
 sky130_fd_sc_hd__xor2_1 \U$$2577  (.A(\t$5721 ),
    .B(net1411),
    .X(booth_b36_m52));
 sky130_fd_sc_hd__a22o_1 \U$$2578  (.A1(net1640),
    .A2(net555),
    .B1(net1632),
    .B2(net828),
    .X(\t$5722 ));
 sky130_fd_sc_hd__xor2_1 \U$$2579  (.A(\t$5722 ),
    .B(net1409),
    .X(booth_b36_m53));
 sky130_fd_sc_hd__xor2_1 \U$$258  (.A(\t$4536 ),
    .B(net1387),
    .X(booth_b2_m57));
 sky130_fd_sc_hd__a22o_1 \U$$2580  (.A1(net1634),
    .A2(net557),
    .B1(net1624),
    .B2(net830),
    .X(\t$5723 ));
 sky130_fd_sc_hd__xor2_1 \U$$2581  (.A(\t$5723 ),
    .B(net1410),
    .X(booth_b36_m54));
 sky130_fd_sc_hd__a22o_1 \U$$2582  (.A1(net1624),
    .A2(net557),
    .B1(net1616),
    .B2(net830),
    .X(\t$5724 ));
 sky130_fd_sc_hd__xor2_1 \U$$2583  (.A(\t$5724 ),
    .B(net1410),
    .X(booth_b36_m55));
 sky130_fd_sc_hd__a22o_1 \U$$2584  (.A1(net1618),
    .A2(net557),
    .B1(net1609),
    .B2(net830),
    .X(\t$5725 ));
 sky130_fd_sc_hd__xor2_1 \U$$2585  (.A(\t$5725 ),
    .B(net1410),
    .X(booth_b36_m56));
 sky130_fd_sc_hd__a22o_1 \U$$2586  (.A1(net1611),
    .A2(net557),
    .B1(net1599),
    .B2(net830),
    .X(\t$5726 ));
 sky130_fd_sc_hd__xor2_1 \U$$2587  (.A(\t$5726 ),
    .B(net1410),
    .X(booth_b36_m57));
 sky130_fd_sc_hd__a22o_1 \U$$2588  (.A1(net1599),
    .A2(net557),
    .B1(net1593),
    .B2(net830),
    .X(\t$5727 ));
 sky130_fd_sc_hd__xor2_1 \U$$2589  (.A(\t$5727 ),
    .B(net1410),
    .X(booth_b36_m58));
 sky130_fd_sc_hd__a22o_1 \U$$259  (.A1(net1596),
    .A2(net622),
    .B1(net1587),
    .B2(net895),
    .X(\t$4537 ));
 sky130_fd_sc_hd__a22o_1 \U$$2590  (.A1(net1593),
    .A2(net557),
    .B1(net1585),
    .B2(net830),
    .X(\t$5728 ));
 sky130_fd_sc_hd__xor2_1 \U$$2591  (.A(\t$5728 ),
    .B(net1410),
    .X(booth_b36_m59));
 sky130_fd_sc_hd__a22o_1 \U$$2592  (.A1(net1585),
    .A2(net557),
    .B1(net1555),
    .B2(net830),
    .X(\t$5729 ));
 sky130_fd_sc_hd__xor2_1 \U$$2593  (.A(\t$5729 ),
    .B(net1410),
    .X(booth_b36_m60));
 sky130_fd_sc_hd__a22o_1 \U$$2594  (.A1(net1557),
    .A2(net558),
    .B1(net1550),
    .B2(net831),
    .X(\t$5730 ));
 sky130_fd_sc_hd__xor2_1 \U$$2595  (.A(\t$5730 ),
    .B(net1410),
    .X(booth_b36_m61));
 sky130_fd_sc_hd__a22o_1 \U$$2596  (.A1(net1550),
    .A2(net558),
    .B1(net1542),
    .B2(net831),
    .X(\t$5731 ));
 sky130_fd_sc_hd__xor2_1 \U$$2597  (.A(\t$5731 ),
    .B(net1411),
    .X(booth_b36_m62));
 sky130_fd_sc_hd__a22o_1 \U$$2598  (.A1(net1542),
    .A2(net558),
    .B1(net1534),
    .B2(net831),
    .X(\t$5732 ));
 sky130_fd_sc_hd__xor2_1 \U$$2599  (.A(\t$5732 ),
    .B(net1411),
    .X(booth_b36_m63));
 sky130_fd_sc_hd__a22o_1 \U$$26  (.A1(net1499),
    .A2(net446),
    .B1(net1224),
    .B2(net688),
    .X(\t$4420 ));
 sky130_fd_sc_hd__xor2_1 \U$$260  (.A(\t$4537 ),
    .B(net1388),
    .X(booth_b2_m58));
 sky130_fd_sc_hd__a22o_1 \U$$2600  (.A1(net1534),
    .A2(net557),
    .B1(net1778),
    .B2(net830),
    .X(\t$5733 ));
 sky130_fd_sc_hd__xor2_1 \U$$2601  (.A(\t$5733 ),
    .B(net1411),
    .X(booth_b36_m64));
 sky130_fd_sc_hd__inv_1 \U$$2602  (.A(net1411),
    .Y(\notsign$5734 ));
 sky130_fd_sc_hd__inv_1 \U$$2603  (.A(net1408),
    .Y(\notblock$5735[0] ));
 sky130_fd_sc_hd__inv_1 \U$$2604  (.A(net32),
    .Y(\notblock$5735[1] ));
 sky130_fd_sc_hd__inv_1 \U$$2605  (.A(net1397),
    .Y(\notblock$5735[2] ));
 sky130_fd_sc_hd__and2_1 \U$$2606  (.A(net1397),
    .B(\notblock$5735[1] ),
    .X(\t$5736 ));
 sky130_fd_sc_hd__a32o_1 \U$$2607  (.A1(\notblock$5735[2] ),
    .A2(net32),
    .A3(net1408),
    .B1(\t$5736 ),
    .B2(\notblock$5735[0] ),
    .X(\sel_0$5737 ));
 sky130_fd_sc_hd__xor2_1 \U$$2608  (.A(net32),
    .B(net1411),
    .X(\sel_1$5738 ));
 sky130_fd_sc_hd__a22o_1 \U$$2609  (.A1(net1779),
    .A2(net543),
    .B1(net1227),
    .B2(net816),
    .X(\t$5739 ));
 sky130_fd_sc_hd__a22o_1 \U$$261  (.A1(net1586),
    .A2(net621),
    .B1(net1578),
    .B2(net894),
    .X(\t$4538 ));
 sky130_fd_sc_hd__xor2_1 \U$$2610  (.A(\t$5739 ),
    .B(net1394),
    .X(booth_b38_m0));
 sky130_fd_sc_hd__a22o_1 \U$$2611  (.A1(net1228),
    .A2(net544),
    .B1(net1123),
    .B2(net817),
    .X(\t$5740 ));
 sky130_fd_sc_hd__xor2_1 \U$$2612  (.A(\t$5740 ),
    .B(net1395),
    .X(booth_b38_m1));
 sky130_fd_sc_hd__a22o_1 \U$$2613  (.A1(net1123),
    .A2(net544),
    .B1(net1033),
    .B2(net817),
    .X(\t$5741 ));
 sky130_fd_sc_hd__xor2_1 \U$$2614  (.A(\t$5741 ),
    .B(net1395),
    .X(booth_b38_m2));
 sky130_fd_sc_hd__a22o_1 \U$$2615  (.A1(net1031),
    .A2(net543),
    .B1(net932),
    .B2(net816),
    .X(\t$5742 ));
 sky130_fd_sc_hd__xor2_1 \U$$2616  (.A(\t$5742 ),
    .B(net1394),
    .X(booth_b38_m3));
 sky130_fd_sc_hd__a22o_1 \U$$2617  (.A1(net932),
    .A2(net543),
    .B1(net1671),
    .B2(net816),
    .X(\t$5743 ));
 sky130_fd_sc_hd__xor2_1 \U$$2618  (.A(\t$5743 ),
    .B(net1394),
    .X(booth_b38_m4));
 sky130_fd_sc_hd__a22o_1 \U$$2619  (.A1(net1673),
    .A2(net543),
    .B1(net1562),
    .B2(net816),
    .X(\t$5744 ));
 sky130_fd_sc_hd__xor2_1 \U$$262  (.A(\t$4538 ),
    .B(net1387),
    .X(booth_b2_m59));
 sky130_fd_sc_hd__xor2_1 \U$$2620  (.A(\t$5744 ),
    .B(net1394),
    .X(booth_b38_m5));
 sky130_fd_sc_hd__a22o_1 \U$$2621  (.A1(net1562),
    .A2(net543),
    .B1(net1520),
    .B2(net816),
    .X(\t$5745 ));
 sky130_fd_sc_hd__xor2_1 \U$$2622  (.A(\t$5745 ),
    .B(net1394),
    .X(booth_b38_m6));
 sky130_fd_sc_hd__a22o_1 \U$$2623  (.A1(net1520),
    .A2(net543),
    .B1(net1512),
    .B2(net816),
    .X(\t$5746 ));
 sky130_fd_sc_hd__xor2_1 \U$$2624  (.A(\t$5746 ),
    .B(net1395),
    .X(booth_b38_m7));
 sky130_fd_sc_hd__a22o_1 \U$$2625  (.A1(net1512),
    .A2(net543),
    .B1(net1504),
    .B2(net816),
    .X(\t$5747 ));
 sky130_fd_sc_hd__xor2_1 \U$$2626  (.A(\t$5747 ),
    .B(net1395),
    .X(booth_b38_m8));
 sky130_fd_sc_hd__a22o_1 \U$$2627  (.A1(net1504),
    .A2(net543),
    .B1(net1495),
    .B2(net816),
    .X(\t$5748 ));
 sky130_fd_sc_hd__xor2_1 \U$$2628  (.A(\t$5748 ),
    .B(net1394),
    .X(booth_b38_m9));
 sky130_fd_sc_hd__a22o_1 \U$$2629  (.A1(net1495),
    .A2(net543),
    .B1(net1220),
    .B2(net816),
    .X(\t$5749 ));
 sky130_fd_sc_hd__a22o_1 \U$$263  (.A1(net1578),
    .A2(net621),
    .B1(net1551),
    .B2(net894),
    .X(\t$4539 ));
 sky130_fd_sc_hd__xor2_1 \U$$2630  (.A(\t$5749 ),
    .B(net1394),
    .X(booth_b38_m10));
 sky130_fd_sc_hd__a22o_1 \U$$2631  (.A1(net1222),
    .A2(net544),
    .B1(net1214),
    .B2(net817),
    .X(\t$5750 ));
 sky130_fd_sc_hd__xor2_1 \U$$2632  (.A(\t$5750 ),
    .B(net1395),
    .X(booth_b38_m11));
 sky130_fd_sc_hd__a22o_1 \U$$2633  (.A1(net1217),
    .A2(net549),
    .B1(net1206),
    .B2(net822),
    .X(\t$5751 ));
 sky130_fd_sc_hd__xor2_1 \U$$2634  (.A(\t$5751 ),
    .B(net1399),
    .X(booth_b38_m12));
 sky130_fd_sc_hd__a22o_1 \U$$2635  (.A1(net1206),
    .A2(net549),
    .B1(net1199),
    .B2(net822),
    .X(\t$5752 ));
 sky130_fd_sc_hd__xor2_1 \U$$2636  (.A(\t$5752 ),
    .B(net1399),
    .X(booth_b38_m13));
 sky130_fd_sc_hd__a22o_1 \U$$2637  (.A1(net1199),
    .A2(net549),
    .B1(net1180),
    .B2(net822),
    .X(\t$5753 ));
 sky130_fd_sc_hd__xor2_1 \U$$2638  (.A(\t$5753 ),
    .B(net1399),
    .X(booth_b38_m14));
 sky130_fd_sc_hd__a22o_1 \U$$2639  (.A1(net1180),
    .A2(net549),
    .B1(net1171),
    .B2(net822),
    .X(\t$5754 ));
 sky130_fd_sc_hd__xor2_1 \U$$264  (.A(\t$4539 ),
    .B(net1387),
    .X(booth_b2_m60));
 sky130_fd_sc_hd__xor2_1 \U$$2640  (.A(\t$5754 ),
    .B(net1399),
    .X(booth_b38_m15));
 sky130_fd_sc_hd__a22o_1 \U$$2641  (.A1(net1171),
    .A2(net549),
    .B1(net1162),
    .B2(net822),
    .X(\t$5755 ));
 sky130_fd_sc_hd__xor2_1 \U$$2642  (.A(\t$5755 ),
    .B(net1399),
    .X(booth_b38_m16));
 sky130_fd_sc_hd__a22o_1 \U$$2643  (.A1(net1162),
    .A2(net549),
    .B1(net1150),
    .B2(net822),
    .X(\t$5756 ));
 sky130_fd_sc_hd__xor2_1 \U$$2644  (.A(\t$5756 ),
    .B(net1399),
    .X(booth_b38_m17));
 sky130_fd_sc_hd__a22o_1 \U$$2645  (.A1(net1150),
    .A2(net549),
    .B1(net1144),
    .B2(net822),
    .X(\t$5757 ));
 sky130_fd_sc_hd__xor2_1 \U$$2646  (.A(\t$5757 ),
    .B(net1399),
    .X(booth_b38_m18));
 sky130_fd_sc_hd__a22o_1 \U$$2647  (.A1(net1143),
    .A2(net544),
    .B1(net1134),
    .B2(net817),
    .X(\t$5758 ));
 sky130_fd_sc_hd__xor2_1 \U$$2648  (.A(\t$5758 ),
    .B(net1402),
    .X(booth_b38_m19));
 sky130_fd_sc_hd__a22o_1 \U$$2649  (.A1(net1134),
    .A2(net544),
    .B1(net1118),
    .B2(net817),
    .X(\t$5759 ));
 sky130_fd_sc_hd__a22o_1 \U$$265  (.A1(net1551),
    .A2(net621),
    .B1(net1543),
    .B2(net894),
    .X(\t$4540 ));
 sky130_fd_sc_hd__xor2_1 \U$$2650  (.A(\t$5759 ),
    .B(net1402),
    .X(booth_b38_m20));
 sky130_fd_sc_hd__a22o_1 \U$$2651  (.A1(net1116),
    .A2(net544),
    .B1(net1107),
    .B2(net817),
    .X(\t$5760 ));
 sky130_fd_sc_hd__xor2_1 \U$$2652  (.A(\t$5760 ),
    .B(net1395),
    .X(booth_b38_m21));
 sky130_fd_sc_hd__a22o_1 \U$$2653  (.A1(net1107),
    .A2(net550),
    .B1(net1098),
    .B2(net823),
    .X(\t$5761 ));
 sky130_fd_sc_hd__xor2_1 \U$$2654  (.A(\t$5761 ),
    .B(net1395),
    .X(booth_b38_m22));
 sky130_fd_sc_hd__a22o_1 \U$$2655  (.A1(net1099),
    .A2(net544),
    .B1(net1093),
    .B2(net817),
    .X(\t$5762 ));
 sky130_fd_sc_hd__xor2_1 \U$$2656  (.A(\t$5762 ),
    .B(net1395),
    .X(booth_b38_m23));
 sky130_fd_sc_hd__a22o_1 \U$$2657  (.A1(net1096),
    .A2(net546),
    .B1(net1087),
    .B2(net819),
    .X(\t$5763 ));
 sky130_fd_sc_hd__xor2_1 \U$$2658  (.A(\t$5763 ),
    .B(net1397),
    .X(booth_b38_m24));
 sky130_fd_sc_hd__a22o_1 \U$$2659  (.A1(net1086),
    .A2(net544),
    .B1(net1076),
    .B2(net817),
    .X(\t$5764 ));
 sky130_fd_sc_hd__xor2_1 \U$$266  (.A(\t$4540 ),
    .B(net1387),
    .X(booth_b2_m61));
 sky130_fd_sc_hd__xor2_1 \U$$2660  (.A(\t$5764 ),
    .B(net1395),
    .X(booth_b38_m25));
 sky130_fd_sc_hd__a22o_1 \U$$2661  (.A1(net1075),
    .A2(net549),
    .B1(net1067),
    .B2(net822),
    .X(\t$5765 ));
 sky130_fd_sc_hd__xor2_1 \U$$2662  (.A(\t$5765 ),
    .B(net1399),
    .X(booth_b38_m26));
 sky130_fd_sc_hd__a22o_1 \U$$2663  (.A1(net1067),
    .A2(net549),
    .B1(net1058),
    .B2(net822),
    .X(\t$5766 ));
 sky130_fd_sc_hd__xor2_1 \U$$2664  (.A(\t$5766 ),
    .B(net1399),
    .X(booth_b38_m27));
 sky130_fd_sc_hd__a22o_1 \U$$2665  (.A1(net1058),
    .A2(net549),
    .B1(net1054),
    .B2(net822),
    .X(\t$5767 ));
 sky130_fd_sc_hd__xor2_1 \U$$2666  (.A(\t$5767 ),
    .B(net1399),
    .X(booth_b38_m28));
 sky130_fd_sc_hd__a22o_1 \U$$2667  (.A1(net1053),
    .A2(net547),
    .B1(net1045),
    .B2(net820),
    .X(\t$5768 ));
 sky130_fd_sc_hd__xor2_1 \U$$2668  (.A(\t$5768 ),
    .B(net1402),
    .X(booth_b38_m29));
 sky130_fd_sc_hd__a22o_1 \U$$2669  (.A1(net1045),
    .A2(net547),
    .B1(net1029),
    .B2(net820),
    .X(\t$5769 ));
 sky130_fd_sc_hd__a22o_1 \U$$267  (.A1(net1543),
    .A2(net621),
    .B1(net1535),
    .B2(net894),
    .X(\t$4541 ));
 sky130_fd_sc_hd__xor2_1 \U$$2670  (.A(\t$5769 ),
    .B(net1400),
    .X(booth_b38_m30));
 sky130_fd_sc_hd__a22o_1 \U$$2671  (.A1(net1029),
    .A2(net547),
    .B1(net1021),
    .B2(net820),
    .X(\t$5770 ));
 sky130_fd_sc_hd__xor2_1 \U$$2672  (.A(\t$5770 ),
    .B(net1400),
    .X(booth_b38_m31));
 sky130_fd_sc_hd__a22o_1 \U$$2673  (.A1(net1019),
    .A2(net546),
    .B1(net1002),
    .B2(net819),
    .X(\t$5771 ));
 sky130_fd_sc_hd__xor2_1 \U$$2674  (.A(\t$5771 ),
    .B(net1397),
    .X(booth_b38_m32));
 sky130_fd_sc_hd__a22o_1 \U$$2675  (.A1(net1002),
    .A2(net546),
    .B1(net994),
    .B2(net819),
    .X(\t$5772 ));
 sky130_fd_sc_hd__xor2_1 \U$$2676  (.A(\t$5772 ),
    .B(net1397),
    .X(booth_b38_m33));
 sky130_fd_sc_hd__a22o_1 \U$$2677  (.A1(net994),
    .A2(net546),
    .B1(net984),
    .B2(net819),
    .X(\t$5773 ));
 sky130_fd_sc_hd__xor2_1 \U$$2678  (.A(\t$5773 ),
    .B(net1397),
    .X(booth_b38_m34));
 sky130_fd_sc_hd__a22o_1 \U$$2679  (.A1(net983),
    .A2(net544),
    .B1(net974),
    .B2(net817),
    .X(\t$5774 ));
 sky130_fd_sc_hd__xor2_1 \U$$268  (.A(\t$4541 ),
    .B(net1388),
    .X(booth_b2_m62));
 sky130_fd_sc_hd__xor2_1 \U$$2680  (.A(\t$5774 ),
    .B(net1394),
    .X(booth_b38_m35));
 sky130_fd_sc_hd__a22o_1 \U$$2681  (.A1(net974),
    .A2(net543),
    .B1(net965),
    .B2(net816),
    .X(\t$5775 ));
 sky130_fd_sc_hd__xor2_1 \U$$2682  (.A(\t$5775 ),
    .B(net1394),
    .X(booth_b38_m36));
 sky130_fd_sc_hd__a22o_1 \U$$2683  (.A1(net966),
    .A2(net545),
    .B1(net959),
    .B2(net818),
    .X(\t$5776 ));
 sky130_fd_sc_hd__xor2_1 \U$$2684  (.A(\t$5776 ),
    .B(net1396),
    .X(booth_b38_m37));
 sky130_fd_sc_hd__a22o_1 \U$$2685  (.A1(net959),
    .A2(net545),
    .B1(net950),
    .B2(net818),
    .X(\t$5777 ));
 sky130_fd_sc_hd__xor2_1 \U$$2686  (.A(\t$5777 ),
    .B(net1396),
    .X(booth_b38_m38));
 sky130_fd_sc_hd__a22o_1 \U$$2687  (.A1(net951),
    .A2(net545),
    .B1(net943),
    .B2(net818),
    .X(\t$5778 ));
 sky130_fd_sc_hd__xor2_1 \U$$2688  (.A(\t$5778 ),
    .B(net1396),
    .X(booth_b38_m39));
 sky130_fd_sc_hd__a22o_1 \U$$2689  (.A1(net943),
    .A2(net546),
    .B1(net927),
    .B2(net819),
    .X(\t$5779 ));
 sky130_fd_sc_hd__a22o_1 \U$$269  (.A1(net1539),
    .A2(net626),
    .B1(net1531),
    .B2(net899),
    .X(\t$4542 ));
 sky130_fd_sc_hd__xor2_1 \U$$2690  (.A(\t$5779 ),
    .B(net1397),
    .X(booth_b38_m40));
 sky130_fd_sc_hd__a22o_1 \U$$2691  (.A1(net926),
    .A2(net545),
    .B1(net1747),
    .B2(net818),
    .X(\t$5780 ));
 sky130_fd_sc_hd__xor2_1 \U$$2692  (.A(\t$5780 ),
    .B(net1396),
    .X(booth_b38_m41));
 sky130_fd_sc_hd__a22o_1 \U$$2693  (.A1(net1748),
    .A2(net546),
    .B1(net1740),
    .B2(net819),
    .X(\t$5781 ));
 sky130_fd_sc_hd__xor2_1 \U$$2694  (.A(\t$5781 ),
    .B(net1397),
    .X(booth_b38_m42));
 sky130_fd_sc_hd__a22o_1 \U$$2695  (.A1(net1740),
    .A2(net545),
    .B1(net1732),
    .B2(net818),
    .X(\t$5782 ));
 sky130_fd_sc_hd__xor2_1 \U$$2696  (.A(\t$5782 ),
    .B(net1396),
    .X(booth_b38_m43));
 sky130_fd_sc_hd__a22o_1 \U$$2697  (.A1(net1731),
    .A2(net546),
    .B1(net1722),
    .B2(net819),
    .X(\t$5783 ));
 sky130_fd_sc_hd__xor2_1 \U$$2698  (.A(\t$5783 ),
    .B(net1396),
    .X(booth_b38_m44));
 sky130_fd_sc_hd__a22o_1 \U$$2699  (.A1(net1722),
    .A2(net545),
    .B1(net1713),
    .B2(net818),
    .X(\t$5784 ));
 sky130_fd_sc_hd__xor2_1 \U$$27  (.A(\t$4420 ),
    .B(net1573),
    .X(booth_b0_m10));
 sky130_fd_sc_hd__xor2_1 \U$$270  (.A(\t$4542 ),
    .B(net1392),
    .X(booth_b2_m63));
 sky130_fd_sc_hd__xor2_1 \U$$2700  (.A(\t$5784 ),
    .B(net1396),
    .X(booth_b38_m45));
 sky130_fd_sc_hd__a22o_1 \U$$2701  (.A1(net1713),
    .A2(net545),
    .B1(net1704),
    .B2(net818),
    .X(\t$5785 ));
 sky130_fd_sc_hd__xor2_1 \U$$2702  (.A(\t$5785 ),
    .B(net1396),
    .X(booth_b38_m46));
 sky130_fd_sc_hd__a22o_1 \U$$2703  (.A1(net1704),
    .A2(net545),
    .B1(net1696),
    .B2(net818),
    .X(\t$5786 ));
 sky130_fd_sc_hd__xor2_1 \U$$2704  (.A(\t$5786 ),
    .B(net1396),
    .X(booth_b38_m47));
 sky130_fd_sc_hd__a22o_1 \U$$2705  (.A1(net1696),
    .A2(net545),
    .B1(net1688),
    .B2(net818),
    .X(\t$5787 ));
 sky130_fd_sc_hd__xor2_1 \U$$2706  (.A(\t$5787 ),
    .B(net1396),
    .X(booth_b38_m48));
 sky130_fd_sc_hd__a22o_1 \U$$2707  (.A1(net1688),
    .A2(net545),
    .B1(net1680),
    .B2(net818),
    .X(\t$5788 ));
 sky130_fd_sc_hd__xor2_1 \U$$2708  (.A(\t$5788 ),
    .B(net1398),
    .X(booth_b38_m49));
 sky130_fd_sc_hd__a22o_1 \U$$2709  (.A1(net1681),
    .A2(net546),
    .B1(net1656),
    .B2(net819),
    .X(\t$5789 ));
 sky130_fd_sc_hd__a22o_1 \U$$271  (.A1(net1531),
    .A2(net626),
    .B1(net1780),
    .B2(net899),
    .X(\t$4543 ));
 sky130_fd_sc_hd__xor2_1 \U$$2710  (.A(\t$5789 ),
    .B(net1397),
    .X(booth_b38_m50));
 sky130_fd_sc_hd__a22o_1 \U$$2711  (.A1(net1656),
    .A2(net546),
    .B1(net1648),
    .B2(net819),
    .X(\t$5790 ));
 sky130_fd_sc_hd__xor2_1 \U$$2712  (.A(\t$5790 ),
    .B(net1397),
    .X(booth_b38_m51));
 sky130_fd_sc_hd__a22o_1 \U$$2713  (.A1(net1651),
    .A2(net548),
    .B1(net1643),
    .B2(net821),
    .X(\t$5791 ));
 sky130_fd_sc_hd__xor2_1 \U$$2714  (.A(\t$5791 ),
    .B(net1401),
    .X(booth_b38_m52));
 sky130_fd_sc_hd__a22o_1 \U$$2715  (.A1(net1643),
    .A2(net548),
    .B1(net1634),
    .B2(net821),
    .X(\t$5792 ));
 sky130_fd_sc_hd__xor2_1 \U$$2716  (.A(\t$5792 ),
    .B(net1401),
    .X(booth_b38_m53));
 sky130_fd_sc_hd__a22o_1 \U$$2717  (.A1(net1635),
    .A2(net547),
    .B1(net1627),
    .B2(net820),
    .X(\t$5793 ));
 sky130_fd_sc_hd__xor2_1 \U$$2718  (.A(\t$5793 ),
    .B(net1400),
    .X(booth_b38_m54));
 sky130_fd_sc_hd__a22o_1 \U$$2719  (.A1(net1627),
    .A2(net547),
    .B1(net1619),
    .B2(net820),
    .X(\t$5794 ));
 sky130_fd_sc_hd__xor2_1 \U$$272  (.A(\t$4543 ),
    .B(net1392),
    .X(booth_b2_m64));
 sky130_fd_sc_hd__xor2_1 \U$$2720  (.A(\t$5794 ),
    .B(net1400),
    .X(booth_b38_m55));
 sky130_fd_sc_hd__a22o_1 \U$$2721  (.A1(net1618),
    .A2(net547),
    .B1(net1609),
    .B2(net820),
    .X(\t$5795 ));
 sky130_fd_sc_hd__xor2_1 \U$$2722  (.A(\t$5795 ),
    .B(net1400),
    .X(booth_b38_m56));
 sky130_fd_sc_hd__a22o_1 \U$$2723  (.A1(net1611),
    .A2(net547),
    .B1(net1603),
    .B2(net820),
    .X(\t$5796 ));
 sky130_fd_sc_hd__xor2_1 \U$$2724  (.A(\t$5796 ),
    .B(net1400),
    .X(booth_b38_m57));
 sky130_fd_sc_hd__a22o_1 \U$$2725  (.A1(net1603),
    .A2(net547),
    .B1(net1593),
    .B2(net820),
    .X(\t$5797 ));
 sky130_fd_sc_hd__xor2_1 \U$$2726  (.A(\t$5797 ),
    .B(net1400),
    .X(booth_b38_m58));
 sky130_fd_sc_hd__a22o_1 \U$$2727  (.A1(net1592),
    .A2(net548),
    .B1(net1584),
    .B2(net821),
    .X(\t$5798 ));
 sky130_fd_sc_hd__xor2_1 \U$$2728  (.A(\t$5798 ),
    .B(net1400),
    .X(booth_b38_m59));
 sky130_fd_sc_hd__a22o_1 \U$$2729  (.A1(net1584),
    .A2(net547),
    .B1(net1557),
    .B2(net820),
    .X(\t$5799 ));
 sky130_fd_sc_hd__inv_1 \U$$273  (.A(net1393),
    .Y(\notsign$4544 ));
 sky130_fd_sc_hd__xor2_1 \U$$2730  (.A(\t$5799 ),
    .B(net1400),
    .X(booth_b38_m60));
 sky130_fd_sc_hd__a22o_1 \U$$2731  (.A1(net1557),
    .A2(net548),
    .B1(net1550),
    .B2(net821),
    .X(\t$5800 ));
 sky130_fd_sc_hd__xor2_1 \U$$2732  (.A(\t$5800 ),
    .B(net1400),
    .X(booth_b38_m61));
 sky130_fd_sc_hd__a22o_1 \U$$2733  (.A1(net1550),
    .A2(net548),
    .B1(net1542),
    .B2(net821),
    .X(\t$5801 ));
 sky130_fd_sc_hd__xor2_1 \U$$2734  (.A(\t$5801 ),
    .B(net1401),
    .X(booth_b38_m62));
 sky130_fd_sc_hd__a22o_1 \U$$2735  (.A1(net1542),
    .A2(net547),
    .B1(net1534),
    .B2(net820),
    .X(\t$5802 ));
 sky130_fd_sc_hd__xor2_1 \U$$2736  (.A(\t$5802 ),
    .B(net1401),
    .X(booth_b38_m63));
 sky130_fd_sc_hd__a22o_1 \U$$2737  (.A1(net1534),
    .A2(net548),
    .B1(net1781),
    .B2(net821),
    .X(\t$5803 ));
 sky130_fd_sc_hd__xor2_1 \U$$2738  (.A(\t$5803 ),
    .B(net1401),
    .X(booth_b38_m64));
 sky130_fd_sc_hd__inv_1 \U$$2739  (.A(net1401),
    .Y(\notsign$5804 ));
 sky130_fd_sc_hd__inv_1 \U$$274  (.A(net1388),
    .Y(\notblock$4545[0] ));
 sky130_fd_sc_hd__inv_1 \U$$2740  (.A(net1398),
    .Y(\notblock$5805[0] ));
 sky130_fd_sc_hd__inv_1 \U$$2741  (.A(net35),
    .Y(\notblock$5805[1] ));
 sky130_fd_sc_hd__inv_1 \U$$2742  (.A(net1378),
    .Y(\notblock$5805[2] ));
 sky130_fd_sc_hd__and2_1 \U$$2743  (.A(net1378),
    .B(\notblock$5805[1] ),
    .X(\t$5806 ));
 sky130_fd_sc_hd__a32o_1 \U$$2744  (.A1(\notblock$5805[2] ),
    .A2(net35),
    .A3(net1398),
    .B1(\t$5806 ),
    .B2(\notblock$5805[0] ),
    .X(\sel_0$5807 ));
 sky130_fd_sc_hd__xor2_1 \U$$2745  (.A(net35),
    .B(net1398),
    .X(\sel_1$5808 ));
 sky130_fd_sc_hd__a22o_1 \U$$2746  (.A1(net1782),
    .A2(net535),
    .B1(net1227),
    .B2(net808),
    .X(\t$5809 ));
 sky130_fd_sc_hd__xor2_1 \U$$2747  (.A(\t$5809 ),
    .B(net1376),
    .X(booth_b40_m0));
 sky130_fd_sc_hd__a22o_1 \U$$2748  (.A1(net1227),
    .A2(net535),
    .B1(net1122),
    .B2(net808),
    .X(\t$5810 ));
 sky130_fd_sc_hd__xor2_1 \U$$2749  (.A(\t$5810 ),
    .B(net1376),
    .X(booth_b40_m1));
 sky130_fd_sc_hd__inv_1 \U$$275  (.A(net45),
    .Y(\notblock$4545[1] ));
 sky130_fd_sc_hd__a22o_1 \U$$2750  (.A1(net1122),
    .A2(net535),
    .B1(net1031),
    .B2(net808),
    .X(\t$5811 ));
 sky130_fd_sc_hd__xor2_1 \U$$2751  (.A(\t$5811 ),
    .B(net1376),
    .X(booth_b40_m2));
 sky130_fd_sc_hd__a22o_1 \U$$2752  (.A1(net1031),
    .A2(net535),
    .B1(net934),
    .B2(net808),
    .X(\t$5812 ));
 sky130_fd_sc_hd__xor2_1 \U$$2753  (.A(\t$5812 ),
    .B(net1376),
    .X(booth_b40_m3));
 sky130_fd_sc_hd__a22o_1 \U$$2754  (.A1(net934),
    .A2(net535),
    .B1(net1673),
    .B2(net808),
    .X(\t$5813 ));
 sky130_fd_sc_hd__xor2_1 \U$$2755  (.A(\t$5813 ),
    .B(net1376),
    .X(booth_b40_m4));
 sky130_fd_sc_hd__a22o_1 \U$$2756  (.A1(net1672),
    .A2(net536),
    .B1(net1562),
    .B2(net809),
    .X(\t$5814 ));
 sky130_fd_sc_hd__xor2_1 \U$$2757  (.A(\t$5814 ),
    .B(net1377),
    .X(booth_b40_m5));
 sky130_fd_sc_hd__a22o_1 \U$$2758  (.A1(net1562),
    .A2(net536),
    .B1(net1521),
    .B2(net809),
    .X(\t$5815 ));
 sky130_fd_sc_hd__xor2_1 \U$$2759  (.A(\t$5815 ),
    .B(net1377),
    .X(booth_b40_m6));
 sky130_fd_sc_hd__inv_1 \U$$276  (.A(net1275),
    .Y(\notblock$4545[2] ));
 sky130_fd_sc_hd__a22o_1 \U$$2760  (.A1(net1522),
    .A2(net535),
    .B1(net1514),
    .B2(net808),
    .X(\t$5816 ));
 sky130_fd_sc_hd__xor2_1 \U$$2761  (.A(\t$5816 ),
    .B(net1376),
    .X(booth_b40_m7));
 sky130_fd_sc_hd__a22o_1 \U$$2762  (.A1(net1512),
    .A2(net535),
    .B1(net1504),
    .B2(net808),
    .X(\t$5817 ));
 sky130_fd_sc_hd__xor2_1 \U$$2763  (.A(\t$5817 ),
    .B(net1376),
    .X(booth_b40_m8));
 sky130_fd_sc_hd__a22o_1 \U$$2764  (.A1(net1506),
    .A2(net536),
    .B1(net1497),
    .B2(net809),
    .X(\t$5818 ));
 sky130_fd_sc_hd__xor2_1 \U$$2765  (.A(\t$5818 ),
    .B(net1377),
    .X(booth_b40_m9));
 sky130_fd_sc_hd__a22o_1 \U$$2766  (.A1(net1500),
    .A2(net539),
    .B1(net1225),
    .B2(net812),
    .X(\t$5819 ));
 sky130_fd_sc_hd__xor2_1 \U$$2767  (.A(\t$5819 ),
    .B(net1381),
    .X(booth_b40_m10));
 sky130_fd_sc_hd__a22o_1 \U$$2768  (.A1(net1225),
    .A2(net539),
    .B1(net1218),
    .B2(net812),
    .X(\t$5820 ));
 sky130_fd_sc_hd__xor2_1 \U$$2769  (.A(\t$5820 ),
    .B(net1381),
    .X(booth_b40_m11));
 sky130_fd_sc_hd__and2_1 \U$$277  (.A(net1275),
    .B(\notblock$4545[1] ),
    .X(\t$4546 ));
 sky130_fd_sc_hd__a22o_1 \U$$2770  (.A1(net1218),
    .A2(net539),
    .B1(net1207),
    .B2(net812),
    .X(\t$5821 ));
 sky130_fd_sc_hd__xor2_1 \U$$2771  (.A(\t$5821 ),
    .B(net1381),
    .X(booth_b40_m12));
 sky130_fd_sc_hd__a22o_1 \U$$2772  (.A1(net1207),
    .A2(net539),
    .B1(net1199),
    .B2(net812),
    .X(\t$5822 ));
 sky130_fd_sc_hd__xor2_1 \U$$2773  (.A(\t$5822 ),
    .B(net1381),
    .X(booth_b40_m13));
 sky130_fd_sc_hd__a22o_1 \U$$2774  (.A1(net1199),
    .A2(net539),
    .B1(net1181),
    .B2(net812),
    .X(\t$5823 ));
 sky130_fd_sc_hd__xor2_1 \U$$2775  (.A(\t$5823 ),
    .B(net1381),
    .X(booth_b40_m14));
 sky130_fd_sc_hd__a22o_1 \U$$2776  (.A1(net1181),
    .A2(net539),
    .B1(net1172),
    .B2(net812),
    .X(\t$5824 ));
 sky130_fd_sc_hd__xor2_1 \U$$2777  (.A(\t$5824 ),
    .B(net1381),
    .X(booth_b40_m15));
 sky130_fd_sc_hd__a22o_1 \U$$2778  (.A1(net1172),
    .A2(net539),
    .B1(net1163),
    .B2(net812),
    .X(\t$5825 ));
 sky130_fd_sc_hd__xor2_1 \U$$2779  (.A(\t$5825 ),
    .B(net1381),
    .X(booth_b40_m16));
 sky130_fd_sc_hd__a32o_4 \U$$278  (.A1(\notblock$4545[2] ),
    .A2(net45),
    .A3(net1388),
    .B1(\t$4546 ),
    .B2(\notblock$4545[0] ),
    .X(\sel_0$4547 ));
 sky130_fd_sc_hd__a22o_1 \U$$2780  (.A1(net1161),
    .A2(net542),
    .B1(net1150),
    .B2(net815),
    .X(\t$5826 ));
 sky130_fd_sc_hd__xor2_1 \U$$2781  (.A(\t$5826 ),
    .B(net1384),
    .X(booth_b40_m17));
 sky130_fd_sc_hd__a22o_1 \U$$2782  (.A1(net1151),
    .A2(net536),
    .B1(net1141),
    .B2(net809),
    .X(\t$5827 ));
 sky130_fd_sc_hd__xor2_1 \U$$2783  (.A(\t$5827 ),
    .B(net1377),
    .X(booth_b40_m18));
 sky130_fd_sc_hd__a22o_1 \U$$2784  (.A1(net1140),
    .A2(net536),
    .B1(net1132),
    .B2(net809),
    .X(\t$5828 ));
 sky130_fd_sc_hd__xor2_1 \U$$2785  (.A(\t$5828 ),
    .B(net1377),
    .X(booth_b40_m19));
 sky130_fd_sc_hd__a22o_1 \U$$2786  (.A1(net1132),
    .A2(net535),
    .B1(net1116),
    .B2(net808),
    .X(\t$5829 ));
 sky130_fd_sc_hd__xor2_1 \U$$2787  (.A(\t$5829 ),
    .B(net1376),
    .X(booth_b40_m20));
 sky130_fd_sc_hd__a22o_1 \U$$2788  (.A1(net1120),
    .A2(net536),
    .B1(net1111),
    .B2(net809),
    .X(\t$5830 ));
 sky130_fd_sc_hd__xor2_1 \U$$2789  (.A(\t$5830 ),
    .B(net1377),
    .X(booth_b40_m21));
 sky130_fd_sc_hd__xor2_4 \U$$279  (.A(net45),
    .B(net1388),
    .X(\sel_1$4548 ));
 sky130_fd_sc_hd__a22o_1 \U$$2790  (.A1(net1110),
    .A2(net536),
    .B1(net1099),
    .B2(net809),
    .X(\t$5831 ));
 sky130_fd_sc_hd__xor2_1 \U$$2791  (.A(\t$5831 ),
    .B(net1377),
    .X(booth_b40_m22));
 sky130_fd_sc_hd__a22o_1 \U$$2792  (.A1(net1102),
    .A2(net538),
    .B1(net1094),
    .B2(net811),
    .X(\t$5832 ));
 sky130_fd_sc_hd__xor2_1 \U$$2793  (.A(\t$5832 ),
    .B(net1380),
    .X(booth_b40_m23));
 sky130_fd_sc_hd__a22o_1 \U$$2794  (.A1(net1092),
    .A2(net539),
    .B1(net1084),
    .B2(net812),
    .X(\t$5833 ));
 sky130_fd_sc_hd__xor2_1 \U$$2795  (.A(\t$5833 ),
    .B(net1381),
    .X(booth_b40_m24));
 sky130_fd_sc_hd__a22o_1 \U$$2796  (.A1(net1084),
    .A2(net539),
    .B1(net1075),
    .B2(net812),
    .X(\t$5834 ));
 sky130_fd_sc_hd__xor2_1 \U$$2797  (.A(\t$5834 ),
    .B(net1381),
    .X(booth_b40_m25));
 sky130_fd_sc_hd__a22o_1 \U$$2798  (.A1(net1078),
    .A2(net542),
    .B1(net1070),
    .B2(net815),
    .X(\t$5835 ));
 sky130_fd_sc_hd__xor2_1 \U$$2799  (.A(\t$5835 ),
    .B(net1381),
    .X(booth_b40_m26));
 sky130_fd_sc_hd__a22o_1 \U$$28  (.A1(net1224),
    .A2(net446),
    .B1(net1216),
    .B2(net688),
    .X(\t$4421 ));
 sky130_fd_sc_hd__a22o_1 \U$$280  (.A1(net1783),
    .A2(net531),
    .B1(net1231),
    .B2(net804),
    .X(\t$4549 ));
 sky130_fd_sc_hd__a22o_1 \U$$2800  (.A1(net1070),
    .A2(net539),
    .B1(net1062),
    .B2(net812),
    .X(\t$5836 ));
 sky130_fd_sc_hd__xor2_1 \U$$2801  (.A(\t$5836 ),
    .B(net1384),
    .X(booth_b40_m27));
 sky130_fd_sc_hd__a22o_1 \U$$2802  (.A1(net1062),
    .A2(net540),
    .B1(net1053),
    .B2(net813),
    .X(\t$5837 ));
 sky130_fd_sc_hd__xor2_1 \U$$2803  (.A(\t$5837 ),
    .B(net1382),
    .X(booth_b40_m28));
 sky130_fd_sc_hd__a22o_1 \U$$2804  (.A1(net1053),
    .A2(net538),
    .B1(net1045),
    .B2(net811),
    .X(\t$5838 ));
 sky130_fd_sc_hd__xor2_1 \U$$2805  (.A(\t$5838 ),
    .B(net1380),
    .X(booth_b40_m29));
 sky130_fd_sc_hd__a22o_1 \U$$2806  (.A1(net1043),
    .A2(net538),
    .B1(net1027),
    .B2(net811),
    .X(\t$5839 ));
 sky130_fd_sc_hd__xor2_1 \U$$2807  (.A(\t$5839 ),
    .B(net1380),
    .X(booth_b40_m30));
 sky130_fd_sc_hd__a22o_1 \U$$2808  (.A1(net1027),
    .A2(net538),
    .B1(net1019),
    .B2(net811),
    .X(\t$5840 ));
 sky130_fd_sc_hd__xor2_1 \U$$2809  (.A(\t$5840 ),
    .B(net1380),
    .X(booth_b40_m31));
 sky130_fd_sc_hd__xor2_1 \U$$281  (.A(\t$4549 ),
    .B(net1277),
    .X(booth_b4_m0));
 sky130_fd_sc_hd__a22o_1 \U$$2810  (.A1(net1016),
    .A2(net535),
    .B1(net999),
    .B2(net808),
    .X(\t$5841 ));
 sky130_fd_sc_hd__xor2_1 \U$$2811  (.A(\t$5841 ),
    .B(net1376),
    .X(booth_b40_m32));
 sky130_fd_sc_hd__a22o_1 \U$$2812  (.A1(net1005),
    .A2(net536),
    .B1(net991),
    .B2(net809),
    .X(\t$5842 ));
 sky130_fd_sc_hd__xor2_1 \U$$2813  (.A(\t$5842 ),
    .B(net1377),
    .X(booth_b40_m33));
 sky130_fd_sc_hd__a22o_1 \U$$2814  (.A1(net91),
    .A2(net535),
    .B1(net983),
    .B2(net808),
    .X(\t$5843 ));
 sky130_fd_sc_hd__xor2_1 \U$$2815  (.A(\t$5843 ),
    .B(net1377),
    .X(booth_b40_m34));
 sky130_fd_sc_hd__a22o_1 \U$$2816  (.A1(net984),
    .A2(net537),
    .B1(net975),
    .B2(net810),
    .X(\t$5844 ));
 sky130_fd_sc_hd__xor2_1 \U$$2817  (.A(\t$5844 ),
    .B(net1378),
    .X(booth_b40_m35));
 sky130_fd_sc_hd__a22o_1 \U$$2818  (.A1(net975),
    .A2(net537),
    .B1(net966),
    .B2(net810),
    .X(\t$5845 ));
 sky130_fd_sc_hd__xor2_1 \U$$2819  (.A(\t$5845 ),
    .B(net1378),
    .X(booth_b40_m36));
 sky130_fd_sc_hd__a22o_1 \U$$282  (.A1(net1232),
    .A2(net531),
    .B1(net1127),
    .B2(net804),
    .X(\t$4550 ));
 sky130_fd_sc_hd__a22o_1 \U$$2820  (.A1(net967),
    .A2(net537),
    .B1(net958),
    .B2(net810),
    .X(\t$5846 ));
 sky130_fd_sc_hd__xor2_1 \U$$2821  (.A(\t$5846 ),
    .B(net1378),
    .X(booth_b40_m37));
 sky130_fd_sc_hd__a22o_1 \U$$2822  (.A1(net958),
    .A2(net537),
    .B1(net951),
    .B2(net810),
    .X(\t$5847 ));
 sky130_fd_sc_hd__xor2_1 \U$$2823  (.A(\t$5847 ),
    .B(net1378),
    .X(booth_b40_m38));
 sky130_fd_sc_hd__a22o_1 \U$$2824  (.A1(net950),
    .A2(net537),
    .B1(net942),
    .B2(net810),
    .X(\t$5848 ));
 sky130_fd_sc_hd__xor2_1 \U$$2825  (.A(\t$5848 ),
    .B(net1378),
    .X(booth_b40_m39));
 sky130_fd_sc_hd__a22o_1 \U$$2826  (.A1(net943),
    .A2(net538),
    .B1(net927),
    .B2(net811),
    .X(\t$5849 ));
 sky130_fd_sc_hd__xor2_1 \U$$2827  (.A(\t$5849 ),
    .B(net1380),
    .X(booth_b40_m40));
 sky130_fd_sc_hd__a22o_1 \U$$2828  (.A1(net927),
    .A2(net538),
    .B1(net1748),
    .B2(net811),
    .X(\t$5850 ));
 sky130_fd_sc_hd__xor2_1 \U$$2829  (.A(\t$5850 ),
    .B(net1380),
    .X(booth_b40_m41));
 sky130_fd_sc_hd__xor2_1 \U$$283  (.A(\t$4550 ),
    .B(net1277),
    .X(booth_b4_m1));
 sky130_fd_sc_hd__a22o_1 \U$$2830  (.A1(net1747),
    .A2(net537),
    .B1(net1739),
    .B2(net810),
    .X(\t$5851 ));
 sky130_fd_sc_hd__xor2_1 \U$$2831  (.A(\t$5851 ),
    .B(net1378),
    .X(booth_b40_m42));
 sky130_fd_sc_hd__a22o_1 \U$$2832  (.A1(net1739),
    .A2(net537),
    .B1(net1731),
    .B2(net810),
    .X(\t$5852 ));
 sky130_fd_sc_hd__xor2_1 \U$$2833  (.A(\t$5852 ),
    .B(net1378),
    .X(booth_b40_m43));
 sky130_fd_sc_hd__a22o_1 \U$$2834  (.A1(net1731),
    .A2(net537),
    .B1(net1722),
    .B2(net810),
    .X(\t$5853 ));
 sky130_fd_sc_hd__xor2_1 \U$$2835  (.A(\t$5853 ),
    .B(net1378),
    .X(booth_b40_m44));
 sky130_fd_sc_hd__a22o_1 \U$$2836  (.A1(net1723),
    .A2(net538),
    .B1(net1714),
    .B2(net811),
    .X(\t$5854 ));
 sky130_fd_sc_hd__xor2_1 \U$$2837  (.A(\t$5854 ),
    .B(net1379),
    .X(booth_b40_m45));
 sky130_fd_sc_hd__a22o_1 \U$$2838  (.A1(net1713),
    .A2(net537),
    .B1(net1704),
    .B2(net810),
    .X(\t$5855 ));
 sky130_fd_sc_hd__xor2_1 \U$$2839  (.A(\t$5855 ),
    .B(net1379),
    .X(booth_b40_m46));
 sky130_fd_sc_hd__a22o_1 \U$$284  (.A1(net1128),
    .A2(net534),
    .B1(net1035),
    .B2(net807),
    .X(\t$4551 ));
 sky130_fd_sc_hd__a22o_1 \U$$2840  (.A1(net1705),
    .A2(net537),
    .B1(net1697),
    .B2(net810),
    .X(\t$5856 ));
 sky130_fd_sc_hd__xor2_1 \U$$2841  (.A(\t$5856 ),
    .B(net1379),
    .X(booth_b40_m47));
 sky130_fd_sc_hd__a22o_1 \U$$2842  (.A1(net1702),
    .A2(net538),
    .B1(net1692),
    .B2(net811),
    .X(\t$5857 ));
 sky130_fd_sc_hd__xor2_1 \U$$2843  (.A(\t$5857 ),
    .B(net1380),
    .X(booth_b40_m48));
 sky130_fd_sc_hd__a22o_1 \U$$2844  (.A1(net1689),
    .A2(net538),
    .B1(net1681),
    .B2(net811),
    .X(\t$5858 ));
 sky130_fd_sc_hd__xor2_1 \U$$2845  (.A(\t$5858 ),
    .B(net1380),
    .X(booth_b40_m49));
 sky130_fd_sc_hd__a22o_1 \U$$2846  (.A1(net1685),
    .A2(net541),
    .B1(net1659),
    .B2(net814),
    .X(\t$5859 ));
 sky130_fd_sc_hd__xor2_1 \U$$2847  (.A(\t$5859 ),
    .B(net1383),
    .X(booth_b40_m50));
 sky130_fd_sc_hd__a22o_1 \U$$2848  (.A1(net1659),
    .A2(net541),
    .B1(net1651),
    .B2(net814),
    .X(\t$5860 ));
 sky130_fd_sc_hd__xor2_1 \U$$2849  (.A(\t$5860 ),
    .B(net1383),
    .X(booth_b40_m51));
 sky130_fd_sc_hd__xor2_1 \U$$285  (.A(\t$4551 ),
    .B(net1277),
    .X(booth_b4_m2));
 sky130_fd_sc_hd__a22o_1 \U$$2850  (.A1(net1652),
    .A2(net540),
    .B1(net1642),
    .B2(net813),
    .X(\t$5861 ));
 sky130_fd_sc_hd__xor2_1 \U$$2851  (.A(\t$5861 ),
    .B(net1382),
    .X(booth_b40_m52));
 sky130_fd_sc_hd__a22o_1 \U$$2852  (.A1(net1644),
    .A2(net540),
    .B1(net1635),
    .B2(net813),
    .X(\t$5862 ));
 sky130_fd_sc_hd__xor2_1 \U$$2853  (.A(\t$5862 ),
    .B(net1382),
    .X(booth_b40_m53));
 sky130_fd_sc_hd__a22o_1 \U$$2854  (.A1(net1635),
    .A2(net540),
    .B1(net1626),
    .B2(net813),
    .X(\t$5863 ));
 sky130_fd_sc_hd__xor2_1 \U$$2855  (.A(\t$5863 ),
    .B(net1382),
    .X(booth_b40_m54));
 sky130_fd_sc_hd__a22o_1 \U$$2856  (.A1(net1627),
    .A2(net540),
    .B1(net1619),
    .B2(net813),
    .X(\t$5864 ));
 sky130_fd_sc_hd__xor2_1 \U$$2857  (.A(\t$5864 ),
    .B(net1382),
    .X(booth_b40_m55));
 sky130_fd_sc_hd__a22o_1 \U$$2858  (.A1(net1619),
    .A2(net540),
    .B1(net1611),
    .B2(net813),
    .X(\t$5865 ));
 sky130_fd_sc_hd__xor2_1 \U$$2859  (.A(\t$5865 ),
    .B(net1382),
    .X(booth_b40_m56));
 sky130_fd_sc_hd__a22o_1 \U$$286  (.A1(net1035),
    .A2(net531),
    .B1(net937),
    .B2(net804),
    .X(\t$4552 ));
 sky130_fd_sc_hd__a22o_1 \U$$2860  (.A1(net1609),
    .A2(net540),
    .B1(net1602),
    .B2(net813),
    .X(\t$5866 ));
 sky130_fd_sc_hd__xor2_1 \U$$2861  (.A(\t$5866 ),
    .B(net1382),
    .X(booth_b40_m57));
 sky130_fd_sc_hd__a22o_1 \U$$2862  (.A1(net1602),
    .A2(net540),
    .B1(net1592),
    .B2(net813),
    .X(\t$5867 ));
 sky130_fd_sc_hd__xor2_1 \U$$2863  (.A(\t$5867 ),
    .B(net1382),
    .X(booth_b40_m58));
 sky130_fd_sc_hd__a22o_1 \U$$2864  (.A1(net1592),
    .A2(net541),
    .B1(net1584),
    .B2(net814),
    .X(\t$5868 ));
 sky130_fd_sc_hd__xor2_1 \U$$2865  (.A(\t$5868 ),
    .B(net1382),
    .X(booth_b40_m59));
 sky130_fd_sc_hd__a22o_1 \U$$2866  (.A1(net1584),
    .A2(net541),
    .B1(net1558),
    .B2(net814),
    .X(\t$5869 ));
 sky130_fd_sc_hd__xor2_1 \U$$2867  (.A(\t$5869 ),
    .B(net1382),
    .X(booth_b40_m60));
 sky130_fd_sc_hd__a22o_1 \U$$2868  (.A1(net1558),
    .A2(net540),
    .B1(net1550),
    .B2(net813),
    .X(\t$5870 ));
 sky130_fd_sc_hd__xor2_1 \U$$2869  (.A(\t$5870 ),
    .B(net1383),
    .X(booth_b40_m61));
 sky130_fd_sc_hd__xor2_1 \U$$287  (.A(\t$4552 ),
    .B(net1277),
    .X(booth_b4_m3));
 sky130_fd_sc_hd__a22o_1 \U$$2870  (.A1(net1550),
    .A2(net540),
    .B1(net1542),
    .B2(net813),
    .X(\t$5871 ));
 sky130_fd_sc_hd__xor2_1 \U$$2871  (.A(\t$5871 ),
    .B(net1383),
    .X(booth_b40_m62));
 sky130_fd_sc_hd__a22o_1 \U$$2872  (.A1(net1540),
    .A2(net541),
    .B1(net1532),
    .B2(net814),
    .X(\t$5872 ));
 sky130_fd_sc_hd__xor2_1 \U$$2873  (.A(\t$5872 ),
    .B(net1383),
    .X(booth_b40_m63));
 sky130_fd_sc_hd__a22o_1 \U$$2874  (.A1(net1532),
    .A2(net541),
    .B1(net1784),
    .B2(net814),
    .X(\t$5873 ));
 sky130_fd_sc_hd__xor2_1 \U$$2875  (.A(\t$5873 ),
    .B(net1383),
    .X(booth_b40_m64));
 sky130_fd_sc_hd__inv_1 \U$$2876  (.A(net1383),
    .Y(\notsign$5874 ));
 sky130_fd_sc_hd__inv_1 \U$$2877  (.A(net1379),
    .Y(\notblock$5875[0] ));
 sky130_fd_sc_hd__inv_1 \U$$2878  (.A(net37),
    .Y(\notblock$5875[1] ));
 sky130_fd_sc_hd__inv_1 \U$$2879  (.A(net1369),
    .Y(\notblock$5875[2] ));
 sky130_fd_sc_hd__a22o_1 \U$$288  (.A1(net937),
    .A2(net531),
    .B1(net1675),
    .B2(net804),
    .X(\t$4553 ));
 sky130_fd_sc_hd__and2_1 \U$$2880  (.A(net1369),
    .B(\notblock$5875[1] ),
    .X(\t$5876 ));
 sky130_fd_sc_hd__a32o_4 \U$$2881  (.A1(\notblock$5875[2] ),
    .A2(net37),
    .A3(net1379),
    .B1(\t$5876 ),
    .B2(\notblock$5875[0] ),
    .X(\sel_0$5877 ));
 sky130_fd_sc_hd__xor2_4 \U$$2882  (.A(net37),
    .B(net1379),
    .X(\sel_1$5878 ));
 sky130_fd_sc_hd__a22o_1 \U$$2883  (.A1(net1785),
    .A2(net519),
    .B1(net1227),
    .B2(net792),
    .X(\t$5879 ));
 sky130_fd_sc_hd__xor2_1 \U$$2884  (.A(\t$5879 ),
    .B(net1367),
    .X(booth_b42_m0));
 sky130_fd_sc_hd__a22o_1 \U$$2885  (.A1(net1227),
    .A2(net519),
    .B1(net1122),
    .B2(net792),
    .X(\t$5880 ));
 sky130_fd_sc_hd__xor2_1 \U$$2886  (.A(\t$5880 ),
    .B(net1367),
    .X(booth_b42_m1));
 sky130_fd_sc_hd__a22o_1 \U$$2887  (.A1(net1124),
    .A2(net519),
    .B1(net1033),
    .B2(net792),
    .X(\t$5881 ));
 sky130_fd_sc_hd__xor2_1 \U$$2888  (.A(\t$5881 ),
    .B(net1367),
    .X(booth_b42_m2));
 sky130_fd_sc_hd__a22o_1 \U$$2889  (.A1(net1033),
    .A2(net520),
    .B1(net934),
    .B2(net793),
    .X(\t$5882 ));
 sky130_fd_sc_hd__xor2_1 \U$$289  (.A(\t$4553 ),
    .B(net1277),
    .X(booth_b4_m4));
 sky130_fd_sc_hd__xor2_1 \U$$2890  (.A(\t$5882 ),
    .B(net1368),
    .X(booth_b42_m3));
 sky130_fd_sc_hd__a22o_1 \U$$2891  (.A1(net935),
    .A2(net520),
    .B1(net1673),
    .B2(net793),
    .X(\t$5883 ));
 sky130_fd_sc_hd__xor2_1 \U$$2892  (.A(\t$5883 ),
    .B(net1368),
    .X(booth_b42_m4));
 sky130_fd_sc_hd__a22o_1 \U$$2893  (.A1(net1673),
    .A2(net519),
    .B1(net1562),
    .B2(net792),
    .X(\t$5884 ));
 sky130_fd_sc_hd__xor2_1 \U$$2894  (.A(\t$5884 ),
    .B(net1367),
    .X(booth_b42_m5));
 sky130_fd_sc_hd__a22o_1 \U$$2895  (.A1(net1562),
    .A2(net519),
    .B1(net1520),
    .B2(net792),
    .X(\t$5885 ));
 sky130_fd_sc_hd__xor2_1 \U$$2896  (.A(\t$5885 ),
    .B(net1367),
    .X(booth_b42_m6));
 sky130_fd_sc_hd__a22o_1 \U$$2897  (.A1(net1522),
    .A2(net519),
    .B1(net1514),
    .B2(net792),
    .X(\t$5886 ));
 sky130_fd_sc_hd__xor2_1 \U$$2898  (.A(\t$5886 ),
    .B(net1367),
    .X(booth_b42_m7));
 sky130_fd_sc_hd__a22o_1 \U$$2899  (.A1(net1516),
    .A2(net523),
    .B1(net1509),
    .B2(net796),
    .X(\t$5887 ));
 sky130_fd_sc_hd__xor2_1 \U$$29  (.A(\t$4421 ),
    .B(net1573),
    .X(booth_b0_m11));
 sky130_fd_sc_hd__a22o_1 \U$$290  (.A1(net1675),
    .A2(net531),
    .B1(net1565),
    .B2(net804),
    .X(\t$4554 ));
 sky130_fd_sc_hd__xor2_1 \U$$2900  (.A(\t$5887 ),
    .B(net1372),
    .X(booth_b42_m8));
 sky130_fd_sc_hd__a22o_1 \U$$2901  (.A1(net1509),
    .A2(net523),
    .B1(net1500),
    .B2(net796),
    .X(\t$5888 ));
 sky130_fd_sc_hd__xor2_1 \U$$2902  (.A(\t$5888 ),
    .B(net1372),
    .X(booth_b42_m9));
 sky130_fd_sc_hd__a22o_1 \U$$2903  (.A1(net1500),
    .A2(net523),
    .B1(net1225),
    .B2(net796),
    .X(\t$5889 ));
 sky130_fd_sc_hd__xor2_1 \U$$2904  (.A(\t$5889 ),
    .B(net1372),
    .X(booth_b42_m10));
 sky130_fd_sc_hd__a22o_1 \U$$2905  (.A1(net1225),
    .A2(net523),
    .B1(net1218),
    .B2(net796),
    .X(\t$5890 ));
 sky130_fd_sc_hd__xor2_1 \U$$2906  (.A(\t$5890 ),
    .B(net1372),
    .X(booth_b42_m11));
 sky130_fd_sc_hd__a22o_1 \U$$2907  (.A1(net1217),
    .A2(net523),
    .B1(net1207),
    .B2(net796),
    .X(\t$5891 ));
 sky130_fd_sc_hd__xor2_1 \U$$2908  (.A(\t$5891 ),
    .B(net1372),
    .X(booth_b42_m12));
 sky130_fd_sc_hd__a22o_1 \U$$2909  (.A1(net1208),
    .A2(net523),
    .B1(net1200),
    .B2(net796),
    .X(\t$5892 ));
 sky130_fd_sc_hd__xor2_1 \U$$291  (.A(\t$4554 ),
    .B(net1277),
    .X(booth_b4_m5));
 sky130_fd_sc_hd__xor2_1 \U$$2910  (.A(\t$5892 ),
    .B(net1372),
    .X(booth_b42_m13));
 sky130_fd_sc_hd__a22o_1 \U$$2911  (.A1(net1200),
    .A2(net523),
    .B1(net1181),
    .B2(net796),
    .X(\t$5893 ));
 sky130_fd_sc_hd__xor2_1 \U$$2912  (.A(\t$5893 ),
    .B(net1372),
    .X(booth_b42_m14));
 sky130_fd_sc_hd__a22o_1 \U$$2913  (.A1(net1179),
    .A2(net526),
    .B1(net1170),
    .B2(net799),
    .X(\t$5894 ));
 sky130_fd_sc_hd__xor2_1 \U$$2914  (.A(\t$5894 ),
    .B(net1375),
    .X(booth_b42_m15));
 sky130_fd_sc_hd__a22o_1 \U$$2915  (.A1(net1168),
    .A2(net520),
    .B1(net1159),
    .B2(net793),
    .X(\t$5895 ));
 sky130_fd_sc_hd__xor2_1 \U$$2916  (.A(\t$5895 ),
    .B(net1368),
    .X(booth_b42_m16));
 sky130_fd_sc_hd__a22o_1 \U$$2917  (.A1(net1158),
    .A2(net520),
    .B1(net1148),
    .B2(net793),
    .X(\t$5896 ));
 sky130_fd_sc_hd__xor2_1 \U$$2918  (.A(\t$5896 ),
    .B(net1368),
    .X(booth_b42_m17));
 sky130_fd_sc_hd__a22o_1 \U$$2919  (.A1(net1151),
    .A2(net519),
    .B1(net1140),
    .B2(net792),
    .X(\t$5897 ));
 sky130_fd_sc_hd__a22o_1 \U$$292  (.A1(net1564),
    .A2(net531),
    .B1(net1523),
    .B2(net804),
    .X(\t$4555 ));
 sky130_fd_sc_hd__xor2_1 \U$$2920  (.A(\t$5897 ),
    .B(net1367),
    .X(booth_b42_m18));
 sky130_fd_sc_hd__a22o_1 \U$$2921  (.A1(net1141),
    .A2(net520),
    .B1(net1136),
    .B2(net793),
    .X(\t$5898 ));
 sky130_fd_sc_hd__xor2_1 \U$$2922  (.A(\t$5898 ),
    .B(net1368),
    .X(booth_b42_m19));
 sky130_fd_sc_hd__a22o_1 \U$$2923  (.A1(net1136),
    .A2(net520),
    .B1(net1120),
    .B2(net793),
    .X(\t$5899 ));
 sky130_fd_sc_hd__xor2_1 \U$$2924  (.A(\t$5899 ),
    .B(net1368),
    .X(booth_b42_m20));
 sky130_fd_sc_hd__a22o_1 \U$$2925  (.A1(net1120),
    .A2(net522),
    .B1(net1111),
    .B2(net795),
    .X(\t$5900 ));
 sky130_fd_sc_hd__xor2_1 \U$$2926  (.A(\t$5900 ),
    .B(net1371),
    .X(booth_b42_m21));
 sky130_fd_sc_hd__a22o_1 \U$$2927  (.A1(net1109),
    .A2(net523),
    .B1(net1101),
    .B2(net796),
    .X(\t$5901 ));
 sky130_fd_sc_hd__xor2_1 \U$$2928  (.A(\t$5901 ),
    .B(net1372),
    .X(booth_b42_m22));
 sky130_fd_sc_hd__a22o_1 \U$$2929  (.A1(net1104),
    .A2(net523),
    .B1(net1092),
    .B2(net796),
    .X(\t$5902 ));
 sky130_fd_sc_hd__xor2_1 \U$$293  (.A(\t$4555 ),
    .B(net1277),
    .X(booth_b4_m6));
 sky130_fd_sc_hd__xor2_1 \U$$2930  (.A(\t$5902 ),
    .B(net1372),
    .X(booth_b42_m23));
 sky130_fd_sc_hd__a22o_1 \U$$2931  (.A1(net1096),
    .A2(net526),
    .B1(net1087),
    .B2(net799),
    .X(\t$5903 ));
 sky130_fd_sc_hd__xor2_1 \U$$2932  (.A(\t$5903 ),
    .B(net1372),
    .X(booth_b42_m24));
 sky130_fd_sc_hd__a22o_1 \U$$2933  (.A1(net1087),
    .A2(net526),
    .B1(net1078),
    .B2(net799),
    .X(\t$5904 ));
 sky130_fd_sc_hd__xor2_1 \U$$2934  (.A(\t$5904 ),
    .B(net1375),
    .X(booth_b42_m25));
 sky130_fd_sc_hd__a22o_1 \U$$2935  (.A1(net1078),
    .A2(net524),
    .B1(net1070),
    .B2(net797),
    .X(\t$5905 ));
 sky130_fd_sc_hd__xor2_1 \U$$2936  (.A(\t$5905 ),
    .B(net1373),
    .X(booth_b42_m26));
 sky130_fd_sc_hd__a22o_1 \U$$2937  (.A1(net1070),
    .A2(net522),
    .B1(net1062),
    .B2(net795),
    .X(\t$5906 ));
 sky130_fd_sc_hd__xor2_1 \U$$2938  (.A(\t$5906 ),
    .B(net1371),
    .X(booth_b42_m27));
 sky130_fd_sc_hd__a22o_1 \U$$2939  (.A1(net1060),
    .A2(net522),
    .B1(net1051),
    .B2(net795),
    .X(\t$5907 ));
 sky130_fd_sc_hd__a22o_1 \U$$294  (.A1(net1523),
    .A2(net531),
    .B1(net1515),
    .B2(net804),
    .X(\t$4556 ));
 sky130_fd_sc_hd__xor2_1 \U$$2940  (.A(\t$5907 ),
    .B(net1371),
    .X(booth_b42_m28));
 sky130_fd_sc_hd__a22o_1 \U$$2941  (.A1(net1051),
    .A2(net520),
    .B1(net1043),
    .B2(net793),
    .X(\t$5908 ));
 sky130_fd_sc_hd__xor2_1 \U$$2942  (.A(\t$5908 ),
    .B(net1368),
    .X(booth_b42_m29));
 sky130_fd_sc_hd__a22o_1 \U$$2943  (.A1(net1040),
    .A2(net519),
    .B1(net1024),
    .B2(net792),
    .X(\t$5909 ));
 sky130_fd_sc_hd__xor2_1 \U$$2944  (.A(\t$5909 ),
    .B(net1367),
    .X(booth_b42_m30));
 sky130_fd_sc_hd__a22o_1 \U$$2945  (.A1(net1024),
    .A2(net519),
    .B1(net1016),
    .B2(net792),
    .X(\t$5910 ));
 sky130_fd_sc_hd__xor2_1 \U$$2946  (.A(\t$5910 ),
    .B(net1367),
    .X(booth_b42_m31));
 sky130_fd_sc_hd__a22o_1 \U$$2947  (.A1(net1022),
    .A2(net519),
    .B1(net1005),
    .B2(net792),
    .X(\t$5911 ));
 sky130_fd_sc_hd__xor2_1 \U$$2948  (.A(\t$5911 ),
    .B(net1368),
    .X(booth_b42_m32));
 sky130_fd_sc_hd__a22o_1 \U$$2949  (.A1(net1002),
    .A2(net521),
    .B1(net994),
    .B2(net794),
    .X(\t$5912 ));
 sky130_fd_sc_hd__xor2_1 \U$$295  (.A(\t$4556 ),
    .B(net1277),
    .X(booth_b4_m7));
 sky130_fd_sc_hd__xor2_1 \U$$2950  (.A(\t$5912 ),
    .B(net1370),
    .X(booth_b42_m33));
 sky130_fd_sc_hd__a22o_1 \U$$2951  (.A1(net994),
    .A2(net521),
    .B1(net984),
    .B2(net794),
    .X(\t$5913 ));
 sky130_fd_sc_hd__xor2_1 \U$$2952  (.A(\t$5913 ),
    .B(net1370),
    .X(booth_b42_m34));
 sky130_fd_sc_hd__a22o_1 \U$$2953  (.A1(net985),
    .A2(net520),
    .B1(net976),
    .B2(net793),
    .X(\t$5914 ));
 sky130_fd_sc_hd__xor2_1 \U$$2954  (.A(\t$5914 ),
    .B(net1368),
    .X(booth_b42_m35));
 sky130_fd_sc_hd__a22o_1 \U$$2955  (.A1(net975),
    .A2(net521),
    .B1(net966),
    .B2(net794),
    .X(\t$5915 ));
 sky130_fd_sc_hd__xor2_1 \U$$2956  (.A(\t$5915 ),
    .B(net1370),
    .X(booth_b42_m36));
 sky130_fd_sc_hd__a22o_1 \U$$2957  (.A1(net966),
    .A2(net521),
    .B1(net959),
    .B2(net794),
    .X(\t$5916 ));
 sky130_fd_sc_hd__xor2_1 \U$$2958  (.A(\t$5916 ),
    .B(net1370),
    .X(booth_b42_m37));
 sky130_fd_sc_hd__a22o_1 \U$$2959  (.A1(net958),
    .A2(net522),
    .B1(net951),
    .B2(net795),
    .X(\t$5917 ));
 sky130_fd_sc_hd__a22o_1 \U$$296  (.A1(net1516),
    .A2(net531),
    .B1(net1509),
    .B2(net804),
    .X(\t$4557 ));
 sky130_fd_sc_hd__xor2_1 \U$$2960  (.A(\t$5917 ),
    .B(net1371),
    .X(booth_b42_m38));
 sky130_fd_sc_hd__a22o_1 \U$$2961  (.A1(net951),
    .A2(net521),
    .B1(net943),
    .B2(net794),
    .X(\t$5918 ));
 sky130_fd_sc_hd__xor2_1 \U$$2962  (.A(\t$5918 ),
    .B(net1369),
    .X(booth_b42_m39));
 sky130_fd_sc_hd__a22o_1 \U$$2963  (.A1(net942),
    .A2(net521),
    .B1(net926),
    .B2(net794),
    .X(\t$5919 ));
 sky130_fd_sc_hd__xor2_1 \U$$2964  (.A(\t$5919 ),
    .B(net1370),
    .X(booth_b42_m40));
 sky130_fd_sc_hd__a22o_1 \U$$2965  (.A1(net926),
    .A2(net522),
    .B1(net1747),
    .B2(net795),
    .X(\t$5920 ));
 sky130_fd_sc_hd__xor2_1 \U$$2966  (.A(\t$5920 ),
    .B(net1369),
    .X(booth_b42_m41));
 sky130_fd_sc_hd__a22o_1 \U$$2967  (.A1(net1747),
    .A2(net521),
    .B1(net1739),
    .B2(net794),
    .X(\t$5921 ));
 sky130_fd_sc_hd__xor2_1 \U$$2968  (.A(\t$5921 ),
    .B(net1369),
    .X(booth_b42_m42));
 sky130_fd_sc_hd__a22o_1 \U$$2969  (.A1(net1740),
    .A2(net521),
    .B1(net1732),
    .B2(net794),
    .X(\t$5922 ));
 sky130_fd_sc_hd__xor2_1 \U$$297  (.A(\t$4557 ),
    .B(net1277),
    .X(booth_b4_m8));
 sky130_fd_sc_hd__xor2_1 \U$$2970  (.A(\t$5922 ),
    .B(net1369),
    .X(booth_b42_m43));
 sky130_fd_sc_hd__a22o_1 \U$$2971  (.A1(net1731),
    .A2(net521),
    .B1(net1722),
    .B2(net794),
    .X(\t$5923 ));
 sky130_fd_sc_hd__xor2_1 \U$$2972  (.A(\t$5923 ),
    .B(net1369),
    .X(booth_b42_m44));
 sky130_fd_sc_hd__a22o_1 \U$$2973  (.A1(net1723),
    .A2(net521),
    .B1(net1714),
    .B2(net794),
    .X(\t$5924 ));
 sky130_fd_sc_hd__xor2_1 \U$$2974  (.A(\t$5924 ),
    .B(net1369),
    .X(booth_b42_m45));
 sky130_fd_sc_hd__a22o_1 \U$$2975  (.A1(net1719),
    .A2(net522),
    .B1(net1710),
    .B2(net795),
    .X(\t$5925 ));
 sky130_fd_sc_hd__xor2_1 \U$$2976  (.A(\t$5925 ),
    .B(net1371),
    .X(booth_b42_m46));
 sky130_fd_sc_hd__a22o_1 \U$$2977  (.A1(net1705),
    .A2(net522),
    .B1(net1697),
    .B2(net795),
    .X(\t$5926 ));
 sky130_fd_sc_hd__xor2_1 \U$$2978  (.A(\t$5926 ),
    .B(net1371),
    .X(booth_b42_m47));
 sky130_fd_sc_hd__a22o_1 \U$$2979  (.A1(net1697),
    .A2(net522),
    .B1(net1689),
    .B2(net795),
    .X(\t$5927 ));
 sky130_fd_sc_hd__a22o_1 \U$$298  (.A1(net1509),
    .A2(net531),
    .B1(net1500),
    .B2(net804),
    .X(\t$4558 ));
 sky130_fd_sc_hd__xor2_1 \U$$2980  (.A(\t$5927 ),
    .B(net1371),
    .X(booth_b42_m48));
 sky130_fd_sc_hd__a22o_1 \U$$2981  (.A1(net1692),
    .A2(net525),
    .B1(net1685),
    .B2(net798),
    .X(\t$5928 ));
 sky130_fd_sc_hd__xor2_1 \U$$2982  (.A(\t$5928 ),
    .B(net1374),
    .X(booth_b42_m49));
 sky130_fd_sc_hd__a22o_1 \U$$2983  (.A1(net1684),
    .A2(net524),
    .B1(net1660),
    .B2(net797),
    .X(\t$5929 ));
 sky130_fd_sc_hd__xor2_1 \U$$2984  (.A(\t$5929 ),
    .B(net1373),
    .X(booth_b42_m50));
 sky130_fd_sc_hd__a22o_1 \U$$2985  (.A1(net1660),
    .A2(net524),
    .B1(net1652),
    .B2(net797),
    .X(\t$5930 ));
 sky130_fd_sc_hd__xor2_1 \U$$2986  (.A(\t$5930 ),
    .B(net1373),
    .X(booth_b42_m51));
 sky130_fd_sc_hd__a22o_1 \U$$2987  (.A1(net1652),
    .A2(net524),
    .B1(net1644),
    .B2(net797),
    .X(\t$5931 ));
 sky130_fd_sc_hd__xor2_1 \U$$2988  (.A(\t$5931 ),
    .B(net1373),
    .X(booth_b42_m52));
 sky130_fd_sc_hd__a22o_1 \U$$2989  (.A1(net1642),
    .A2(net523),
    .B1(net1637),
    .B2(net796),
    .X(\t$5932 ));
 sky130_fd_sc_hd__xor2_1 \U$$299  (.A(\t$4558 ),
    .B(net1278),
    .X(booth_b4_m9));
 sky130_fd_sc_hd__xor2_1 \U$$2990  (.A(\t$5932 ),
    .B(net1375),
    .X(booth_b42_m53));
 sky130_fd_sc_hd__a22o_1 \U$$2991  (.A1(net1637),
    .A2(net524),
    .B1(net1627),
    .B2(net797),
    .X(\t$5933 ));
 sky130_fd_sc_hd__xor2_1 \U$$2992  (.A(\t$5933 ),
    .B(net1373),
    .X(booth_b42_m54));
 sky130_fd_sc_hd__a22o_1 \U$$2993  (.A1(net1626),
    .A2(net524),
    .B1(net1618),
    .B2(net797),
    .X(\t$5934 ));
 sky130_fd_sc_hd__xor2_1 \U$$2994  (.A(\t$5934 ),
    .B(net1373),
    .X(booth_b42_m55));
 sky130_fd_sc_hd__a22o_1 \U$$2995  (.A1(net1618),
    .A2(net524),
    .B1(net1609),
    .B2(net797),
    .X(\t$5935 ));
 sky130_fd_sc_hd__xor2_1 \U$$2996  (.A(\t$5935 ),
    .B(net1373),
    .X(booth_b42_m56));
 sky130_fd_sc_hd__a22o_1 \U$$2997  (.A1(net1609),
    .A2(net525),
    .B1(net1602),
    .B2(net798),
    .X(\t$5936 ));
 sky130_fd_sc_hd__xor2_1 \U$$2998  (.A(\t$5936 ),
    .B(net1373),
    .X(booth_b42_m57));
 sky130_fd_sc_hd__a22o_1 \U$$2999  (.A1(net1602),
    .A2(net524),
    .B1(net1592),
    .B2(net797),
    .X(\t$5937 ));
 sky130_fd_sc_hd__and2_1 \U$$3  (.A(net1571),
    .B(\notblock[1] ),
    .X(t));
 sky130_fd_sc_hd__a22o_1 \U$$30  (.A1(net1218),
    .A2(net446),
    .B1(net1207),
    .B2(net688),
    .X(\t$4422 ));
 sky130_fd_sc_hd__a22o_1 \U$$300  (.A1(net1496),
    .A2(net532),
    .B1(net1221),
    .B2(net805),
    .X(\t$4559 ));
 sky130_fd_sc_hd__xor2_1 \U$$3000  (.A(\t$5937 ),
    .B(net1373),
    .X(booth_b42_m58));
 sky130_fd_sc_hd__a22o_1 \U$$3001  (.A1(net1592),
    .A2(net525),
    .B1(net1584),
    .B2(net798),
    .X(\t$5938 ));
 sky130_fd_sc_hd__xor2_1 \U$$3002  (.A(\t$5938 ),
    .B(net1373),
    .X(booth_b42_m59));
 sky130_fd_sc_hd__a22o_1 \U$$3003  (.A1(net1585),
    .A2(net524),
    .B1(net1558),
    .B2(net797),
    .X(\t$5939 ));
 sky130_fd_sc_hd__xor2_1 \U$$3004  (.A(\t$5939 ),
    .B(net1374),
    .X(booth_b42_m60));
 sky130_fd_sc_hd__a22o_1 \U$$3005  (.A1(net1556),
    .A2(net525),
    .B1(net1548),
    .B2(net798),
    .X(\t$5940 ));
 sky130_fd_sc_hd__xor2_1 \U$$3006  (.A(\t$5940 ),
    .B(net1374),
    .X(booth_b42_m61));
 sky130_fd_sc_hd__a22o_1 \U$$3007  (.A1(net1548),
    .A2(net525),
    .B1(net1540),
    .B2(net798),
    .X(\t$5941 ));
 sky130_fd_sc_hd__xor2_1 \U$$3008  (.A(\t$5941 ),
    .B(net1374),
    .X(booth_b42_m62));
 sky130_fd_sc_hd__a22o_1 \U$$3009  (.A1(net1542),
    .A2(net524),
    .B1(net1534),
    .B2(net797),
    .X(\t$5942 ));
 sky130_fd_sc_hd__xor2_1 \U$$301  (.A(\t$4559 ),
    .B(net1279),
    .X(booth_b4_m10));
 sky130_fd_sc_hd__xor2_1 \U$$3010  (.A(\t$5942 ),
    .B(net1374),
    .X(booth_b42_m63));
 sky130_fd_sc_hd__a22o_1 \U$$3011  (.A1(net1532),
    .A2(net525),
    .B1(net1786),
    .B2(net798),
    .X(\t$5943 ));
 sky130_fd_sc_hd__xor2_1 \U$$3012  (.A(\t$5943 ),
    .B(net1374),
    .X(booth_b42_m64));
 sky130_fd_sc_hd__inv_1 \U$$3013  (.A(net1374),
    .Y(\notsign$5944 ));
 sky130_fd_sc_hd__inv_1 \U$$3014  (.A(net1369),
    .Y(\notblock$5945[0] ));
 sky130_fd_sc_hd__inv_1 \U$$3015  (.A(net39),
    .Y(\notblock$5945[1] ));
 sky130_fd_sc_hd__inv_1 \U$$3016  (.A(net1359),
    .Y(\notblock$5945[2] ));
 sky130_fd_sc_hd__and2_1 \U$$3017  (.A(net1359),
    .B(\notblock$5945[1] ),
    .X(\t$5946 ));
 sky130_fd_sc_hd__a32o_1 \U$$3018  (.A1(\notblock$5945[2] ),
    .A2(net39),
    .A3(net1369),
    .B1(\t$5946 ),
    .B2(\notblock$5945[0] ),
    .X(\sel_0$5947 ));
 sky130_fd_sc_hd__xor2_1 \U$$3019  (.A(net39),
    .B(net1370),
    .X(\sel_1$5948 ));
 sky130_fd_sc_hd__a22o_1 \U$$302  (.A1(net1221),
    .A2(net532),
    .B1(net1211),
    .B2(net805),
    .X(\t$4560 ));
 sky130_fd_sc_hd__a22o_1 \U$$3020  (.A1(net1787),
    .A2(net510),
    .B1(net1229),
    .B2(net783),
    .X(\t$5949 ));
 sky130_fd_sc_hd__xor2_1 \U$$3021  (.A(\t$5949 ),
    .B(net1357),
    .X(booth_b44_m0));
 sky130_fd_sc_hd__a22o_1 \U$$3022  (.A1(net1228),
    .A2(net511),
    .B1(net1124),
    .B2(net784),
    .X(\t$5950 ));
 sky130_fd_sc_hd__xor2_1 \U$$3023  (.A(\t$5950 ),
    .B(net1358),
    .X(booth_b44_m1));
 sky130_fd_sc_hd__a22o_1 \U$$3024  (.A1(net1125),
    .A2(net511),
    .B1(net1034),
    .B2(net784),
    .X(\t$5951 ));
 sky130_fd_sc_hd__xor2_1 \U$$3025  (.A(\t$5951 ),
    .B(net1358),
    .X(booth_b44_m2));
 sky130_fd_sc_hd__a22o_1 \U$$3026  (.A1(net1034),
    .A2(net510),
    .B1(net935),
    .B2(net783),
    .X(\t$5952 ));
 sky130_fd_sc_hd__xor2_1 \U$$3027  (.A(\t$5952 ),
    .B(net1357),
    .X(booth_b44_m3));
 sky130_fd_sc_hd__a22o_1 \U$$3028  (.A1(net935),
    .A2(net510),
    .B1(net1673),
    .B2(net783),
    .X(\t$5953 ));
 sky130_fd_sc_hd__xor2_1 \U$$3029  (.A(\t$5953 ),
    .B(net1357),
    .X(booth_b44_m4));
 sky130_fd_sc_hd__xor2_1 \U$$303  (.A(\t$4560 ),
    .B(net1279),
    .X(booth_b4_m11));
 sky130_fd_sc_hd__a22o_1 \U$$3030  (.A1(net1674),
    .A2(net510),
    .B1(net1563),
    .B2(net783),
    .X(\t$5954 ));
 sky130_fd_sc_hd__xor2_1 \U$$3031  (.A(\t$5954 ),
    .B(net1357),
    .X(booth_b44_m5));
 sky130_fd_sc_hd__a22o_1 \U$$3032  (.A1(net1565),
    .A2(net514),
    .B1(net1524),
    .B2(net787),
    .X(\t$5955 ));
 sky130_fd_sc_hd__xor2_1 \U$$3033  (.A(\t$5955 ),
    .B(net1362),
    .X(booth_b44_m6));
 sky130_fd_sc_hd__a22o_1 \U$$3034  (.A1(net1524),
    .A2(net514),
    .B1(net1516),
    .B2(net787),
    .X(\t$5956 ));
 sky130_fd_sc_hd__xor2_1 \U$$3035  (.A(\t$5956 ),
    .B(net1362),
    .X(booth_b44_m7));
 sky130_fd_sc_hd__a22o_1 \U$$3036  (.A1(net1516),
    .A2(net514),
    .B1(net1509),
    .B2(net787),
    .X(\t$5957 ));
 sky130_fd_sc_hd__xor2_1 \U$$3037  (.A(\t$5957 ),
    .B(net1362),
    .X(booth_b44_m8));
 sky130_fd_sc_hd__a22o_1 \U$$3038  (.A1(net1509),
    .A2(net514),
    .B1(net1500),
    .B2(net787),
    .X(\t$5958 ));
 sky130_fd_sc_hd__xor2_1 \U$$3039  (.A(\t$5958 ),
    .B(net1362),
    .X(booth_b44_m9));
 sky130_fd_sc_hd__a22o_1 \U$$304  (.A1(net1211),
    .A2(net528),
    .B1(net1203),
    .B2(net801),
    .X(\t$4561 ));
 sky130_fd_sc_hd__a22o_1 \U$$3040  (.A1(net1501),
    .A2(net514),
    .B1(net1226),
    .B2(net787),
    .X(\t$5959 ));
 sky130_fd_sc_hd__xor2_1 \U$$3041  (.A(\t$5959 ),
    .B(net1362),
    .X(booth_b44_m10));
 sky130_fd_sc_hd__a22o_1 \U$$3042  (.A1(net1226),
    .A2(net514),
    .B1(net1217),
    .B2(net787),
    .X(\t$5960 ));
 sky130_fd_sc_hd__xor2_1 \U$$3043  (.A(\t$5960 ),
    .B(net1362),
    .X(booth_b44_m11));
 sky130_fd_sc_hd__a22o_1 \U$$3044  (.A1(net1217),
    .A2(net514),
    .B1(net1208),
    .B2(net787),
    .X(\t$5961 ));
 sky130_fd_sc_hd__xor2_1 \U$$3045  (.A(\t$5961 ),
    .B(net1362),
    .X(booth_b44_m12));
 sky130_fd_sc_hd__a22o_1 \U$$3046  (.A1(net1206),
    .A2(net517),
    .B1(net1198),
    .B2(net790),
    .X(\t$5962 ));
 sky130_fd_sc_hd__xor2_1 \U$$3047  (.A(\t$5962 ),
    .B(net1363),
    .X(booth_b44_m13));
 sky130_fd_sc_hd__a22o_1 \U$$3048  (.A1(net1196),
    .A2(net511),
    .B1(net1178),
    .B2(net784),
    .X(\t$5963 ));
 sky130_fd_sc_hd__xor2_1 \U$$3049  (.A(\t$5963 ),
    .B(net1358),
    .X(booth_b44_m14));
 sky130_fd_sc_hd__xor2_1 \U$$305  (.A(\t$4561 ),
    .B(net1274),
    .X(booth_b4_m12));
 sky130_fd_sc_hd__a22o_1 \U$$3050  (.A1(net1176),
    .A2(net511),
    .B1(net1167),
    .B2(net784),
    .X(\t$5964 ));
 sky130_fd_sc_hd__xor2_1 \U$$3051  (.A(\t$5964 ),
    .B(net1358),
    .X(booth_b44_m15));
 sky130_fd_sc_hd__a22o_1 \U$$3052  (.A1(net1165),
    .A2(net510),
    .B1(net1156),
    .B2(net783),
    .X(\t$5965 ));
 sky130_fd_sc_hd__xor2_1 \U$$3053  (.A(\t$5965 ),
    .B(net1357),
    .X(booth_b44_m16));
 sky130_fd_sc_hd__a22o_1 \U$$3054  (.A1(net1159),
    .A2(net510),
    .B1(net1151),
    .B2(net783),
    .X(\t$5966 ));
 sky130_fd_sc_hd__xor2_1 \U$$3055  (.A(\t$5966 ),
    .B(net1358),
    .X(booth_b44_m17));
 sky130_fd_sc_hd__a22o_1 \U$$3056  (.A1(net1151),
    .A2(net511),
    .B1(net1142),
    .B2(net784),
    .X(\t$5967 ));
 sky130_fd_sc_hd__xor2_1 \U$$3057  (.A(\t$5967 ),
    .B(net1358),
    .X(booth_b44_m18));
 sky130_fd_sc_hd__a22o_1 \U$$3058  (.A1(net1142),
    .A2(net513),
    .B1(net1135),
    .B2(net786),
    .X(\t$5968 ));
 sky130_fd_sc_hd__xor2_1 \U$$3059  (.A(\t$5968 ),
    .B(net1360),
    .X(booth_b44_m19));
 sky130_fd_sc_hd__a22o_1 \U$$306  (.A1(net1203),
    .A2(net528),
    .B1(net1194),
    .B2(net801),
    .X(\t$4562 ));
 sky130_fd_sc_hd__a22o_1 \U$$3060  (.A1(net1137),
    .A2(net514),
    .B1(net1121),
    .B2(net787),
    .X(\t$5969 ));
 sky130_fd_sc_hd__xor2_1 \U$$3061  (.A(\t$5969 ),
    .B(net1362),
    .X(booth_b44_m20));
 sky130_fd_sc_hd__a22o_1 \U$$3062  (.A1(net1121),
    .A2(net514),
    .B1(net1113),
    .B2(net787),
    .X(\t$5970 ));
 sky130_fd_sc_hd__xor2_1 \U$$3063  (.A(\t$5970 ),
    .B(net1362),
    .X(booth_b44_m21));
 sky130_fd_sc_hd__a22o_1 \U$$3064  (.A1(net1113),
    .A2(net517),
    .B1(net1104),
    .B2(net790),
    .X(\t$5971 ));
 sky130_fd_sc_hd__xor2_1 \U$$3065  (.A(\t$5971 ),
    .B(net1362),
    .X(booth_b44_m22));
 sky130_fd_sc_hd__a22o_1 \U$$3066  (.A1(net1104),
    .A2(net517),
    .B1(net1096),
    .B2(net790),
    .X(\t$5972 ));
 sky130_fd_sc_hd__xor2_1 \U$$3067  (.A(\t$5972 ),
    .B(net1363),
    .X(booth_b44_m23));
 sky130_fd_sc_hd__a22o_1 \U$$3068  (.A1(net1096),
    .A2(net515),
    .B1(net1087),
    .B2(net788),
    .X(\t$5973 ));
 sky130_fd_sc_hd__xor2_1 \U$$3069  (.A(\t$5973 ),
    .B(net1363),
    .X(booth_b44_m24));
 sky130_fd_sc_hd__xor2_1 \U$$307  (.A(\t$4562 ),
    .B(net1274),
    .X(booth_b4_m13));
 sky130_fd_sc_hd__a22o_1 \U$$3070  (.A1(net1087),
    .A2(net511),
    .B1(net1078),
    .B2(net784),
    .X(\t$5974 ));
 sky130_fd_sc_hd__xor2_1 \U$$3071  (.A(\t$5974 ),
    .B(net1358),
    .X(booth_b44_m25));
 sky130_fd_sc_hd__a22o_1 \U$$3072  (.A1(net1076),
    .A2(net513),
    .B1(net1068),
    .B2(net786),
    .X(\t$5975 ));
 sky130_fd_sc_hd__xor2_1 \U$$3073  (.A(\t$5975 ),
    .B(net1360),
    .X(booth_b44_m26));
 sky130_fd_sc_hd__a22o_1 \U$$3074  (.A1(net1068),
    .A2(net511),
    .B1(net1060),
    .B2(net784),
    .X(\t$5976 ));
 sky130_fd_sc_hd__xor2_1 \U$$3075  (.A(\t$5976 ),
    .B(net1358),
    .X(booth_b44_m27));
 sky130_fd_sc_hd__a22o_1 \U$$3076  (.A1(net1059),
    .A2(net510),
    .B1(net1048),
    .B2(net783),
    .X(\t$5977 ));
 sky130_fd_sc_hd__xor2_1 \U$$3077  (.A(\t$5977 ),
    .B(net1357),
    .X(booth_b44_m28));
 sky130_fd_sc_hd__a22o_1 \U$$3078  (.A1(net1048),
    .A2(net510),
    .B1(net1040),
    .B2(net783),
    .X(\t$5978 ));
 sky130_fd_sc_hd__xor2_1 \U$$3079  (.A(\t$5978 ),
    .B(net1357),
    .X(booth_b44_m29));
 sky130_fd_sc_hd__a22o_1 \U$$308  (.A1(net1194),
    .A2(net528),
    .B1(net1175),
    .B2(net801),
    .X(\t$4563 ));
 sky130_fd_sc_hd__a22o_1 \U$$3080  (.A1(net1046),
    .A2(net510),
    .B1(net1030),
    .B2(net783),
    .X(\t$5979 ));
 sky130_fd_sc_hd__xor2_1 \U$$3081  (.A(\t$5979 ),
    .B(net1357),
    .X(booth_b44_m30));
 sky130_fd_sc_hd__a22o_1 \U$$3082  (.A1(net1027),
    .A2(net512),
    .B1(net1019),
    .B2(net785),
    .X(\t$5980 ));
 sky130_fd_sc_hd__xor2_1 \U$$3083  (.A(\t$5980 ),
    .B(net1359),
    .X(booth_b44_m31));
 sky130_fd_sc_hd__a22o_1 \U$$3084  (.A1(net1019),
    .A2(net512),
    .B1(net1002),
    .B2(net785),
    .X(\t$5981 ));
 sky130_fd_sc_hd__xor2_1 \U$$3085  (.A(\t$5981 ),
    .B(net1359),
    .X(booth_b44_m32));
 sky130_fd_sc_hd__a22o_1 \U$$3086  (.A1(net1002),
    .A2(net510),
    .B1(net994),
    .B2(net783),
    .X(\t$5982 ));
 sky130_fd_sc_hd__xor2_1 \U$$3087  (.A(\t$5982 ),
    .B(net1357),
    .X(booth_b44_m33));
 sky130_fd_sc_hd__a22o_1 \U$$3088  (.A1(net994),
    .A2(net512),
    .B1(net985),
    .B2(net785),
    .X(\t$5983 ));
 sky130_fd_sc_hd__xor2_1 \U$$3089  (.A(\t$5983 ),
    .B(net1359),
    .X(booth_b44_m34));
 sky130_fd_sc_hd__xor2_1 \U$$309  (.A(\t$4563 ),
    .B(net1274),
    .X(booth_b4_m14));
 sky130_fd_sc_hd__a22o_1 \U$$3090  (.A1(net985),
    .A2(net513),
    .B1(net976),
    .B2(net786),
    .X(\t$5984 ));
 sky130_fd_sc_hd__xor2_1 \U$$3091  (.A(\t$5984 ),
    .B(net1360),
    .X(booth_b44_m35));
 sky130_fd_sc_hd__a22o_1 \U$$3092  (.A1(net976),
    .A2(net513),
    .B1(net967),
    .B2(net786),
    .X(\t$5985 ));
 sky130_fd_sc_hd__xor2_1 \U$$3093  (.A(\t$5985 ),
    .B(net1360),
    .X(booth_b44_m36));
 sky130_fd_sc_hd__a22o_1 \U$$3094  (.A1(net967),
    .A2(net512),
    .B1(net958),
    .B2(net785),
    .X(\t$5986 ));
 sky130_fd_sc_hd__xor2_1 \U$$3095  (.A(\t$5986 ),
    .B(net1359),
    .X(booth_b44_m37));
 sky130_fd_sc_hd__a22o_1 \U$$3096  (.A1(net959),
    .A2(net512),
    .B1(net950),
    .B2(net785),
    .X(\t$5987 ));
 sky130_fd_sc_hd__xor2_1 \U$$3097  (.A(\t$5987 ),
    .B(net1359),
    .X(booth_b44_m38));
 sky130_fd_sc_hd__a22o_1 \U$$3098  (.A1(net950),
    .A2(net512),
    .B1(net942),
    .B2(net785),
    .X(\t$5988 ));
 sky130_fd_sc_hd__xor2_1 \U$$3099  (.A(\t$5988 ),
    .B(net1359),
    .X(booth_b44_m39));
 sky130_fd_sc_hd__xor2_1 \U$$31  (.A(\t$4422 ),
    .B(net1573),
    .X(booth_b0_m12));
 sky130_fd_sc_hd__a22o_1 \U$$310  (.A1(net1179),
    .A2(net532),
    .B1(net1166),
    .B2(net805),
    .X(\t$4564 ));
 sky130_fd_sc_hd__a22o_1 \U$$3100  (.A1(net942),
    .A2(net512),
    .B1(net926),
    .B2(net785),
    .X(\t$5989 ));
 sky130_fd_sc_hd__xor2_1 \U$$3101  (.A(\t$5989 ),
    .B(net1359),
    .X(booth_b44_m40));
 sky130_fd_sc_hd__a22o_1 \U$$3102  (.A1(net926),
    .A2(net512),
    .B1(net1747),
    .B2(net785),
    .X(\t$5990 ));
 sky130_fd_sc_hd__xor2_1 \U$$3103  (.A(\t$5990 ),
    .B(net1359),
    .X(booth_b44_m41));
 sky130_fd_sc_hd__a22o_1 \U$$3104  (.A1(net1747),
    .A2(net512),
    .B1(net1739),
    .B2(net785),
    .X(\t$5991 ));
 sky130_fd_sc_hd__xor2_1 \U$$3105  (.A(\t$5991 ),
    .B(net1361),
    .X(booth_b44_m42));
 sky130_fd_sc_hd__a22o_1 \U$$3106  (.A1(net1740),
    .A2(net512),
    .B1(net1732),
    .B2(net785),
    .X(\t$5992 ));
 sky130_fd_sc_hd__xor2_1 \U$$3107  (.A(\t$5992 ),
    .B(net1361),
    .X(booth_b44_m43));
 sky130_fd_sc_hd__a22o_1 \U$$3108  (.A1(net1735),
    .A2(net513),
    .B1(net1727),
    .B2(net786),
    .X(\t$5993 ));
 sky130_fd_sc_hd__xor2_1 \U$$3109  (.A(\t$5993 ),
    .B(net1360),
    .X(booth_b44_m44));
 sky130_fd_sc_hd__xor2_1 \U$$311  (.A(\t$4564 ),
    .B(net1279),
    .X(booth_b4_m15));
 sky130_fd_sc_hd__a22o_1 \U$$3110  (.A1(net1723),
    .A2(net513),
    .B1(net1714),
    .B2(net786),
    .X(\t$5994 ));
 sky130_fd_sc_hd__xor2_1 \U$$3111  (.A(\t$5994 ),
    .B(net1360),
    .X(booth_b44_m45));
 sky130_fd_sc_hd__a22o_1 \U$$3112  (.A1(net1714),
    .A2(net513),
    .B1(net1705),
    .B2(net786),
    .X(\t$5995 ));
 sky130_fd_sc_hd__xor2_1 \U$$3113  (.A(\t$5995 ),
    .B(net1360),
    .X(booth_b44_m46));
 sky130_fd_sc_hd__a22o_1 \U$$3114  (.A1(net1708),
    .A2(net515),
    .B1(net1700),
    .B2(net788),
    .X(\t$5996 ));
 sky130_fd_sc_hd__xor2_1 \U$$3115  (.A(\t$5996 ),
    .B(net1364),
    .X(booth_b44_m47));
 sky130_fd_sc_hd__a22o_1 \U$$3116  (.A1(net1700),
    .A2(net515),
    .B1(net1693),
    .B2(net788),
    .X(\t$5997 ));
 sky130_fd_sc_hd__xor2_1 \U$$3117  (.A(\t$5997 ),
    .B(net1364),
    .X(booth_b44_m48));
 sky130_fd_sc_hd__a22o_1 \U$$3118  (.A1(net1693),
    .A2(net515),
    .B1(net1684),
    .B2(net788),
    .X(\t$5998 ));
 sky130_fd_sc_hd__xor2_1 \U$$3119  (.A(\t$5998 ),
    .B(net1364),
    .X(booth_b44_m49));
 sky130_fd_sc_hd__a22o_1 \U$$312  (.A1(net1170),
    .A2(net532),
    .B1(net1161),
    .B2(net805),
    .X(\t$4565 ));
 sky130_fd_sc_hd__a22o_1 \U$$3120  (.A1(net1684),
    .A2(net515),
    .B1(net1660),
    .B2(net788),
    .X(\t$5999 ));
 sky130_fd_sc_hd__xor2_1 \U$$3121  (.A(\t$5999 ),
    .B(net1364),
    .X(booth_b44_m50));
 sky130_fd_sc_hd__a22o_1 \U$$3122  (.A1(net1658),
    .A2(net514),
    .B1(net1650),
    .B2(net787),
    .X(\t$6000 ));
 sky130_fd_sc_hd__xor2_1 \U$$3123  (.A(\t$6000 ),
    .B(net1363),
    .X(booth_b44_m51));
 sky130_fd_sc_hd__a22o_1 \U$$3124  (.A1(net1650),
    .A2(net515),
    .B1(net1642),
    .B2(net788),
    .X(\t$6001 ));
 sky130_fd_sc_hd__xor2_1 \U$$3125  (.A(\t$6001 ),
    .B(net1364),
    .X(booth_b44_m52));
 sky130_fd_sc_hd__a22o_1 \U$$3126  (.A1(net1644),
    .A2(net515),
    .B1(net1635),
    .B2(net788),
    .X(\t$6002 ));
 sky130_fd_sc_hd__xor2_1 \U$$3127  (.A(\t$6002 ),
    .B(net1364),
    .X(booth_b44_m53));
 sky130_fd_sc_hd__a22o_1 \U$$3128  (.A1(net1635),
    .A2(net516),
    .B1(net1626),
    .B2(net789),
    .X(\t$6003 ));
 sky130_fd_sc_hd__xor2_1 \U$$3129  (.A(\t$6003 ),
    .B(net1364),
    .X(booth_b44_m54));
 sky130_fd_sc_hd__xor2_1 \U$$313  (.A(\t$4565 ),
    .B(net1279),
    .X(booth_b4_m16));
 sky130_fd_sc_hd__a22o_1 \U$$3130  (.A1(net1626),
    .A2(net516),
    .B1(net1618),
    .B2(net789),
    .X(\t$6004 ));
 sky130_fd_sc_hd__xor2_1 \U$$3131  (.A(\t$6004 ),
    .B(net1364),
    .X(booth_b44_m55));
 sky130_fd_sc_hd__a22o_1 \U$$3132  (.A1(net1618),
    .A2(net515),
    .B1(net1609),
    .B2(net788),
    .X(\t$6005 ));
 sky130_fd_sc_hd__xor2_1 \U$$3133  (.A(\t$6005 ),
    .B(net1364),
    .X(booth_b44_m56));
 sky130_fd_sc_hd__a22o_1 \U$$3134  (.A1(net1609),
    .A2(net516),
    .B1(net1602),
    .B2(net789),
    .X(\t$6006 ));
 sky130_fd_sc_hd__xor2_1 \U$$3135  (.A(\t$6006 ),
    .B(net1365),
    .X(booth_b44_m57));
 sky130_fd_sc_hd__a22o_1 \U$$3136  (.A1(net1602),
    .A2(net516),
    .B1(net1593),
    .B2(net789),
    .X(\t$6007 ));
 sky130_fd_sc_hd__xor2_1 \U$$3137  (.A(\t$6007 ),
    .B(net1365),
    .X(booth_b44_m58));
 sky130_fd_sc_hd__a22o_1 \U$$3138  (.A1(net1590),
    .A2(net513),
    .B1(net1582),
    .B2(net786),
    .X(\t$6008 ));
 sky130_fd_sc_hd__xor2_1 \U$$3139  (.A(\t$6008 ),
    .B(net1360),
    .X(booth_b44_m59));
 sky130_fd_sc_hd__a22o_1 \U$$314  (.A1(net1161),
    .A2(net532),
    .B1(net1149),
    .B2(net805),
    .X(\t$4566 ));
 sky130_fd_sc_hd__a22o_1 \U$$3140  (.A1(net1585),
    .A2(net515),
    .B1(net1558),
    .B2(net788),
    .X(\t$6009 ));
 sky130_fd_sc_hd__xor2_1 \U$$3141  (.A(\t$6009 ),
    .B(net1364),
    .X(booth_b44_m60));
 sky130_fd_sc_hd__a22o_1 \U$$3142  (.A1(net1558),
    .A2(net515),
    .B1(net1550),
    .B2(net788),
    .X(\t$6010 ));
 sky130_fd_sc_hd__xor2_1 \U$$3143  (.A(\t$6010 ),
    .B(net1365),
    .X(booth_b44_m61));
 sky130_fd_sc_hd__a22o_1 \U$$3144  (.A1(net1548),
    .A2(net516),
    .B1(net1540),
    .B2(net789),
    .X(\t$6011 ));
 sky130_fd_sc_hd__xor2_1 \U$$3145  (.A(\t$6011 ),
    .B(net1365),
    .X(booth_b44_m62));
 sky130_fd_sc_hd__a22o_1 \U$$3146  (.A1(net1539),
    .A2(net516),
    .B1(net1531),
    .B2(net789),
    .X(\t$6012 ));
 sky130_fd_sc_hd__xor2_1 \U$$3147  (.A(\t$6012 ),
    .B(net1365),
    .X(booth_b44_m63));
 sky130_fd_sc_hd__a22o_1 \U$$3148  (.A1(net1532),
    .A2(net513),
    .B1(net1788),
    .B2(net786),
    .X(\t$6013 ));
 sky130_fd_sc_hd__xor2_1 \U$$3149  (.A(\t$6013 ),
    .B(net1360),
    .X(booth_b44_m64));
 sky130_fd_sc_hd__xor2_1 \U$$315  (.A(\t$4566 ),
    .B(net1279),
    .X(booth_b4_m17));
 sky130_fd_sc_hd__inv_1 \U$$3150  (.A(net1360),
    .Y(\notsign$6014 ));
 sky130_fd_sc_hd__inv_1 \U$$3151  (.A(net1361),
    .Y(\notblock$6015[0] ));
 sky130_fd_sc_hd__inv_1 \U$$3152  (.A(net41),
    .Y(\notblock$6015[1] ));
 sky130_fd_sc_hd__inv_1 \U$$3153  (.A(net1350),
    .Y(\notblock$6015[2] ));
 sky130_fd_sc_hd__and2_1 \U$$3154  (.A(net1350),
    .B(\notblock$6015[1] ),
    .X(\t$6016 ));
 sky130_fd_sc_hd__a32o_1 \U$$3155  (.A1(\notblock$6015[2] ),
    .A2(net41),
    .A3(net1361),
    .B1(\t$6016 ),
    .B2(\notblock$6015[0] ),
    .X(\sel_0$6017 ));
 sky130_fd_sc_hd__xor2_1 \U$$3156  (.A(net41),
    .B(net1361),
    .X(\sel_1$6018 ));
 sky130_fd_sc_hd__a22o_1 \U$$3157  (.A1(net1789),
    .A2(net502),
    .B1(net1229),
    .B2(net775),
    .X(\t$6019 ));
 sky130_fd_sc_hd__xor2_1 \U$$3158  (.A(\t$6019 ),
    .B(net1349),
    .X(booth_b46_m0));
 sky130_fd_sc_hd__a22o_1 \U$$3159  (.A1(net1229),
    .A2(net501),
    .B1(net1125),
    .B2(net774),
    .X(\t$6020 ));
 sky130_fd_sc_hd__a22o_1 \U$$316  (.A1(net1149),
    .A2(net532),
    .B1(net1143),
    .B2(net805),
    .X(\t$4567 ));
 sky130_fd_sc_hd__xor2_1 \U$$3160  (.A(\t$6020 ),
    .B(net1348),
    .X(booth_b46_m1));
 sky130_fd_sc_hd__a22o_1 \U$$3161  (.A1(net1125),
    .A2(net501),
    .B1(net1034),
    .B2(net774),
    .X(\t$6021 ));
 sky130_fd_sc_hd__xor2_1 \U$$3162  (.A(\t$6021 ),
    .B(net1348),
    .X(booth_b46_m2));
 sky130_fd_sc_hd__a22o_1 \U$$3163  (.A1(net1034),
    .A2(net501),
    .B1(net935),
    .B2(net774),
    .X(\t$6022 ));
 sky130_fd_sc_hd__xor2_1 \U$$3164  (.A(\t$6022 ),
    .B(net1348),
    .X(booth_b46_m3));
 sky130_fd_sc_hd__a22o_1 \U$$3165  (.A1(net938),
    .A2(net505),
    .B1(net1677),
    .B2(net778),
    .X(\t$6023 ));
 sky130_fd_sc_hd__xor2_1 \U$$3166  (.A(\t$6023 ),
    .B(net1353),
    .X(booth_b46_m4));
 sky130_fd_sc_hd__a22o_1 \U$$3167  (.A1(net1678),
    .A2(net505),
    .B1(net1567),
    .B2(net778),
    .X(\t$6024 ));
 sky130_fd_sc_hd__xor2_1 \U$$3168  (.A(\t$6024 ),
    .B(net1353),
    .X(booth_b46_m5));
 sky130_fd_sc_hd__a22o_1 \U$$3169  (.A1(net1566),
    .A2(net505),
    .B1(net1526),
    .B2(net778),
    .X(\t$6025 ));
 sky130_fd_sc_hd__xor2_1 \U$$317  (.A(\t$4567 ),
    .B(net1279),
    .X(booth_b4_m18));
 sky130_fd_sc_hd__xor2_1 \U$$3170  (.A(\t$6025 ),
    .B(net1353),
    .X(booth_b46_m6));
 sky130_fd_sc_hd__a22o_1 \U$$3171  (.A1(net1525),
    .A2(net505),
    .B1(net1517),
    .B2(net778),
    .X(\t$6026 ));
 sky130_fd_sc_hd__xor2_1 \U$$3172  (.A(\t$6026 ),
    .B(net1353),
    .X(booth_b46_m7));
 sky130_fd_sc_hd__a22o_1 \U$$3173  (.A1(net1517),
    .A2(net505),
    .B1(net1510),
    .B2(net778),
    .X(\t$6027 ));
 sky130_fd_sc_hd__xor2_1 \U$$3174  (.A(\t$6027 ),
    .B(net1353),
    .X(booth_b46_m8));
 sky130_fd_sc_hd__a22o_1 \U$$3175  (.A1(net1510),
    .A2(net505),
    .B1(net1501),
    .B2(net778),
    .X(\t$6028 ));
 sky130_fd_sc_hd__xor2_1 \U$$3176  (.A(\t$6028 ),
    .B(net1353),
    .X(booth_b46_m9));
 sky130_fd_sc_hd__a22o_1 \U$$3177  (.A1(net1501),
    .A2(net506),
    .B1(net1226),
    .B2(net779),
    .X(\t$6029 ));
 sky130_fd_sc_hd__xor2_1 \U$$3178  (.A(\t$6029 ),
    .B(net1354),
    .X(booth_b46_m10));
 sky130_fd_sc_hd__a22o_1 \U$$3179  (.A1(net1226),
    .A2(net506),
    .B1(net1217),
    .B2(net779),
    .X(\t$6030 ));
 sky130_fd_sc_hd__a22o_1 \U$$318  (.A1(net1143),
    .A2(net532),
    .B1(net1133),
    .B2(net805),
    .X(\t$4568 ));
 sky130_fd_sc_hd__xor2_1 \U$$3180  (.A(\t$6030 ),
    .B(net1354),
    .X(booth_b46_m11));
 sky130_fd_sc_hd__a22o_1 \U$$3181  (.A1(net1212),
    .A2(net502),
    .B1(net1204),
    .B2(net775),
    .X(\t$6031 ));
 sky130_fd_sc_hd__xor2_1 \U$$3182  (.A(\t$6031 ),
    .B(net1349),
    .X(booth_b46_m12));
 sky130_fd_sc_hd__a22o_1 \U$$3183  (.A1(net1202),
    .A2(net501),
    .B1(net1193),
    .B2(net774),
    .X(\t$6032 ));
 sky130_fd_sc_hd__xor2_1 \U$$3184  (.A(\t$6032 ),
    .B(net1348),
    .X(booth_b46_m13));
 sky130_fd_sc_hd__a22o_1 \U$$3185  (.A1(net1193),
    .A2(net501),
    .B1(net1177),
    .B2(net774),
    .X(\t$6033 ));
 sky130_fd_sc_hd__xor2_1 \U$$3186  (.A(\t$6033 ),
    .B(net1348),
    .X(booth_b46_m14));
 sky130_fd_sc_hd__a22o_1 \U$$3187  (.A1(net1177),
    .A2(net501),
    .B1(net1168),
    .B2(net774),
    .X(\t$6034 ));
 sky130_fd_sc_hd__xor2_1 \U$$3188  (.A(\t$6034 ),
    .B(net1348),
    .X(booth_b46_m15));
 sky130_fd_sc_hd__a22o_1 \U$$3189  (.A1(net1168),
    .A2(net502),
    .B1(net1160),
    .B2(net775),
    .X(\t$6035 ));
 sky130_fd_sc_hd__xor2_1 \U$$319  (.A(\t$4568 ),
    .B(net1279),
    .X(booth_b4_m19));
 sky130_fd_sc_hd__xor2_1 \U$$3190  (.A(\t$6035 ),
    .B(net1349),
    .X(booth_b46_m16));
 sky130_fd_sc_hd__a22o_1 \U$$3191  (.A1(net1159),
    .A2(net501),
    .B1(net1151),
    .B2(net774),
    .X(\t$6036 ));
 sky130_fd_sc_hd__xor2_1 \U$$3192  (.A(\t$6036 ),
    .B(net1349),
    .X(booth_b46_m17));
 sky130_fd_sc_hd__a22o_1 \U$$3193  (.A1(net1153),
    .A2(net505),
    .B1(net1145),
    .B2(net778),
    .X(\t$6037 ));
 sky130_fd_sc_hd__xor2_1 \U$$3194  (.A(\t$6037 ),
    .B(net1353),
    .X(booth_b46_m18));
 sky130_fd_sc_hd__a22o_1 \U$$3195  (.A1(net1145),
    .A2(net505),
    .B1(net1137),
    .B2(net778),
    .X(\t$6038 ));
 sky130_fd_sc_hd__xor2_1 \U$$3196  (.A(\t$6038 ),
    .B(net1353),
    .X(booth_b46_m19));
 sky130_fd_sc_hd__a22o_1 \U$$3197  (.A1(net1137),
    .A2(net505),
    .B1(net1121),
    .B2(net778),
    .X(\t$6039 ));
 sky130_fd_sc_hd__xor2_1 \U$$3198  (.A(\t$6039 ),
    .B(net1353),
    .X(booth_b46_m20));
 sky130_fd_sc_hd__a22o_1 \U$$3199  (.A1(net1121),
    .A2(net506),
    .B1(net1113),
    .B2(net779),
    .X(\t$6040 ));
 sky130_fd_sc_hd__a22o_1 \U$$32  (.A1(net1207),
    .A2(net447),
    .B1(net1199),
    .B2(net689),
    .X(\t$4423 ));
 sky130_fd_sc_hd__a22o_1 \U$$320  (.A1(net1131),
    .A2(net528),
    .B1(net1115),
    .B2(net801),
    .X(\t$4569 ));
 sky130_fd_sc_hd__xor2_1 \U$$3200  (.A(\t$6040 ),
    .B(net1353),
    .X(booth_b46_m21));
 sky130_fd_sc_hd__a22o_1 \U$$3201  (.A1(net1113),
    .A2(net506),
    .B1(net1104),
    .B2(net779),
    .X(\t$6041 ));
 sky130_fd_sc_hd__xor2_1 \U$$3202  (.A(\t$6041 ),
    .B(net1354),
    .X(booth_b46_m22));
 sky130_fd_sc_hd__a22o_1 \U$$3203  (.A1(net1104),
    .A2(net506),
    .B1(net1096),
    .B2(net779),
    .X(\t$6042 ));
 sky130_fd_sc_hd__xor2_1 \U$$3204  (.A(\t$6042 ),
    .B(net1354),
    .X(booth_b46_m23));
 sky130_fd_sc_hd__a22o_1 \U$$3205  (.A1(net1094),
    .A2(net504),
    .B1(net1086),
    .B2(net777),
    .X(\t$6043 ));
 sky130_fd_sc_hd__xor2_1 \U$$3206  (.A(\t$6043 ),
    .B(net1350),
    .X(booth_b46_m24));
 sky130_fd_sc_hd__a22o_1 \U$$3207  (.A1(net1086),
    .A2(net502),
    .B1(net1076),
    .B2(net775),
    .X(\t$6044 ));
 sky130_fd_sc_hd__xor2_1 \U$$3208  (.A(\t$6044 ),
    .B(net1349),
    .X(booth_b46_m25));
 sky130_fd_sc_hd__a22o_1 \U$$3209  (.A1(net1073),
    .A2(net501),
    .B1(net1065),
    .B2(net774),
    .X(\t$6045 ));
 sky130_fd_sc_hd__xor2_1 \U$$321  (.A(\t$4569 ),
    .B(net1274),
    .X(booth_b4_m20));
 sky130_fd_sc_hd__xor2_1 \U$$3210  (.A(\t$6045 ),
    .B(net1348),
    .X(booth_b46_m26));
 sky130_fd_sc_hd__a22o_1 \U$$3211  (.A1(net1065),
    .A2(net501),
    .B1(net1059),
    .B2(net774),
    .X(\t$6046 ));
 sky130_fd_sc_hd__xor2_1 \U$$3212  (.A(\t$6046 ),
    .B(net1348),
    .X(booth_b46_m27));
 sky130_fd_sc_hd__a22o_1 \U$$3213  (.A1(net1059),
    .A2(net501),
    .B1(net1054),
    .B2(net774),
    .X(\t$6047 ));
 sky130_fd_sc_hd__xor2_1 \U$$3214  (.A(\t$6047 ),
    .B(net1348),
    .X(booth_b46_m28));
 sky130_fd_sc_hd__a22o_1 \U$$3215  (.A1(net1051),
    .A2(net503),
    .B1(net1043),
    .B2(net776),
    .X(\t$6048 ));
 sky130_fd_sc_hd__xor2_1 \U$$3216  (.A(\t$6048 ),
    .B(net1351),
    .X(booth_b46_m29));
 sky130_fd_sc_hd__a22o_1 \U$$3217  (.A1(net1043),
    .A2(net503),
    .B1(net1027),
    .B2(net776),
    .X(\t$6049 ));
 sky130_fd_sc_hd__xor2_1 \U$$3218  (.A(\t$6049 ),
    .B(net1351),
    .X(booth_b46_m30));
 sky130_fd_sc_hd__a22o_1 \U$$3219  (.A1(net1027),
    .A2(net502),
    .B1(net1019),
    .B2(net775),
    .X(\t$6050 ));
 sky130_fd_sc_hd__a22o_1 \U$$322  (.A1(net1114),
    .A2(net528),
    .B1(net1105),
    .B2(net801),
    .X(\t$4570 ));
 sky130_fd_sc_hd__xor2_1 \U$$3220  (.A(\t$6050 ),
    .B(net1349),
    .X(booth_b46_m31));
 sky130_fd_sc_hd__a22o_1 \U$$3221  (.A1(net1019),
    .A2(net503),
    .B1(net1002),
    .B2(net776),
    .X(\t$6051 ));
 sky130_fd_sc_hd__xor2_1 \U$$3222  (.A(\t$6051 ),
    .B(net1351),
    .X(booth_b46_m32));
 sky130_fd_sc_hd__a22o_1 \U$$3223  (.A1(net1002),
    .A2(net504),
    .B1(net994),
    .B2(net777),
    .X(\t$6052 ));
 sky130_fd_sc_hd__xor2_1 \U$$3224  (.A(\t$6052 ),
    .B(net1350),
    .X(booth_b46_m33));
 sky130_fd_sc_hd__a22o_1 \U$$3225  (.A1(net994),
    .A2(net504),
    .B1(net985),
    .B2(net777),
    .X(\t$6053 ));
 sky130_fd_sc_hd__xor2_1 \U$$3226  (.A(\t$6053 ),
    .B(net1350),
    .X(booth_b46_m34));
 sky130_fd_sc_hd__a22o_1 \U$$3227  (.A1(net985),
    .A2(net503),
    .B1(net976),
    .B2(net776),
    .X(\t$6054 ));
 sky130_fd_sc_hd__xor2_1 \U$$3228  (.A(\t$6054 ),
    .B(net1351),
    .X(booth_b46_m35));
 sky130_fd_sc_hd__a22o_1 \U$$3229  (.A1(net975),
    .A2(net503),
    .B1(net966),
    .B2(net776),
    .X(\t$6055 ));
 sky130_fd_sc_hd__xor2_1 \U$$323  (.A(\t$4570 ),
    .B(net1274),
    .X(booth_b4_m21));
 sky130_fd_sc_hd__xor2_1 \U$$3230  (.A(\t$6055 ),
    .B(net1351),
    .X(booth_b46_m36));
 sky130_fd_sc_hd__a22o_1 \U$$3231  (.A1(net966),
    .A2(net503),
    .B1(net959),
    .B2(net776),
    .X(\t$6056 ));
 sky130_fd_sc_hd__xor2_1 \U$$3232  (.A(\t$6056 ),
    .B(net1351),
    .X(booth_b46_m37));
 sky130_fd_sc_hd__a22o_1 \U$$3233  (.A1(net959),
    .A2(net503),
    .B1(net950),
    .B2(net776),
    .X(\t$6057 ));
 sky130_fd_sc_hd__xor2_1 \U$$3234  (.A(\t$6057 ),
    .B(net1351),
    .X(booth_b46_m38));
 sky130_fd_sc_hd__a22o_1 \U$$3235  (.A1(net950),
    .A2(net503),
    .B1(net942),
    .B2(net776),
    .X(\t$6058 ));
 sky130_fd_sc_hd__xor2_1 \U$$3236  (.A(\t$6058 ),
    .B(net1351),
    .X(booth_b46_m39));
 sky130_fd_sc_hd__a22o_1 \U$$3237  (.A1(net942),
    .A2(net503),
    .B1(net926),
    .B2(net776),
    .X(\t$6059 ));
 sky130_fd_sc_hd__xor2_1 \U$$3238  (.A(\t$6059 ),
    .B(net1351),
    .X(booth_b46_m40));
 sky130_fd_sc_hd__a22o_1 \U$$3239  (.A1(net927),
    .A2(net503),
    .B1(net1748),
    .B2(net776),
    .X(\t$6060 ));
 sky130_fd_sc_hd__a22o_1 \U$$324  (.A1(net1105),
    .A2(net527),
    .B1(net1097),
    .B2(net800),
    .X(\t$4571 ));
 sky130_fd_sc_hd__xor2_1 \U$$3240  (.A(\t$6060 ),
    .B(net1351),
    .X(booth_b46_m41));
 sky130_fd_sc_hd__a22o_1 \U$$3241  (.A1(net1748),
    .A2(net504),
    .B1(net1740),
    .B2(net777),
    .X(\t$6061 ));
 sky130_fd_sc_hd__xor2_1 \U$$3242  (.A(\t$6061 ),
    .B(net1350),
    .X(booth_b46_m42));
 sky130_fd_sc_hd__a22o_1 \U$$3243  (.A1(net1740),
    .A2(net504),
    .B1(net1732),
    .B2(net777),
    .X(\t$6062 ));
 sky130_fd_sc_hd__xor2_1 \U$$3244  (.A(\t$6062 ),
    .B(net1350),
    .X(booth_b46_m43));
 sky130_fd_sc_hd__a22o_1 \U$$3245  (.A1(net1735),
    .A2(net508),
    .B1(net1727),
    .B2(net781),
    .X(\t$6063 ));
 sky130_fd_sc_hd__xor2_1 \U$$3246  (.A(\t$6063 ),
    .B(net1356),
    .X(booth_b46_m44));
 sky130_fd_sc_hd__a22o_1 \U$$3247  (.A1(net1726),
    .A2(net507),
    .B1(net1717),
    .B2(net780),
    .X(\t$6064 ));
 sky130_fd_sc_hd__xor2_1 \U$$3248  (.A(\t$6064 ),
    .B(net1355),
    .X(booth_b46_m45));
 sky130_fd_sc_hd__a22o_1 \U$$3249  (.A1(net1717),
    .A2(net507),
    .B1(net1708),
    .B2(net780),
    .X(\t$6065 ));
 sky130_fd_sc_hd__xor2_1 \U$$325  (.A(\t$4571 ),
    .B(net1273),
    .X(booth_b4_m22));
 sky130_fd_sc_hd__xor2_1 \U$$3250  (.A(\t$6065 ),
    .B(net1355),
    .X(booth_b46_m46));
 sky130_fd_sc_hd__a22o_1 \U$$3251  (.A1(net1708),
    .A2(net507),
    .B1(net1700),
    .B2(net780),
    .X(\t$6066 ));
 sky130_fd_sc_hd__xor2_1 \U$$3252  (.A(\t$6066 ),
    .B(net1355),
    .X(booth_b46_m47));
 sky130_fd_sc_hd__a22o_1 \U$$3253  (.A1(net1700),
    .A2(net507),
    .B1(net1693),
    .B2(net780),
    .X(\t$6067 ));
 sky130_fd_sc_hd__xor2_1 \U$$3254  (.A(\t$6067 ),
    .B(net1355),
    .X(booth_b46_m48));
 sky130_fd_sc_hd__a22o_1 \U$$3255  (.A1(net1691),
    .A2(net505),
    .B1(net1683),
    .B2(net778),
    .X(\t$6068 ));
 sky130_fd_sc_hd__xor2_1 \U$$3256  (.A(\t$6068 ),
    .B(net1354),
    .X(booth_b46_m49));
 sky130_fd_sc_hd__a22o_1 \U$$3257  (.A1(net1684),
    .A2(net507),
    .B1(net1660),
    .B2(net780),
    .X(\t$6069 ));
 sky130_fd_sc_hd__xor2_1 \U$$3258  (.A(\t$6069 ),
    .B(net1355),
    .X(booth_b46_m50));
 sky130_fd_sc_hd__a22o_1 \U$$3259  (.A1(net1660),
    .A2(net507),
    .B1(net1652),
    .B2(net780),
    .X(\t$6070 ));
 sky130_fd_sc_hd__a22o_1 \U$$326  (.A1(net1097),
    .A2(net527),
    .B1(net1088),
    .B2(net800),
    .X(\t$4572 ));
 sky130_fd_sc_hd__xor2_1 \U$$3260  (.A(\t$6070 ),
    .B(net1355),
    .X(booth_b46_m51));
 sky130_fd_sc_hd__a22o_1 \U$$3261  (.A1(net1652),
    .A2(net507),
    .B1(net1644),
    .B2(net780),
    .X(\t$6071 ));
 sky130_fd_sc_hd__xor2_1 \U$$3262  (.A(\t$6071 ),
    .B(net1355),
    .X(booth_b46_m52));
 sky130_fd_sc_hd__a22o_1 \U$$3263  (.A1(net1644),
    .A2(net508),
    .B1(net1635),
    .B2(net781),
    .X(\t$6072 ));
 sky130_fd_sc_hd__xor2_1 \U$$3264  (.A(\t$6072 ),
    .B(net1355),
    .X(booth_b46_m53));
 sky130_fd_sc_hd__a22o_1 \U$$3265  (.A1(net1635),
    .A2(net508),
    .B1(net1626),
    .B2(net781),
    .X(\t$6073 ));
 sky130_fd_sc_hd__xor2_1 \U$$3266  (.A(\t$6073 ),
    .B(net1355),
    .X(booth_b46_m54));
 sky130_fd_sc_hd__a22o_1 \U$$3267  (.A1(net1626),
    .A2(net508),
    .B1(net1618),
    .B2(net781),
    .X(\t$6074 ));
 sky130_fd_sc_hd__xor2_1 \U$$3268  (.A(\t$6074 ),
    .B(net1355),
    .X(booth_b46_m55));
 sky130_fd_sc_hd__a22o_1 \U$$3269  (.A1(net1618),
    .A2(net507),
    .B1(net1609),
    .B2(net780),
    .X(\t$6075 ));
 sky130_fd_sc_hd__xor2_1 \U$$327  (.A(\t$4572 ),
    .B(net1273),
    .X(booth_b4_m23));
 sky130_fd_sc_hd__xor2_1 \U$$3270  (.A(\t$6075 ),
    .B(net1356),
    .X(booth_b46_m56));
 sky130_fd_sc_hd__a22o_1 \U$$3271  (.A1(net1608),
    .A2(net504),
    .B1(net1600),
    .B2(net777),
    .X(\t$6076 ));
 sky130_fd_sc_hd__xor2_1 \U$$3272  (.A(\t$6076 ),
    .B(net1350),
    .X(booth_b46_m57));
 sky130_fd_sc_hd__a22o_1 \U$$3273  (.A1(net1602),
    .A2(net507),
    .B1(net1593),
    .B2(net780),
    .X(\t$6077 ));
 sky130_fd_sc_hd__xor2_1 \U$$3274  (.A(\t$6077 ),
    .B(net1356),
    .X(booth_b46_m58));
 sky130_fd_sc_hd__a22o_1 \U$$3275  (.A1(net1593),
    .A2(net507),
    .B1(net1585),
    .B2(net780),
    .X(\t$6078 ));
 sky130_fd_sc_hd__xor2_1 \U$$3276  (.A(\t$6078 ),
    .B(net1356),
    .X(booth_b46_m59));
 sky130_fd_sc_hd__a22o_1 \U$$3277  (.A1(net1583),
    .A2(net508),
    .B1(net1556),
    .B2(net781),
    .X(\t$6079 ));
 sky130_fd_sc_hd__xor2_1 \U$$3278  (.A(\t$6079 ),
    .B(net1356),
    .X(booth_b46_m60));
 sky130_fd_sc_hd__a22o_1 \U$$3279  (.A1(net1555),
    .A2(net508),
    .B1(net1547),
    .B2(net781),
    .X(\t$6080 ));
 sky130_fd_sc_hd__a22o_1 \U$$328  (.A1(net1088),
    .A2(net527),
    .B1(net1080),
    .B2(net800),
    .X(\t$4573 ));
 sky130_fd_sc_hd__xor2_1 \U$$3280  (.A(\t$6080 ),
    .B(net1356),
    .X(booth_b46_m61));
 sky130_fd_sc_hd__a22o_1 \U$$3281  (.A1(net1548),
    .A2(net508),
    .B1(net1540),
    .B2(net781),
    .X(\t$6081 ));
 sky130_fd_sc_hd__xor2_1 \U$$3282  (.A(\t$6081 ),
    .B(net1356),
    .X(booth_b46_m62));
 sky130_fd_sc_hd__a22o_1 \U$$3283  (.A1(net1540),
    .A2(net508),
    .B1(net1532),
    .B2(net781),
    .X(\t$6082 ));
 sky130_fd_sc_hd__xor2_1 \U$$3284  (.A(\t$6082 ),
    .B(net1356),
    .X(booth_b46_m63));
 sky130_fd_sc_hd__a22o_1 \U$$3285  (.A1(net1532),
    .A2(net504),
    .B1(net1790),
    .B2(net777),
    .X(\t$6083 ));
 sky130_fd_sc_hd__xor2_1 \U$$3286  (.A(\t$6083 ),
    .B(net1350),
    .X(booth_b46_m64));
 sky130_fd_sc_hd__inv_1 \U$$3287  (.A(net1356),
    .Y(\notsign$6084 ));
 sky130_fd_sc_hd__inv_1 \U$$3288  (.A(net1350),
    .Y(\notblock$6085[0] ));
 sky130_fd_sc_hd__inv_1 \U$$3289  (.A(net43),
    .Y(\notblock$6085[1] ));
 sky130_fd_sc_hd__xor2_1 \U$$329  (.A(\t$4573 ),
    .B(net1273),
    .X(booth_b4_m24));
 sky130_fd_sc_hd__inv_1 \U$$3290  (.A(net1340),
    .Y(\notblock$6085[2] ));
 sky130_fd_sc_hd__and2_1 \U$$3291  (.A(net1340),
    .B(\notblock$6085[1] ),
    .X(\t$6086 ));
 sky130_fd_sc_hd__a32o_2 \U$$3292  (.A1(\notblock$6085[2] ),
    .A2(net43),
    .A3(net1352),
    .B1(\t$6086 ),
    .B2(\notblock$6085[0] ),
    .X(\sel_0$6087 ));
 sky130_fd_sc_hd__xor2_4 \U$$3293  (.A(net43),
    .B(net1352),
    .X(\sel_1$6088 ));
 sky130_fd_sc_hd__a22o_1 \U$$3294  (.A1(net1791),
    .A2(net493),
    .B1(net1229),
    .B2(net766),
    .X(\t$6089 ));
 sky130_fd_sc_hd__xor2_1 \U$$3295  (.A(\t$6089 ),
    .B(net1338),
    .X(booth_b48_m0));
 sky130_fd_sc_hd__a22o_1 \U$$3296  (.A1(net1229),
    .A2(net493),
    .B1(net1125),
    .B2(net766),
    .X(\t$6090 ));
 sky130_fd_sc_hd__xor2_1 \U$$3297  (.A(\t$6090 ),
    .B(net1338),
    .X(booth_b48_m1));
 sky130_fd_sc_hd__a22o_1 \U$$3298  (.A1(net1125),
    .A2(net493),
    .B1(net1034),
    .B2(net766),
    .X(\t$6091 ));
 sky130_fd_sc_hd__xor2_1 \U$$3299  (.A(\t$6091 ),
    .B(net1339),
    .X(booth_b48_m2));
 sky130_fd_sc_hd__xor2_1 \U$$33  (.A(\t$4423 ),
    .B(net1574),
    .X(booth_b0_m13));
 sky130_fd_sc_hd__a22o_1 \U$$330  (.A1(net1080),
    .A2(net527),
    .B1(net1071),
    .B2(net800),
    .X(\t$4574 ));
 sky130_fd_sc_hd__a22o_1 \U$$3300  (.A1(net1034),
    .A2(net496),
    .B1(net935),
    .B2(net769),
    .X(\t$6092 ));
 sky130_fd_sc_hd__xor2_1 \U$$3301  (.A(\t$6092 ),
    .B(net1339),
    .X(booth_b48_m3));
 sky130_fd_sc_hd__a22o_1 \U$$3302  (.A1(net938),
    .A2(net497),
    .B1(net1678),
    .B2(net770),
    .X(\t$6093 ));
 sky130_fd_sc_hd__xor2_1 \U$$3303  (.A(\t$6093 ),
    .B(net1343),
    .X(booth_b48_m4));
 sky130_fd_sc_hd__a22o_1 \U$$3304  (.A1(net1677),
    .A2(net497),
    .B1(net1566),
    .B2(net770),
    .X(\t$6094 ));
 sky130_fd_sc_hd__xor2_1 \U$$3305  (.A(\t$6094 ),
    .B(net1343),
    .X(booth_b48_m5));
 sky130_fd_sc_hd__a22o_1 \U$$3306  (.A1(net1566),
    .A2(net497),
    .B1(net1525),
    .B2(net770),
    .X(\t$6095 ));
 sky130_fd_sc_hd__xor2_1 \U$$3307  (.A(\t$6095 ),
    .B(net1343),
    .X(booth_b48_m6));
 sky130_fd_sc_hd__a22o_1 \U$$3308  (.A1(net1525),
    .A2(net497),
    .B1(net1517),
    .B2(net770),
    .X(\t$6096 ));
 sky130_fd_sc_hd__xor2_1 \U$$3309  (.A(\t$6096 ),
    .B(net1343),
    .X(booth_b48_m7));
 sky130_fd_sc_hd__xor2_1 \U$$331  (.A(\t$4574 ),
    .B(net1273),
    .X(booth_b4_m25));
 sky130_fd_sc_hd__a22o_1 \U$$3310  (.A1(net1517),
    .A2(net500),
    .B1(net1510),
    .B2(net773),
    .X(\t$6097 ));
 sky130_fd_sc_hd__xor2_1 \U$$3311  (.A(\t$6097 ),
    .B(net1346),
    .X(booth_b48_m8));
 sky130_fd_sc_hd__a22o_1 \U$$3312  (.A1(net1510),
    .A2(net500),
    .B1(net1501),
    .B2(net773),
    .X(\t$6098 ));
 sky130_fd_sc_hd__xor2_1 \U$$3313  (.A(\t$6098 ),
    .B(net1346),
    .X(booth_b48_m9));
 sky130_fd_sc_hd__a22o_1 \U$$3314  (.A1(net1497),
    .A2(net496),
    .B1(net1223),
    .B2(net769),
    .X(\t$6099 ));
 sky130_fd_sc_hd__xor2_1 \U$$3315  (.A(\t$6099 ),
    .B(net1339),
    .X(booth_b48_m10));
 sky130_fd_sc_hd__a22o_1 \U$$3316  (.A1(net1222),
    .A2(net493),
    .B1(net1214),
    .B2(net766),
    .X(\t$6100 ));
 sky130_fd_sc_hd__xor2_1 \U$$3317  (.A(\t$6100 ),
    .B(net1338),
    .X(booth_b48_m11));
 sky130_fd_sc_hd__a22o_1 \U$$3318  (.A1(net1214),
    .A2(net493),
    .B1(net1202),
    .B2(net766),
    .X(\t$6101 ));
 sky130_fd_sc_hd__xor2_1 \U$$3319  (.A(\t$6101 ),
    .B(net1338),
    .X(booth_b48_m12));
 sky130_fd_sc_hd__a22o_1 \U$$332  (.A1(net1071),
    .A2(net527),
    .B1(net1063),
    .B2(net800),
    .X(\t$4575 ));
 sky130_fd_sc_hd__a22o_1 \U$$3320  (.A1(net1205),
    .A2(net493),
    .B1(net1196),
    .B2(net766),
    .X(\t$6102 ));
 sky130_fd_sc_hd__xor2_1 \U$$3321  (.A(\t$6102 ),
    .B(net1338),
    .X(booth_b48_m13));
 sky130_fd_sc_hd__a22o_1 \U$$3322  (.A1(net1196),
    .A2(net496),
    .B1(net1178),
    .B2(net769),
    .X(\t$6103 ));
 sky130_fd_sc_hd__xor2_1 \U$$3323  (.A(\t$6103 ),
    .B(net1339),
    .X(booth_b48_m14));
 sky130_fd_sc_hd__a22o_1 \U$$3324  (.A1(net1177),
    .A2(net493),
    .B1(net1168),
    .B2(net766),
    .X(\t$6104 ));
 sky130_fd_sc_hd__xor2_1 \U$$3325  (.A(\t$6104 ),
    .B(net1338),
    .X(booth_b48_m15));
 sky130_fd_sc_hd__a22o_1 \U$$3326  (.A1(net1172),
    .A2(net497),
    .B1(net1163),
    .B2(net770),
    .X(\t$6105 ));
 sky130_fd_sc_hd__xor2_1 \U$$3327  (.A(\t$6105 ),
    .B(net1343),
    .X(booth_b48_m16));
 sky130_fd_sc_hd__a22o_1 \U$$3328  (.A1(net1163),
    .A2(net497),
    .B1(net1153),
    .B2(net770),
    .X(\t$6106 ));
 sky130_fd_sc_hd__xor2_1 \U$$3329  (.A(\t$6106 ),
    .B(net1343),
    .X(booth_b48_m17));
 sky130_fd_sc_hd__xor2_1 \U$$333  (.A(\t$4575 ),
    .B(net1273),
    .X(booth_b4_m26));
 sky130_fd_sc_hd__a22o_1 \U$$3330  (.A1(net1153),
    .A2(net497),
    .B1(net1145),
    .B2(net770),
    .X(\t$6107 ));
 sky130_fd_sc_hd__xor2_1 \U$$3331  (.A(\t$6107 ),
    .B(net1343),
    .X(booth_b48_m18));
 sky130_fd_sc_hd__a22o_1 \U$$3332  (.A1(net1145),
    .A2(net497),
    .B1(net1137),
    .B2(net770),
    .X(\t$6108 ));
 sky130_fd_sc_hd__xor2_1 \U$$3333  (.A(\t$6108 ),
    .B(net1343),
    .X(booth_b48_m19));
 sky130_fd_sc_hd__a22o_1 \U$$3334  (.A1(net1137),
    .A2(net497),
    .B1(net1121),
    .B2(net770),
    .X(\t$6109 ));
 sky130_fd_sc_hd__xor2_1 \U$$3335  (.A(\t$6109 ),
    .B(net1343),
    .X(booth_b48_m20));
 sky130_fd_sc_hd__a22o_1 \U$$3336  (.A1(net1121),
    .A2(net500),
    .B1(net1113),
    .B2(net773),
    .X(\t$6110 ));
 sky130_fd_sc_hd__xor2_1 \U$$3337  (.A(\t$6110 ),
    .B(net1343),
    .X(booth_b48_m21));
 sky130_fd_sc_hd__a22o_1 \U$$3338  (.A1(net1111),
    .A2(net495),
    .B1(net1102),
    .B2(net768),
    .X(\t$6111 ));
 sky130_fd_sc_hd__xor2_1 \U$$3339  (.A(\t$6111 ),
    .B(net1340),
    .X(booth_b48_m22));
 sky130_fd_sc_hd__a22o_1 \U$$334  (.A1(net1063),
    .A2(net527),
    .B1(net1055),
    .B2(net800),
    .X(\t$4576 ));
 sky130_fd_sc_hd__a22o_1 \U$$3340  (.A1(net1102),
    .A2(net496),
    .B1(net1094),
    .B2(net769),
    .X(\t$6112 ));
 sky130_fd_sc_hd__xor2_1 \U$$3341  (.A(\t$6112 ),
    .B(net1339),
    .X(booth_b48_m23));
 sky130_fd_sc_hd__a22o_1 \U$$3342  (.A1(net1090),
    .A2(net493),
    .B1(net1082),
    .B2(net766),
    .X(\t$6113 ));
 sky130_fd_sc_hd__xor2_1 \U$$3343  (.A(\t$6113 ),
    .B(net1338),
    .X(booth_b48_m24));
 sky130_fd_sc_hd__a22o_1 \U$$3344  (.A1(net1082),
    .A2(net493),
    .B1(net1073),
    .B2(net766),
    .X(\t$6114 ));
 sky130_fd_sc_hd__xor2_1 \U$$3345  (.A(\t$6114 ),
    .B(net1338),
    .X(booth_b48_m25));
 sky130_fd_sc_hd__a22o_1 \U$$3346  (.A1(net1073),
    .A2(net493),
    .B1(net1065),
    .B2(net766),
    .X(\t$6115 ));
 sky130_fd_sc_hd__xor2_1 \U$$3347  (.A(\t$6115 ),
    .B(net1338),
    .X(booth_b48_m26));
 sky130_fd_sc_hd__a22o_1 \U$$3348  (.A1(net1068),
    .A2(net494),
    .B1(net1060),
    .B2(net767),
    .X(\t$6116 ));
 sky130_fd_sc_hd__xor2_1 \U$$3349  (.A(\t$6116 ),
    .B(net1341),
    .X(booth_b48_m27));
 sky130_fd_sc_hd__xor2_1 \U$$335  (.A(\t$4576 ),
    .B(net1273),
    .X(booth_b4_m27));
 sky130_fd_sc_hd__a22o_1 \U$$3350  (.A1(net1060),
    .A2(net494),
    .B1(net1051),
    .B2(net767),
    .X(\t$6117 ));
 sky130_fd_sc_hd__xor2_1 \U$$3351  (.A(\t$6117 ),
    .B(net1341),
    .X(booth_b48_m28));
 sky130_fd_sc_hd__a22o_1 \U$$3352  (.A1(net1051),
    .A2(net495),
    .B1(net1043),
    .B2(net768),
    .X(\t$6118 ));
 sky130_fd_sc_hd__xor2_1 \U$$3353  (.A(\t$6118 ),
    .B(net1340),
    .X(booth_b48_m29));
 sky130_fd_sc_hd__a22o_1 \U$$3354  (.A1(net1043),
    .A2(net494),
    .B1(net1027),
    .B2(net767),
    .X(\t$6119 ));
 sky130_fd_sc_hd__xor2_1 \U$$3355  (.A(\t$6119 ),
    .B(net1341),
    .X(booth_b48_m30));
 sky130_fd_sc_hd__a22o_1 \U$$3356  (.A1(net1027),
    .A2(net494),
    .B1(net1019),
    .B2(net767),
    .X(\t$6120 ));
 sky130_fd_sc_hd__xor2_1 \U$$3357  (.A(\t$6120 ),
    .B(net1340),
    .X(booth_b48_m31));
 sky130_fd_sc_hd__a22o_1 \U$$3358  (.A1(net1019),
    .A2(net495),
    .B1(net1002),
    .B2(net768),
    .X(\t$6121 ));
 sky130_fd_sc_hd__xor2_1 \U$$3359  (.A(\t$6121 ),
    .B(net1340),
    .X(booth_b48_m32));
 sky130_fd_sc_hd__a22o_1 \U$$336  (.A1(net1056),
    .A2(net528),
    .B1(net1048),
    .B2(net801),
    .X(\t$4577 ));
 sky130_fd_sc_hd__a22o_1 \U$$3360  (.A1(net1002),
    .A2(net494),
    .B1(net995),
    .B2(net767),
    .X(\t$6122 ));
 sky130_fd_sc_hd__xor2_1 \U$$3361  (.A(\t$6122 ),
    .B(net1341),
    .X(booth_b48_m33));
 sky130_fd_sc_hd__a22o_1 \U$$3362  (.A1(net994),
    .A2(net494),
    .B1(net984),
    .B2(net767),
    .X(\t$6123 ));
 sky130_fd_sc_hd__xor2_1 \U$$3363  (.A(\t$6123 ),
    .B(net1341),
    .X(booth_b48_m34));
 sky130_fd_sc_hd__a22o_1 \U$$3364  (.A1(net984),
    .A2(net494),
    .B1(net975),
    .B2(net767),
    .X(\t$6124 ));
 sky130_fd_sc_hd__xor2_1 \U$$3365  (.A(\t$6124 ),
    .B(net1341),
    .X(booth_b48_m35));
 sky130_fd_sc_hd__a22o_1 \U$$3366  (.A1(net975),
    .A2(net494),
    .B1(net966),
    .B2(net767),
    .X(\t$6125 ));
 sky130_fd_sc_hd__xor2_1 \U$$3367  (.A(\t$6125 ),
    .B(net1341),
    .X(booth_b48_m36));
 sky130_fd_sc_hd__a22o_1 \U$$3368  (.A1(net966),
    .A2(net495),
    .B1(net959),
    .B2(net768),
    .X(\t$6126 ));
 sky130_fd_sc_hd__xor2_1 \U$$3369  (.A(\t$6126 ),
    .B(net1341),
    .X(booth_b48_m37));
 sky130_fd_sc_hd__xor2_1 \U$$337  (.A(\t$4577 ),
    .B(net1276),
    .X(booth_b4_m28));
 sky130_fd_sc_hd__a22o_1 \U$$3370  (.A1(net959),
    .A2(net494),
    .B1(net950),
    .B2(net767),
    .X(\t$6127 ));
 sky130_fd_sc_hd__xor2_1 \U$$3371  (.A(\t$6127 ),
    .B(net1341),
    .X(booth_b48_m38));
 sky130_fd_sc_hd__a22o_1 \U$$3372  (.A1(net951),
    .A2(net494),
    .B1(net943),
    .B2(net767),
    .X(\t$6128 ));
 sky130_fd_sc_hd__xor2_1 \U$$3373  (.A(\t$6128 ),
    .B(net1341),
    .X(booth_b48_m39));
 sky130_fd_sc_hd__a22o_1 \U$$3374  (.A1(net943),
    .A2(net495),
    .B1(net927),
    .B2(net768),
    .X(\t$6129 ));
 sky130_fd_sc_hd__xor2_1 \U$$3375  (.A(\t$6129 ),
    .B(net1342),
    .X(booth_b48_m40));
 sky130_fd_sc_hd__a22o_1 \U$$3376  (.A1(net927),
    .A2(net495),
    .B1(net1748),
    .B2(net768),
    .X(\t$6130 ));
 sky130_fd_sc_hd__xor2_1 \U$$3377  (.A(\t$6130 ),
    .B(net1340),
    .X(booth_b48_m41));
 sky130_fd_sc_hd__a22o_1 \U$$3378  (.A1(net1751),
    .A2(net499),
    .B1(net1743),
    .B2(net772),
    .X(\t$6131 ));
 sky130_fd_sc_hd__xor2_1 \U$$3379  (.A(\t$6131 ),
    .B(net1345),
    .X(booth_b48_m42));
 sky130_fd_sc_hd__a22o_1 \U$$338  (.A1(net1050),
    .A2(net531),
    .B1(net1042),
    .B2(net804),
    .X(\t$4578 ));
 sky130_fd_sc_hd__a22o_1 \U$$3380  (.A1(net1742),
    .A2(net498),
    .B1(net1734),
    .B2(net771),
    .X(\t$6132 ));
 sky130_fd_sc_hd__xor2_1 \U$$3381  (.A(\t$6132 ),
    .B(net1344),
    .X(booth_b48_m43));
 sky130_fd_sc_hd__a22o_1 \U$$3382  (.A1(net1734),
    .A2(net498),
    .B1(net1726),
    .B2(net771),
    .X(\t$6133 ));
 sky130_fd_sc_hd__xor2_1 \U$$3383  (.A(\t$6133 ),
    .B(net1344),
    .X(booth_b48_m44));
 sky130_fd_sc_hd__a22o_1 \U$$3384  (.A1(net1726),
    .A2(net498),
    .B1(net1717),
    .B2(net771),
    .X(\t$6134 ));
 sky130_fd_sc_hd__xor2_1 \U$$3385  (.A(\t$6134 ),
    .B(net1344),
    .X(booth_b48_m45));
 sky130_fd_sc_hd__a22o_1 \U$$3386  (.A1(net1717),
    .A2(net498),
    .B1(net1708),
    .B2(net771),
    .X(\t$6135 ));
 sky130_fd_sc_hd__xor2_1 \U$$3387  (.A(\t$6135 ),
    .B(net1344),
    .X(booth_b48_m46));
 sky130_fd_sc_hd__a22o_1 \U$$3388  (.A1(net1706),
    .A2(net497),
    .B1(net1698),
    .B2(net770),
    .X(\t$6136 ));
 sky130_fd_sc_hd__xor2_1 \U$$3389  (.A(\t$6136 ),
    .B(net1346),
    .X(booth_b48_m47));
 sky130_fd_sc_hd__xor2_1 \U$$339  (.A(\t$4578 ),
    .B(net1277),
    .X(booth_b4_m29));
 sky130_fd_sc_hd__a22o_1 \U$$3390  (.A1(net1700),
    .A2(net498),
    .B1(net1693),
    .B2(net771),
    .X(\t$6137 ));
 sky130_fd_sc_hd__xor2_1 \U$$3391  (.A(\t$6137 ),
    .B(net1344),
    .X(booth_b48_m48));
 sky130_fd_sc_hd__a22o_1 \U$$3392  (.A1(net1693),
    .A2(net498),
    .B1(net1684),
    .B2(net771),
    .X(\t$6138 ));
 sky130_fd_sc_hd__xor2_1 \U$$3393  (.A(\t$6138 ),
    .B(net1344),
    .X(booth_b48_m49));
 sky130_fd_sc_hd__a22o_1 \U$$3394  (.A1(net1684),
    .A2(net498),
    .B1(net1660),
    .B2(net771),
    .X(\t$6139 ));
 sky130_fd_sc_hd__xor2_1 \U$$3395  (.A(\t$6139 ),
    .B(net1344),
    .X(booth_b48_m50));
 sky130_fd_sc_hd__a22o_1 \U$$3396  (.A1(net1660),
    .A2(net498),
    .B1(net1652),
    .B2(net771),
    .X(\t$6140 ));
 sky130_fd_sc_hd__xor2_1 \U$$3397  (.A(\t$6140 ),
    .B(net1344),
    .X(booth_b48_m51));
 sky130_fd_sc_hd__a22o_1 \U$$3398  (.A1(net1652),
    .A2(net498),
    .B1(net1644),
    .B2(net771),
    .X(\t$6141 ));
 sky130_fd_sc_hd__xor2_1 \U$$3399  (.A(\t$6141 ),
    .B(net1344),
    .X(booth_b48_m52));
 sky130_fd_sc_hd__a22o_1 \U$$34  (.A1(net1194),
    .A2(net448),
    .B1(net1175),
    .B2(net690),
    .X(\t$4424 ));
 sky130_fd_sc_hd__a22o_1 \U$$340  (.A1(net1042),
    .A2(net534),
    .B1(net1026),
    .B2(net807),
    .X(\t$4579 ));
 sky130_fd_sc_hd__a22o_1 \U$$3400  (.A1(net1644),
    .A2(net499),
    .B1(net1636),
    .B2(net772),
    .X(\t$6142 ));
 sky130_fd_sc_hd__xor2_1 \U$$3401  (.A(\t$6142 ),
    .B(net1346),
    .X(booth_b48_m53));
 sky130_fd_sc_hd__a22o_1 \U$$3402  (.A1(net1636),
    .A2(net499),
    .B1(net1626),
    .B2(net772),
    .X(\t$6143 ));
 sky130_fd_sc_hd__xor2_1 \U$$3403  (.A(\t$6143 ),
    .B(net1345),
    .X(booth_b48_m54));
 sky130_fd_sc_hd__a22o_1 \U$$3404  (.A1(net1624),
    .A2(net495),
    .B1(net1616),
    .B2(net768),
    .X(\t$6144 ));
 sky130_fd_sc_hd__xor2_1 \U$$3405  (.A(\t$6144 ),
    .B(net1340),
    .X(booth_b48_m55));
 sky130_fd_sc_hd__a22o_1 \U$$3406  (.A1(net1618),
    .A2(net498),
    .B1(net1609),
    .B2(net771),
    .X(\t$6145 ));
 sky130_fd_sc_hd__xor2_1 \U$$3407  (.A(\t$6145 ),
    .B(net1344),
    .X(booth_b48_m56));
 sky130_fd_sc_hd__a22o_1 \U$$3408  (.A1(net1609),
    .A2(net499),
    .B1(net1603),
    .B2(net772),
    .X(\t$6146 ));
 sky130_fd_sc_hd__xor2_1 \U$$3409  (.A(\t$6146 ),
    .B(net1345),
    .X(booth_b48_m57));
 sky130_fd_sc_hd__xor2_1 \U$$341  (.A(\t$4579 ),
    .B(net1278),
    .X(booth_b4_m30));
 sky130_fd_sc_hd__a22o_1 \U$$3410  (.A1(net1600),
    .A2(net499),
    .B1(net1591),
    .B2(net772),
    .X(\t$6147 ));
 sky130_fd_sc_hd__xor2_1 \U$$3411  (.A(\t$6147 ),
    .B(net1345),
    .X(booth_b48_m58));
 sky130_fd_sc_hd__a22o_1 \U$$3412  (.A1(net1591),
    .A2(net495),
    .B1(net1583),
    .B2(net768),
    .X(\t$6148 ));
 sky130_fd_sc_hd__xor2_1 \U$$3413  (.A(\t$6148 ),
    .B(net1340),
    .X(booth_b48_m59));
 sky130_fd_sc_hd__a22o_1 \U$$3414  (.A1(net1583),
    .A2(net499),
    .B1(net1556),
    .B2(net772),
    .X(\t$6149 ));
 sky130_fd_sc_hd__xor2_1 \U$$3415  (.A(\t$6149 ),
    .B(net1345),
    .X(booth_b48_m60));
 sky130_fd_sc_hd__a22o_1 \U$$3416  (.A1(net1556),
    .A2(net499),
    .B1(net1548),
    .B2(net772),
    .X(\t$6150 ));
 sky130_fd_sc_hd__xor2_1 \U$$3417  (.A(\t$6150 ),
    .B(net1345),
    .X(booth_b48_m61));
 sky130_fd_sc_hd__a22o_1 \U$$3418  (.A1(net1548),
    .A2(net495),
    .B1(net1540),
    .B2(net768),
    .X(\t$6151 ));
 sky130_fd_sc_hd__xor2_1 \U$$3419  (.A(\t$6151 ),
    .B(net1340),
    .X(booth_b48_m62));
 sky130_fd_sc_hd__a22o_1 \U$$342  (.A1(net1026),
    .A2(net534),
    .B1(net1018),
    .B2(net807),
    .X(\t$4580 ));
 sky130_fd_sc_hd__a22o_1 \U$$3420  (.A1(net1541),
    .A2(net499),
    .B1(net1532),
    .B2(net772),
    .X(\t$6152 ));
 sky130_fd_sc_hd__xor2_1 \U$$3421  (.A(\t$6152 ),
    .B(net1345),
    .X(booth_b48_m63));
 sky130_fd_sc_hd__a22o_1 \U$$3422  (.A1(net1533),
    .A2(net499),
    .B1(net1792),
    .B2(net772),
    .X(\t$6153 ));
 sky130_fd_sc_hd__xor2_1 \U$$3423  (.A(\t$6153 ),
    .B(net1345),
    .X(booth_b48_m64));
 sky130_fd_sc_hd__inv_1 \U$$3424  (.A(net1345),
    .Y(\notsign$6154 ));
 sky130_fd_sc_hd__inv_1 \U$$3425  (.A(net1342),
    .Y(\notblock$6155[0] ));
 sky130_fd_sc_hd__inv_1 \U$$3426  (.A(net46),
    .Y(\notblock$6155[1] ));
 sky130_fd_sc_hd__inv_1 \U$$3427  (.A(net1330),
    .Y(\notblock$6155[2] ));
 sky130_fd_sc_hd__and2_1 \U$$3428  (.A(net1330),
    .B(\notblock$6155[1] ),
    .X(\t$6156 ));
 sky130_fd_sc_hd__a32o_2 \U$$3429  (.A1(\notblock$6155[2] ),
    .A2(net46),
    .A3(net1342),
    .B1(\t$6156 ),
    .B2(\notblock$6155[0] ),
    .X(\sel_0$6157 ));
 sky130_fd_sc_hd__xor2_1 \U$$343  (.A(\t$4580 ),
    .B(net1278),
    .X(booth_b4_m31));
 sky130_fd_sc_hd__xor2_4 \U$$3430  (.A(net46),
    .B(net1342),
    .X(\sel_1$6158 ));
 sky130_fd_sc_hd__a22o_1 \U$$3431  (.A1(net1793),
    .A2(net484),
    .B1(net1228),
    .B2(net757),
    .X(\t$6159 ));
 sky130_fd_sc_hd__xor2_1 \U$$3432  (.A(\t$6159 ),
    .B(net1329),
    .X(booth_b50_m0));
 sky130_fd_sc_hd__a22o_1 \U$$3433  (.A1(net1229),
    .A2(net484),
    .B1(net1124),
    .B2(net757),
    .X(\t$6160 ));
 sky130_fd_sc_hd__xor2_1 \U$$3434  (.A(\t$6160 ),
    .B(net1329),
    .X(booth_b50_m1));
 sky130_fd_sc_hd__a22o_1 \U$$3435  (.A1(net1129),
    .A2(net488),
    .B1(net1037),
    .B2(net761),
    .X(\t$6161 ));
 sky130_fd_sc_hd__xor2_1 \U$$3436  (.A(\t$6161 ),
    .B(net1333),
    .X(booth_b50_m2));
 sky130_fd_sc_hd__a22o_1 \U$$3437  (.A1(net1037),
    .A2(net488),
    .B1(net938),
    .B2(net761),
    .X(\t$6162 ));
 sky130_fd_sc_hd__xor2_1 \U$$3438  (.A(\t$6162 ),
    .B(net1333),
    .X(booth_b50_m3));
 sky130_fd_sc_hd__a22o_1 \U$$3439  (.A1(net938),
    .A2(net488),
    .B1(net1677),
    .B2(net761),
    .X(\t$6163 ));
 sky130_fd_sc_hd__a22o_1 \U$$344  (.A1(net1017),
    .A2(net532),
    .B1(net1000),
    .B2(net805),
    .X(\t$4581 ));
 sky130_fd_sc_hd__xor2_1 \U$$3440  (.A(\t$6163 ),
    .B(net1333),
    .X(booth_b50_m4));
 sky130_fd_sc_hd__a22o_1 \U$$3441  (.A1(net1677),
    .A2(net488),
    .B1(net1566),
    .B2(net761),
    .X(\t$6164 ));
 sky130_fd_sc_hd__xor2_1 \U$$3442  (.A(\t$6164 ),
    .B(net1333),
    .X(booth_b50_m5));
 sky130_fd_sc_hd__a22o_1 \U$$3443  (.A1(net1566),
    .A2(net492),
    .B1(net1525),
    .B2(net765),
    .X(\t$6165 ));
 sky130_fd_sc_hd__xor2_1 \U$$3444  (.A(\t$6165 ),
    .B(net1337),
    .X(booth_b50_m6));
 sky130_fd_sc_hd__a22o_1 \U$$3445  (.A1(net1525),
    .A2(net492),
    .B1(net1517),
    .B2(net765),
    .X(\t$6166 ));
 sky130_fd_sc_hd__xor2_1 \U$$3446  (.A(\t$6166 ),
    .B(net1337),
    .X(booth_b50_m7));
 sky130_fd_sc_hd__a22o_1 \U$$3447  (.A1(net1514),
    .A2(net487),
    .B1(net1506),
    .B2(net760),
    .X(\t$6167 ));
 sky130_fd_sc_hd__xor2_1 \U$$3448  (.A(\t$6167 ),
    .B(net1332),
    .X(booth_b50_m8));
 sky130_fd_sc_hd__a22o_1 \U$$3449  (.A1(net1507),
    .A2(net484),
    .B1(net1498),
    .B2(net757),
    .X(\t$6168 ));
 sky130_fd_sc_hd__xor2_1 \U$$345  (.A(\t$4581 ),
    .B(net1279),
    .X(booth_b4_m32));
 sky130_fd_sc_hd__xor2_1 \U$$3450  (.A(\t$6168 ),
    .B(net1329),
    .X(booth_b50_m9));
 sky130_fd_sc_hd__a22o_1 \U$$3451  (.A1(net1498),
    .A2(net484),
    .B1(net1222),
    .B2(net757),
    .X(\t$6169 ));
 sky130_fd_sc_hd__xor2_1 \U$$3452  (.A(\t$6169 ),
    .B(net1329),
    .X(booth_b50_m10));
 sky130_fd_sc_hd__a22o_1 \U$$3453  (.A1(net1222),
    .A2(net484),
    .B1(net1214),
    .B2(net757),
    .X(\t$6170 ));
 sky130_fd_sc_hd__xor2_1 \U$$3454  (.A(\t$6170 ),
    .B(net1329),
    .X(booth_b50_m11));
 sky130_fd_sc_hd__a22o_1 \U$$3455  (.A1(net1214),
    .A2(net487),
    .B1(net1205),
    .B2(net760),
    .X(\t$6171 ));
 sky130_fd_sc_hd__xor2_1 \U$$3456  (.A(\t$6171 ),
    .B(net1332),
    .X(booth_b50_m12));
 sky130_fd_sc_hd__a22o_1 \U$$3457  (.A1(net1205),
    .A2(net484),
    .B1(net1196),
    .B2(net757),
    .X(\t$6172 ));
 sky130_fd_sc_hd__xor2_1 \U$$3458  (.A(\t$6172 ),
    .B(net1329),
    .X(booth_b50_m13));
 sky130_fd_sc_hd__a22o_1 \U$$3459  (.A1(net1200),
    .A2(net488),
    .B1(net1181),
    .B2(net761),
    .X(\t$6173 ));
 sky130_fd_sc_hd__a22o_1 \U$$346  (.A1(net998),
    .A2(net527),
    .B1(net990),
    .B2(net800),
    .X(\t$4582 ));
 sky130_fd_sc_hd__xor2_1 \U$$3460  (.A(\t$6173 ),
    .B(net1333),
    .X(booth_b50_m14));
 sky130_fd_sc_hd__a22o_1 \U$$3461  (.A1(net1181),
    .A2(net488),
    .B1(net1172),
    .B2(net761),
    .X(\t$6174 ));
 sky130_fd_sc_hd__xor2_1 \U$$3462  (.A(\t$6174 ),
    .B(net1333),
    .X(booth_b50_m15));
 sky130_fd_sc_hd__a22o_1 \U$$3463  (.A1(net1172),
    .A2(net488),
    .B1(net1163),
    .B2(net761),
    .X(\t$6175 ));
 sky130_fd_sc_hd__xor2_1 \U$$3464  (.A(\t$6175 ),
    .B(net1333),
    .X(booth_b50_m16));
 sky130_fd_sc_hd__a22o_1 \U$$3465  (.A1(net1163),
    .A2(net488),
    .B1(net1153),
    .B2(net761),
    .X(\t$6176 ));
 sky130_fd_sc_hd__xor2_1 \U$$3466  (.A(\t$6176 ),
    .B(net1333),
    .X(booth_b50_m17));
 sky130_fd_sc_hd__a22o_1 \U$$3467  (.A1(net1153),
    .A2(net488),
    .B1(net1145),
    .B2(net761),
    .X(\t$6177 ));
 sky130_fd_sc_hd__xor2_1 \U$$3468  (.A(\t$6177 ),
    .B(net1333),
    .X(booth_b50_m18));
 sky130_fd_sc_hd__a22o_1 \U$$3469  (.A1(net1145),
    .A2(net488),
    .B1(net1137),
    .B2(net761),
    .X(\t$6178 ));
 sky130_fd_sc_hd__xor2_1 \U$$347  (.A(\t$4582 ),
    .B(net1273),
    .X(booth_b4_m33));
 sky130_fd_sc_hd__xor2_1 \U$$3470  (.A(\t$6178 ),
    .B(net1333),
    .X(booth_b50_m19));
 sky130_fd_sc_hd__a22o_1 \U$$3471  (.A1(net1135),
    .A2(net486),
    .B1(net1119),
    .B2(net759),
    .X(\t$6179 ));
 sky130_fd_sc_hd__xor2_1 \U$$3472  (.A(\t$6179 ),
    .B(net1330),
    .X(booth_b50_m20));
 sky130_fd_sc_hd__a22o_1 \U$$3473  (.A1(net1120),
    .A2(net487),
    .B1(net1111),
    .B2(net760),
    .X(\t$6180 ));
 sky130_fd_sc_hd__xor2_1 \U$$3474  (.A(\t$6180 ),
    .B(net1332),
    .X(booth_b50_m21));
 sky130_fd_sc_hd__a22o_1 \U$$3475  (.A1(net1107),
    .A2(net484),
    .B1(net1098),
    .B2(net757),
    .X(\t$6181 ));
 sky130_fd_sc_hd__xor2_1 \U$$3476  (.A(\t$6181 ),
    .B(net1329),
    .X(booth_b50_m22));
 sky130_fd_sc_hd__a22o_1 \U$$3477  (.A1(net1102),
    .A2(net484),
    .B1(net1090),
    .B2(net757),
    .X(\t$6182 ));
 sky130_fd_sc_hd__xor2_1 \U$$3478  (.A(\t$6182 ),
    .B(net1329),
    .X(booth_b50_m23));
 sky130_fd_sc_hd__a22o_1 \U$$3479  (.A1(net1090),
    .A2(net484),
    .B1(net1082),
    .B2(net757),
    .X(\t$6183 ));
 sky130_fd_sc_hd__a22o_1 \U$$348  (.A1(net991),
    .A2(net528),
    .B1(net983),
    .B2(net801),
    .X(\t$4583 ));
 sky130_fd_sc_hd__xor2_1 \U$$3480  (.A(\t$6183 ),
    .B(net1329),
    .X(booth_b50_m24));
 sky130_fd_sc_hd__a22o_1 \U$$3481  (.A1(net1086),
    .A2(net485),
    .B1(net1076),
    .B2(net758),
    .X(\t$6184 ));
 sky130_fd_sc_hd__xor2_1 \U$$3482  (.A(\t$6184 ),
    .B(net1331),
    .X(booth_b50_m25));
 sky130_fd_sc_hd__a22o_1 \U$$3483  (.A1(net1076),
    .A2(net484),
    .B1(net1068),
    .B2(net757),
    .X(\t$6185 ));
 sky130_fd_sc_hd__xor2_1 \U$$3484  (.A(\t$6185 ),
    .B(net1329),
    .X(booth_b50_m26));
 sky130_fd_sc_hd__a22o_1 \U$$3485  (.A1(net1068),
    .A2(net486),
    .B1(net1060),
    .B2(net759),
    .X(\t$6186 ));
 sky130_fd_sc_hd__xor2_1 \U$$3486  (.A(\t$6186 ),
    .B(net1330),
    .X(booth_b50_m27));
 sky130_fd_sc_hd__a22o_1 \U$$3487  (.A1(net1060),
    .A2(net485),
    .B1(net1051),
    .B2(net758),
    .X(\t$6187 ));
 sky130_fd_sc_hd__xor2_1 \U$$3488  (.A(\t$6187 ),
    .B(net1331),
    .X(booth_b50_m28));
 sky130_fd_sc_hd__a22o_1 \U$$3489  (.A1(net1051),
    .A2(net485),
    .B1(net1043),
    .B2(net758),
    .X(\t$6188 ));
 sky130_fd_sc_hd__xor2_1 \U$$349  (.A(\t$4583 ),
    .B(net1276),
    .X(booth_b4_m34));
 sky130_fd_sc_hd__xor2_1 \U$$3490  (.A(\t$6188 ),
    .B(net1331),
    .X(booth_b50_m29));
 sky130_fd_sc_hd__a22o_1 \U$$3491  (.A1(net1043),
    .A2(net486),
    .B1(net1027),
    .B2(net759),
    .X(\t$6189 ));
 sky130_fd_sc_hd__xor2_1 \U$$3492  (.A(\t$6189 ),
    .B(net1330),
    .X(booth_b50_m30));
 sky130_fd_sc_hd__a22o_1 \U$$3493  (.A1(net1027),
    .A2(net485),
    .B1(net1019),
    .B2(net758),
    .X(\t$6190 ));
 sky130_fd_sc_hd__xor2_1 \U$$3494  (.A(\t$6190 ),
    .B(net1331),
    .X(booth_b50_m31));
 sky130_fd_sc_hd__a22o_1 \U$$3495  (.A1(net1019),
    .A2(net485),
    .B1(net1002),
    .B2(net758),
    .X(\t$6191 ));
 sky130_fd_sc_hd__xor2_1 \U$$3496  (.A(\t$6191 ),
    .B(net1331),
    .X(booth_b50_m32));
 sky130_fd_sc_hd__a22o_1 \U$$3497  (.A1(net1003),
    .A2(net485),
    .B1(net995),
    .B2(net758),
    .X(\t$6192 ));
 sky130_fd_sc_hd__xor2_1 \U$$3498  (.A(\t$6192 ),
    .B(net1331),
    .X(booth_b50_m33));
 sky130_fd_sc_hd__a22o_1 \U$$3499  (.A1(net995),
    .A2(net485),
    .B1(net984),
    .B2(net758),
    .X(\t$6193 ));
 sky130_fd_sc_hd__xor2_1 \U$$35  (.A(\t$4424 ),
    .B(net1575),
    .X(booth_b0_m14));
 sky130_fd_sc_hd__a22o_1 \U$$350  (.A1(net986),
    .A2(net532),
    .B1(net974),
    .B2(net805),
    .X(\t$4584 ));
 sky130_fd_sc_hd__xor2_1 \U$$3500  (.A(\t$6193 ),
    .B(net1331),
    .X(booth_b50_m34));
 sky130_fd_sc_hd__a22o_1 \U$$3501  (.A1(net984),
    .A2(net485),
    .B1(net975),
    .B2(net758),
    .X(\t$6194 ));
 sky130_fd_sc_hd__xor2_1 \U$$3502  (.A(\t$6194 ),
    .B(net1331),
    .X(booth_b50_m35));
 sky130_fd_sc_hd__a22o_1 \U$$3503  (.A1(net975),
    .A2(net485),
    .B1(net966),
    .B2(net758),
    .X(\t$6195 ));
 sky130_fd_sc_hd__xor2_1 \U$$3504  (.A(\t$6195 ),
    .B(net1331),
    .X(booth_b50_m36));
 sky130_fd_sc_hd__a22o_1 \U$$3505  (.A1(net967),
    .A2(net485),
    .B1(net958),
    .B2(net758),
    .X(\t$6196 ));
 sky130_fd_sc_hd__xor2_1 \U$$3506  (.A(\t$6196 ),
    .B(net1331),
    .X(booth_b50_m37));
 sky130_fd_sc_hd__a22o_1 \U$$3507  (.A1(net959),
    .A2(net486),
    .B1(net951),
    .B2(net759),
    .X(\t$6197 ));
 sky130_fd_sc_hd__xor2_1 \U$$3508  (.A(\t$6197 ),
    .B(net1330),
    .X(booth_b50_m38));
 sky130_fd_sc_hd__a22o_1 \U$$3509  (.A1(net951),
    .A2(net486),
    .B1(net943),
    .B2(net759),
    .X(\t$6198 ));
 sky130_fd_sc_hd__xor2_1 \U$$351  (.A(\t$4584 ),
    .B(net1279),
    .X(booth_b4_m35));
 sky130_fd_sc_hd__xor2_1 \U$$3510  (.A(\t$6198 ),
    .B(net1330),
    .X(booth_b50_m39));
 sky130_fd_sc_hd__a22o_1 \U$$3511  (.A1(net946),
    .A2(net489),
    .B1(net930),
    .B2(net762),
    .X(\t$6199 ));
 sky130_fd_sc_hd__xor2_1 \U$$3512  (.A(\t$6199 ),
    .B(net1334),
    .X(booth_b50_m40));
 sky130_fd_sc_hd__a22o_1 \U$$3513  (.A1(net929),
    .A2(net490),
    .B1(net1750),
    .B2(net763),
    .X(\t$6200 ));
 sky130_fd_sc_hd__xor2_1 \U$$3514  (.A(\t$6200 ),
    .B(net1335),
    .X(booth_b50_m41));
 sky130_fd_sc_hd__a22o_1 \U$$3515  (.A1(net1750),
    .A2(net489),
    .B1(net1742),
    .B2(net762),
    .X(\t$6201 ));
 sky130_fd_sc_hd__xor2_1 \U$$3516  (.A(\t$6201 ),
    .B(net1334),
    .X(booth_b50_m42));
 sky130_fd_sc_hd__a22o_1 \U$$3517  (.A1(net1742),
    .A2(net490),
    .B1(net1734),
    .B2(net763),
    .X(\t$6202 ));
 sky130_fd_sc_hd__xor2_1 \U$$3518  (.A(\t$6202 ),
    .B(net1335),
    .X(booth_b50_m43));
 sky130_fd_sc_hd__a22o_1 \U$$3519  (.A1(net1735),
    .A2(net489),
    .B1(net1727),
    .B2(net762),
    .X(\t$6203 ));
 sky130_fd_sc_hd__a22o_1 \U$$352  (.A1(net973),
    .A2(net527),
    .B1(net964),
    .B2(net800),
    .X(\t$4585 ));
 sky130_fd_sc_hd__xor2_1 \U$$3520  (.A(\t$6203 ),
    .B(net1334),
    .X(booth_b50_m44));
 sky130_fd_sc_hd__a22o_1 \U$$3521  (.A1(net1725),
    .A2(net492),
    .B1(net1715),
    .B2(net765),
    .X(\t$6204 ));
 sky130_fd_sc_hd__xor2_1 \U$$3522  (.A(\t$6204 ),
    .B(net1337),
    .X(booth_b50_m45));
 sky130_fd_sc_hd__a22o_1 \U$$3523  (.A1(net1717),
    .A2(net490),
    .B1(net1708),
    .B2(net763),
    .X(\t$6205 ));
 sky130_fd_sc_hd__xor2_1 \U$$3524  (.A(\t$6205 ),
    .B(net1335),
    .X(booth_b50_m46));
 sky130_fd_sc_hd__a22o_1 \U$$3525  (.A1(net1708),
    .A2(net490),
    .B1(net1700),
    .B2(net763),
    .X(\t$6206 ));
 sky130_fd_sc_hd__xor2_1 \U$$3526  (.A(\t$6206 ),
    .B(net1335),
    .X(booth_b50_m47));
 sky130_fd_sc_hd__a22o_1 \U$$3527  (.A1(net1700),
    .A2(net490),
    .B1(net1693),
    .B2(net763),
    .X(\t$6207 ));
 sky130_fd_sc_hd__xor2_1 \U$$3528  (.A(\t$6207 ),
    .B(net1335),
    .X(booth_b50_m48));
 sky130_fd_sc_hd__a22o_1 \U$$3529  (.A1(net1693),
    .A2(net490),
    .B1(net1684),
    .B2(net763),
    .X(\t$6208 ));
 sky130_fd_sc_hd__xor2_1 \U$$353  (.A(\t$4585 ),
    .B(net1273),
    .X(booth_b4_m36));
 sky130_fd_sc_hd__xor2_1 \U$$3530  (.A(\t$6208 ),
    .B(net1335),
    .X(booth_b50_m49));
 sky130_fd_sc_hd__a22o_1 \U$$3531  (.A1(net1686),
    .A2(net490),
    .B1(net1661),
    .B2(net763),
    .X(\t$6209 ));
 sky130_fd_sc_hd__xor2_1 \U$$3532  (.A(\t$6209 ),
    .B(net1335),
    .X(booth_b50_m50));
 sky130_fd_sc_hd__a22o_1 \U$$3533  (.A1(net1661),
    .A2(net491),
    .B1(net1653),
    .B2(net764),
    .X(\t$6210 ));
 sky130_fd_sc_hd__xor2_1 \U$$3534  (.A(\t$6210 ),
    .B(net1335),
    .X(booth_b50_m51));
 sky130_fd_sc_hd__a22o_1 \U$$3535  (.A1(net1653),
    .A2(net491),
    .B1(net1645),
    .B2(net764),
    .X(\t$6211 ));
 sky130_fd_sc_hd__xor2_1 \U$$3536  (.A(\t$6211 ),
    .B(net1336),
    .X(booth_b50_m52));
 sky130_fd_sc_hd__a22o_1 \U$$3537  (.A1(net1644),
    .A2(net490),
    .B1(net1635),
    .B2(net763),
    .X(\t$6212 ));
 sky130_fd_sc_hd__xor2_1 \U$$3538  (.A(\t$6212 ),
    .B(net1335),
    .X(booth_b50_m53));
 sky130_fd_sc_hd__a22o_1 \U$$3539  (.A1(net1635),
    .A2(net490),
    .B1(net1626),
    .B2(net763),
    .X(\t$6213 ));
 sky130_fd_sc_hd__a22o_1 \U$$354  (.A1(net964),
    .A2(net527),
    .B1(net956),
    .B2(net800),
    .X(\t$4586 ));
 sky130_fd_sc_hd__xor2_1 \U$$3540  (.A(\t$6213 ),
    .B(net1335),
    .X(booth_b50_m54));
 sky130_fd_sc_hd__a22o_1 \U$$3541  (.A1(net1627),
    .A2(net490),
    .B1(net1618),
    .B2(net763),
    .X(\t$6214 ));
 sky130_fd_sc_hd__xor2_1 \U$$3542  (.A(\t$6214 ),
    .B(net1336),
    .X(booth_b50_m55));
 sky130_fd_sc_hd__a22o_1 \U$$3543  (.A1(net1616),
    .A2(net489),
    .B1(net1608),
    .B2(net762),
    .X(\t$6215 ));
 sky130_fd_sc_hd__xor2_1 \U$$3544  (.A(\t$6215 ),
    .B(net1334),
    .X(booth_b50_m56));
 sky130_fd_sc_hd__a22o_1 \U$$3545  (.A1(net1608),
    .A2(net486),
    .B1(net1600),
    .B2(net759),
    .X(\t$6216 ));
 sky130_fd_sc_hd__xor2_1 \U$$3546  (.A(\t$6216 ),
    .B(net1330),
    .X(booth_b50_m57));
 sky130_fd_sc_hd__a22o_1 \U$$3547  (.A1(net1600),
    .A2(net489),
    .B1(net1591),
    .B2(net762),
    .X(\t$6217 ));
 sky130_fd_sc_hd__xor2_1 \U$$3548  (.A(\t$6217 ),
    .B(net1334),
    .X(booth_b50_m58));
 sky130_fd_sc_hd__a22o_1 \U$$3549  (.A1(net1591),
    .A2(net489),
    .B1(net1583),
    .B2(net762),
    .X(\t$6218 ));
 sky130_fd_sc_hd__xor2_1 \U$$355  (.A(\t$4586 ),
    .B(net1273),
    .X(booth_b4_m37));
 sky130_fd_sc_hd__xor2_1 \U$$3550  (.A(\t$6218 ),
    .B(net1334),
    .X(booth_b50_m59));
 sky130_fd_sc_hd__a22o_1 \U$$3551  (.A1(net1583),
    .A2(net489),
    .B1(net1556),
    .B2(net762),
    .X(\t$6219 ));
 sky130_fd_sc_hd__xor2_1 \U$$3552  (.A(\t$6219 ),
    .B(net1334),
    .X(booth_b50_m60));
 sky130_fd_sc_hd__a22o_1 \U$$3553  (.A1(net1556),
    .A2(net491),
    .B1(net1549),
    .B2(net764),
    .X(\t$6220 ));
 sky130_fd_sc_hd__xor2_1 \U$$3554  (.A(\t$6220 ),
    .B(net1334),
    .X(booth_b50_m61));
 sky130_fd_sc_hd__a22o_1 \U$$3555  (.A1(net1549),
    .A2(net489),
    .B1(net1541),
    .B2(net762),
    .X(\t$6221 ));
 sky130_fd_sc_hd__xor2_1 \U$$3556  (.A(\t$6221 ),
    .B(net1334),
    .X(booth_b50_m62));
 sky130_fd_sc_hd__a22o_1 \U$$3557  (.A1(net1541),
    .A2(net489),
    .B1(net1533),
    .B2(net762),
    .X(\t$6222 ));
 sky130_fd_sc_hd__xor2_1 \U$$3558  (.A(\t$6222 ),
    .B(net1334),
    .X(booth_b50_m63));
 sky130_fd_sc_hd__a22o_1 \U$$3559  (.A1(net1533),
    .A2(net489),
    .B1(net1794),
    .B2(net762),
    .X(\t$6223 ));
 sky130_fd_sc_hd__a22o_1 \U$$356  (.A1(net956),
    .A2(net527),
    .B1(net948),
    .B2(net800),
    .X(\t$4587 ));
 sky130_fd_sc_hd__xor2_1 \U$$3560  (.A(\t$6223 ),
    .B(net1336),
    .X(booth_b50_m64));
 sky130_fd_sc_hd__inv_1 \U$$3561  (.A(net1330),
    .Y(\notsign$6224 ));
 sky130_fd_sc_hd__inv_1 \U$$3562  (.A(net1330),
    .Y(\notblock$6225[0] ));
 sky130_fd_sc_hd__inv_1 \U$$3563  (.A(net48),
    .Y(\notblock$6225[1] ));
 sky130_fd_sc_hd__inv_1 \U$$3564  (.A(net1321),
    .Y(\notblock$6225[2] ));
 sky130_fd_sc_hd__and2_1 \U$$3565  (.A(net1321),
    .B(\notblock$6225[1] ),
    .X(\t$6226 ));
 sky130_fd_sc_hd__a32o_4 \U$$3566  (.A1(\notblock$6225[2] ),
    .A2(net48),
    .A3(net1332),
    .B1(\t$6226 ),
    .B2(\notblock$6225[0] ),
    .X(\sel_0$6227 ));
 sky130_fd_sc_hd__xor2_4 \U$$3567  (.A(net48),
    .B(net1332),
    .X(\sel_1$6228 ));
 sky130_fd_sc_hd__a22o_1 \U$$3568  (.A1(net1795),
    .A2(net479),
    .B1(net1233),
    .B2(net752),
    .X(\t$6229 ));
 sky130_fd_sc_hd__xor2_1 \U$$3569  (.A(\t$6229 ),
    .B(net1319),
    .X(booth_b52_m0));
 sky130_fd_sc_hd__xor2_1 \U$$357  (.A(\t$4587 ),
    .B(net1273),
    .X(booth_b4_m38));
 sky130_fd_sc_hd__a22o_1 \U$$3570  (.A1(net1233),
    .A2(net480),
    .B1(net1129),
    .B2(net753),
    .X(\t$6230 ));
 sky130_fd_sc_hd__xor2_1 \U$$3571  (.A(\t$6230 ),
    .B(net1324),
    .X(booth_b52_m1));
 sky130_fd_sc_hd__a22o_1 \U$$3572  (.A1(net1129),
    .A2(net480),
    .B1(net1037),
    .B2(net753),
    .X(\t$6231 ));
 sky130_fd_sc_hd__xor2_1 \U$$3573  (.A(\t$6231 ),
    .B(net1324),
    .X(booth_b52_m2));
 sky130_fd_sc_hd__a22o_1 \U$$3574  (.A1(net1037),
    .A2(net480),
    .B1(net938),
    .B2(net753),
    .X(\t$6232 ));
 sky130_fd_sc_hd__xor2_1 \U$$3575  (.A(\t$6232 ),
    .B(net1324),
    .X(booth_b52_m3));
 sky130_fd_sc_hd__a22o_1 \U$$3576  (.A1(net938),
    .A2(net481),
    .B1(net1677),
    .B2(net754),
    .X(\t$6233 ));
 sky130_fd_sc_hd__xor2_1 \U$$3577  (.A(\t$6233 ),
    .B(net1325),
    .X(booth_b52_m4));
 sky130_fd_sc_hd__a22o_1 \U$$3578  (.A1(net1677),
    .A2(net481),
    .B1(net1566),
    .B2(net754),
    .X(\t$6234 ));
 sky130_fd_sc_hd__xor2_1 \U$$3579  (.A(\t$6234 ),
    .B(net1325),
    .X(booth_b52_m5));
 sky130_fd_sc_hd__a22o_1 \U$$358  (.A1(net948),
    .A2(net529),
    .B1(net940),
    .B2(net802),
    .X(\t$4588 ));
 sky130_fd_sc_hd__a22o_1 \U$$3580  (.A1(net1566),
    .A2(net481),
    .B1(net1525),
    .B2(net754),
    .X(\t$6235 ));
 sky130_fd_sc_hd__xor2_1 \U$$3581  (.A(\t$6235 ),
    .B(net1325),
    .X(booth_b52_m6));
 sky130_fd_sc_hd__a22o_1 \U$$3582  (.A1(net1522),
    .A2(net476),
    .B1(net1514),
    .B2(net749),
    .X(\t$6236 ));
 sky130_fd_sc_hd__xor2_1 \U$$3583  (.A(\t$6236 ),
    .B(net1319),
    .X(booth_b52_m7));
 sky130_fd_sc_hd__a22o_1 \U$$3584  (.A1(net1514),
    .A2(net476),
    .B1(net1507),
    .B2(net749),
    .X(\t$6237 ));
 sky130_fd_sc_hd__xor2_1 \U$$3585  (.A(\t$6237 ),
    .B(net1319),
    .X(booth_b52_m8));
 sky130_fd_sc_hd__a22o_1 \U$$3586  (.A1(net1507),
    .A2(net479),
    .B1(net1498),
    .B2(net752),
    .X(\t$6238 ));
 sky130_fd_sc_hd__xor2_1 \U$$3587  (.A(\t$6238 ),
    .B(net1319),
    .X(booth_b52_m9));
 sky130_fd_sc_hd__a22o_1 \U$$3588  (.A1(net1498),
    .A2(net479),
    .B1(net1222),
    .B2(net752),
    .X(\t$6239 ));
 sky130_fd_sc_hd__xor2_1 \U$$3589  (.A(\t$6239 ),
    .B(net1320),
    .X(booth_b52_m10));
 sky130_fd_sc_hd__xor2_1 \U$$359  (.A(\t$4588 ),
    .B(net1274),
    .X(booth_b4_m39));
 sky130_fd_sc_hd__a22o_1 \U$$3590  (.A1(net1222),
    .A2(net476),
    .B1(net1215),
    .B2(net749),
    .X(\t$6240 ));
 sky130_fd_sc_hd__xor2_1 \U$$3591  (.A(\t$6240 ),
    .B(net1320),
    .X(booth_b52_m11));
 sky130_fd_sc_hd__a22o_1 \U$$3592  (.A1(net1217),
    .A2(net480),
    .B1(net1208),
    .B2(net753),
    .X(\t$6241 ));
 sky130_fd_sc_hd__xor2_1 \U$$3593  (.A(\t$6241 ),
    .B(net1324),
    .X(booth_b52_m12));
 sky130_fd_sc_hd__a22o_1 \U$$3594  (.A1(net1208),
    .A2(net480),
    .B1(net1200),
    .B2(net753),
    .X(\t$6242 ));
 sky130_fd_sc_hd__xor2_1 \U$$3595  (.A(\t$6242 ),
    .B(net1324),
    .X(booth_b52_m13));
 sky130_fd_sc_hd__a22o_1 \U$$3596  (.A1(net1200),
    .A2(net480),
    .B1(net1181),
    .B2(net753),
    .X(\t$6243 ));
 sky130_fd_sc_hd__xor2_1 \U$$3597  (.A(\t$6243 ),
    .B(net1324),
    .X(booth_b52_m14));
 sky130_fd_sc_hd__a22o_1 \U$$3598  (.A1(net1181),
    .A2(net480),
    .B1(net1172),
    .B2(net753),
    .X(\t$6244 ));
 sky130_fd_sc_hd__xor2_1 \U$$3599  (.A(\t$6244 ),
    .B(net1324),
    .X(booth_b52_m15));
 sky130_fd_sc_hd__a22o_1 \U$$36  (.A1(net1175),
    .A2(net443),
    .B1(net1166),
    .B2(net685),
    .X(\t$4425 ));
 sky130_fd_sc_hd__a22o_1 \U$$360  (.A1(net940),
    .A2(net529),
    .B1(net924),
    .B2(net802),
    .X(\t$4589 ));
 sky130_fd_sc_hd__a22o_1 \U$$3600  (.A1(net1172),
    .A2(net481),
    .B1(net1163),
    .B2(net754),
    .X(\t$6245 ));
 sky130_fd_sc_hd__xor2_1 \U$$3601  (.A(\t$6245 ),
    .B(net1324),
    .X(booth_b52_m16));
 sky130_fd_sc_hd__a22o_1 \U$$3602  (.A1(net1163),
    .A2(net480),
    .B1(net1153),
    .B2(net753),
    .X(\t$6246 ));
 sky130_fd_sc_hd__xor2_1 \U$$3603  (.A(\t$6246 ),
    .B(net1324),
    .X(booth_b52_m17));
 sky130_fd_sc_hd__a22o_1 \U$$3604  (.A1(net1151),
    .A2(net479),
    .B1(net1142),
    .B2(net752),
    .X(\t$6247 ));
 sky130_fd_sc_hd__xor2_1 \U$$3605  (.A(\t$6247 ),
    .B(net1320),
    .X(booth_b52_m18));
 sky130_fd_sc_hd__a22o_1 \U$$3606  (.A1(net1142),
    .A2(net476),
    .B1(net1136),
    .B2(net749),
    .X(\t$6248 ));
 sky130_fd_sc_hd__xor2_1 \U$$3607  (.A(\t$6248 ),
    .B(net1320),
    .X(booth_b52_m19));
 sky130_fd_sc_hd__a22o_1 \U$$3608  (.A1(net1136),
    .A2(net476),
    .B1(net1120),
    .B2(net749),
    .X(\t$6249 ));
 sky130_fd_sc_hd__xor2_1 \U$$3609  (.A(\t$6249 ),
    .B(net1319),
    .X(booth_b52_m20));
 sky130_fd_sc_hd__xor2_1 \U$$361  (.A(\t$4589 ),
    .B(net1276),
    .X(booth_b4_m40));
 sky130_fd_sc_hd__a22o_1 \U$$3610  (.A1(net1120),
    .A2(net476),
    .B1(net1111),
    .B2(net749),
    .X(\t$6250 ));
 sky130_fd_sc_hd__xor2_1 \U$$3611  (.A(\t$6250 ),
    .B(net1319),
    .X(booth_b52_m21));
 sky130_fd_sc_hd__a22o_1 \U$$3612  (.A1(net1111),
    .A2(net476),
    .B1(net1102),
    .B2(net749),
    .X(\t$6251 ));
 sky130_fd_sc_hd__xor2_1 \U$$3613  (.A(\t$6251 ),
    .B(net1319),
    .X(booth_b52_m22));
 sky130_fd_sc_hd__a22o_1 \U$$3614  (.A1(net1102),
    .A2(net476),
    .B1(net1094),
    .B2(net749),
    .X(\t$6252 ));
 sky130_fd_sc_hd__xor2_1 \U$$3615  (.A(\t$6252 ),
    .B(net1319),
    .X(booth_b52_m23));
 sky130_fd_sc_hd__a22o_1 \U$$3616  (.A1(net1094),
    .A2(net476),
    .B1(net1086),
    .B2(net749),
    .X(\t$6253 ));
 sky130_fd_sc_hd__xor2_1 \U$$3617  (.A(\t$6253 ),
    .B(net1319),
    .X(booth_b52_m24));
 sky130_fd_sc_hd__a22o_1 \U$$3618  (.A1(net1085),
    .A2(net478),
    .B1(net1076),
    .B2(net751),
    .X(\t$6254 ));
 sky130_fd_sc_hd__xor2_1 \U$$3619  (.A(\t$6254 ),
    .B(net1322),
    .X(booth_b52_m25));
 sky130_fd_sc_hd__a22o_1 \U$$362  (.A1(net925),
    .A2(net530),
    .B1(net1746),
    .B2(net803),
    .X(\t$4590 ));
 sky130_fd_sc_hd__a22o_1 \U$$3620  (.A1(net1076),
    .A2(net476),
    .B1(net1068),
    .B2(net749),
    .X(\t$6255 ));
 sky130_fd_sc_hd__xor2_1 \U$$3621  (.A(\t$6255 ),
    .B(net1319),
    .X(booth_b52_m26));
 sky130_fd_sc_hd__a22o_1 \U$$3622  (.A1(net1068),
    .A2(net478),
    .B1(net1060),
    .B2(net751),
    .X(\t$6256 ));
 sky130_fd_sc_hd__xor2_1 \U$$3623  (.A(\t$6256 ),
    .B(net1322),
    .X(booth_b52_m27));
 sky130_fd_sc_hd__a22o_1 \U$$3624  (.A1(net1060),
    .A2(net477),
    .B1(net1051),
    .B2(net750),
    .X(\t$6257 ));
 sky130_fd_sc_hd__xor2_1 \U$$3625  (.A(\t$6257 ),
    .B(net1321),
    .X(booth_b52_m28));
 sky130_fd_sc_hd__a22o_1 \U$$3626  (.A1(net1052),
    .A2(net477),
    .B1(net1044),
    .B2(net750),
    .X(\t$6258 ));
 sky130_fd_sc_hd__xor2_1 \U$$3627  (.A(\t$6258 ),
    .B(net1323),
    .X(booth_b52_m29));
 sky130_fd_sc_hd__a22o_1 \U$$3628  (.A1(net1043),
    .A2(net477),
    .B1(net1027),
    .B2(net750),
    .X(\t$6259 ));
 sky130_fd_sc_hd__xor2_1 \U$$3629  (.A(\t$6259 ),
    .B(net1323),
    .X(booth_b52_m30));
 sky130_fd_sc_hd__xor2_1 \U$$363  (.A(\t$4590 ),
    .B(net1276),
    .X(booth_b4_m41));
 sky130_fd_sc_hd__a22o_1 \U$$3630  (.A1(net1028),
    .A2(net477),
    .B1(net1020),
    .B2(net750),
    .X(\t$6260 ));
 sky130_fd_sc_hd__xor2_1 \U$$3631  (.A(\t$6260 ),
    .B(net1323),
    .X(booth_b52_m31));
 sky130_fd_sc_hd__a22o_1 \U$$3632  (.A1(net1020),
    .A2(net477),
    .B1(net1003),
    .B2(net750),
    .X(\t$6261 ));
 sky130_fd_sc_hd__xor2_1 \U$$3633  (.A(\t$6261 ),
    .B(net1323),
    .X(booth_b52_m32));
 sky130_fd_sc_hd__a22o_1 \U$$3634  (.A1(net1003),
    .A2(net477),
    .B1(net995),
    .B2(net750),
    .X(\t$6262 ));
 sky130_fd_sc_hd__xor2_1 \U$$3635  (.A(\t$6262 ),
    .B(net1323),
    .X(booth_b52_m33));
 sky130_fd_sc_hd__a22o_1 \U$$3636  (.A1(net995),
    .A2(net477),
    .B1(net984),
    .B2(net750),
    .X(\t$6263 ));
 sky130_fd_sc_hd__xor2_1 \U$$3637  (.A(\t$6263 ),
    .B(net1323),
    .X(booth_b52_m34));
 sky130_fd_sc_hd__a22o_1 \U$$3638  (.A1(net985),
    .A2(net477),
    .B1(net976),
    .B2(net750),
    .X(\t$6264 ));
 sky130_fd_sc_hd__xor2_1 \U$$3639  (.A(\t$6264 ),
    .B(net1321),
    .X(booth_b52_m35));
 sky130_fd_sc_hd__a22o_1 \U$$364  (.A1(net1745),
    .A2(net529),
    .B1(net1737),
    .B2(net802),
    .X(\t$4591 ));
 sky130_fd_sc_hd__a22o_1 \U$$3640  (.A1(net979),
    .A2(net478),
    .B1(net970),
    .B2(net751),
    .X(\t$6265 ));
 sky130_fd_sc_hd__xor2_1 \U$$3641  (.A(\t$6265 ),
    .B(net1321),
    .X(booth_b52_m36));
 sky130_fd_sc_hd__a22o_1 \U$$3642  (.A1(net967),
    .A2(net478),
    .B1(net958),
    .B2(net751),
    .X(\t$6266 ));
 sky130_fd_sc_hd__xor2_1 \U$$3643  (.A(\t$6266 ),
    .B(net1322),
    .X(booth_b52_m37));
 sky130_fd_sc_hd__a22o_1 \U$$3644  (.A1(net962),
    .A2(net483),
    .B1(net954),
    .B2(net756),
    .X(\t$6267 ));
 sky130_fd_sc_hd__xor2_1 \U$$3645  (.A(\t$6267 ),
    .B(net1327),
    .X(booth_b52_m38));
 sky130_fd_sc_hd__a22o_1 \U$$3646  (.A1(net953),
    .A2(net480),
    .B1(net945),
    .B2(net753),
    .X(\t$6268 ));
 sky130_fd_sc_hd__xor2_1 \U$$3647  (.A(\t$6268 ),
    .B(net1324),
    .X(booth_b52_m39));
 sky130_fd_sc_hd__a22o_1 \U$$3648  (.A1(net945),
    .A2(net482),
    .B1(net929),
    .B2(net755),
    .X(\t$6269 ));
 sky130_fd_sc_hd__xor2_1 \U$$3649  (.A(\t$6269 ),
    .B(net1326),
    .X(booth_b52_m40));
 sky130_fd_sc_hd__xor2_1 \U$$365  (.A(\t$4591 ),
    .B(net1274),
    .X(booth_b4_m42));
 sky130_fd_sc_hd__a22o_1 \U$$3650  (.A1(net930),
    .A2(net478),
    .B1(net1751),
    .B2(net751),
    .X(\t$6270 ));
 sky130_fd_sc_hd__xor2_1 \U$$3651  (.A(\t$6270 ),
    .B(net1322),
    .X(booth_b52_m41));
 sky130_fd_sc_hd__a22o_1 \U$$3652  (.A1(net1751),
    .A2(net481),
    .B1(net1743),
    .B2(net754),
    .X(\t$6271 ));
 sky130_fd_sc_hd__xor2_1 \U$$3653  (.A(\t$6271 ),
    .B(net1325),
    .X(booth_b52_m42));
 sky130_fd_sc_hd__a22o_1 \U$$3654  (.A1(net1741),
    .A2(net480),
    .B1(net1733),
    .B2(net753),
    .X(\t$6272 ));
 sky130_fd_sc_hd__xor2_1 \U$$3655  (.A(\t$6272 ),
    .B(net1325),
    .X(booth_b52_m43));
 sky130_fd_sc_hd__a22o_1 \U$$3656  (.A1(net1734),
    .A2(net482),
    .B1(net1726),
    .B2(net755),
    .X(\t$6273 ));
 sky130_fd_sc_hd__xor2_1 \U$$3657  (.A(\t$6273 ),
    .B(net1326),
    .X(booth_b52_m44));
 sky130_fd_sc_hd__a22o_1 \U$$3658  (.A1(net1726),
    .A2(net482),
    .B1(net1717),
    .B2(net755),
    .X(\t$6274 ));
 sky130_fd_sc_hd__xor2_1 \U$$3659  (.A(\t$6274 ),
    .B(net1326),
    .X(booth_b52_m45));
 sky130_fd_sc_hd__a22o_1 \U$$366  (.A1(net1737),
    .A2(net529),
    .B1(net1729),
    .B2(net802),
    .X(\t$4592 ));
 sky130_fd_sc_hd__a22o_1 \U$$3660  (.A1(net1717),
    .A2(\sel_0$6227 ),
    .B1(net1708),
    .B2(\sel_1$6228 ),
    .X(\t$6275 ));
 sky130_fd_sc_hd__xor2_1 \U$$3661  (.A(\t$6275 ),
    .B(net1326),
    .X(booth_b52_m46));
 sky130_fd_sc_hd__a22o_1 \U$$3662  (.A1(net1708),
    .A2(net482),
    .B1(net1700),
    .B2(net755),
    .X(\t$6276 ));
 sky130_fd_sc_hd__xor2_1 \U$$3663  (.A(\t$6276 ),
    .B(net1326),
    .X(booth_b52_m47));
 sky130_fd_sc_hd__a22o_1 \U$$3664  (.A1(net1701),
    .A2(net482),
    .B1(net1694),
    .B2(net755),
    .X(\t$6277 ));
 sky130_fd_sc_hd__xor2_1 \U$$3665  (.A(\t$6277 ),
    .B(net1326),
    .X(booth_b52_m48));
 sky130_fd_sc_hd__a22o_1 \U$$3666  (.A1(net1694),
    .A2(net482),
    .B1(net1686),
    .B2(net755),
    .X(\t$6278 ));
 sky130_fd_sc_hd__xor2_1 \U$$3667  (.A(\t$6278 ),
    .B(net1326),
    .X(booth_b52_m49));
 sky130_fd_sc_hd__a22o_1 \U$$3668  (.A1(net1686),
    .A2(net482),
    .B1(net1661),
    .B2(net755),
    .X(\t$6279 ));
 sky130_fd_sc_hd__xor2_1 \U$$3669  (.A(\t$6279 ),
    .B(net1328),
    .X(booth_b52_m50));
 sky130_fd_sc_hd__xor2_1 \U$$367  (.A(\t$4592 ),
    .B(net1274),
    .X(booth_b4_m43));
 sky130_fd_sc_hd__a22o_1 \U$$3670  (.A1(net1660),
    .A2(net482),
    .B1(net1652),
    .B2(net755),
    .X(\t$6280 ));
 sky130_fd_sc_hd__xor2_1 \U$$3671  (.A(\t$6280 ),
    .B(net1326),
    .X(booth_b52_m51));
 sky130_fd_sc_hd__a22o_1 \U$$3672  (.A1(net1652),
    .A2(net482),
    .B1(net1644),
    .B2(net755),
    .X(\t$6281 ));
 sky130_fd_sc_hd__xor2_1 \U$$3673  (.A(\t$6281 ),
    .B(net1326),
    .X(booth_b52_m52));
 sky130_fd_sc_hd__a22o_1 \U$$3674  (.A1(net1644),
    .A2(net482),
    .B1(net1635),
    .B2(net755),
    .X(\t$6282 ));
 sky130_fd_sc_hd__xor2_1 \U$$3675  (.A(\t$6282 ),
    .B(net1326),
    .X(booth_b52_m53));
 sky130_fd_sc_hd__a22o_1 \U$$3676  (.A1(net1634),
    .A2(net483),
    .B1(net1624),
    .B2(net756),
    .X(\t$6283 ));
 sky130_fd_sc_hd__xor2_1 \U$$3677  (.A(\t$6283 ),
    .B(net1327),
    .X(booth_b52_m54));
 sky130_fd_sc_hd__a22o_1 \U$$3678  (.A1(net1624),
    .A2(net478),
    .B1(net1616),
    .B2(net751),
    .X(\t$6284 ));
 sky130_fd_sc_hd__xor2_1 \U$$3679  (.A(\t$6284 ),
    .B(net1322),
    .X(booth_b52_m55));
 sky130_fd_sc_hd__a22o_1 \U$$368  (.A1(net1729),
    .A2(net529),
    .B1(net1720),
    .B2(net802),
    .X(\t$4593 ));
 sky130_fd_sc_hd__a22o_1 \U$$3680  (.A1(net1616),
    .A2(net483),
    .B1(net1608),
    .B2(net756),
    .X(\t$6285 ));
 sky130_fd_sc_hd__xor2_1 \U$$3681  (.A(\t$6285 ),
    .B(net1327),
    .X(booth_b52_m56));
 sky130_fd_sc_hd__a22o_1 \U$$3682  (.A1(net1608),
    .A2(net483),
    .B1(net1600),
    .B2(net756),
    .X(\t$6286 ));
 sky130_fd_sc_hd__xor2_1 \U$$3683  (.A(\t$6286 ),
    .B(net1327),
    .X(booth_b52_m57));
 sky130_fd_sc_hd__a22o_1 \U$$3684  (.A1(net1600),
    .A2(net483),
    .B1(net1591),
    .B2(net756),
    .X(\t$6287 ));
 sky130_fd_sc_hd__xor2_1 \U$$3685  (.A(\t$6287 ),
    .B(net1327),
    .X(booth_b52_m58));
 sky130_fd_sc_hd__a22o_1 \U$$3686  (.A1(net1591),
    .A2(net483),
    .B1(net1583),
    .B2(net756),
    .X(\t$6288 ));
 sky130_fd_sc_hd__xor2_1 \U$$3687  (.A(\t$6288 ),
    .B(net1327),
    .X(booth_b52_m59));
 sky130_fd_sc_hd__a22o_1 \U$$3688  (.A1(net1583),
    .A2(net483),
    .B1(net1556),
    .B2(net756),
    .X(\t$6289 ));
 sky130_fd_sc_hd__xor2_1 \U$$3689  (.A(\t$6289 ),
    .B(net1327),
    .X(booth_b52_m60));
 sky130_fd_sc_hd__xor2_1 \U$$369  (.A(\t$4593 ),
    .B(net1274),
    .X(booth_b4_m44));
 sky130_fd_sc_hd__a22o_1 \U$$3690  (.A1(net1556),
    .A2(net483),
    .B1(net1549),
    .B2(net756),
    .X(\t$6290 ));
 sky130_fd_sc_hd__xor2_1 \U$$3691  (.A(\t$6290 ),
    .B(net1327),
    .X(booth_b52_m61));
 sky130_fd_sc_hd__a22o_1 \U$$3692  (.A1(net1549),
    .A2(net483),
    .B1(net1541),
    .B2(net756),
    .X(\t$6291 ));
 sky130_fd_sc_hd__xor2_1 \U$$3693  (.A(\t$6291 ),
    .B(net1327),
    .X(booth_b52_m62));
 sky130_fd_sc_hd__a22o_1 \U$$3694  (.A1(net1537),
    .A2(net477),
    .B1(net1529),
    .B2(net750),
    .X(\t$6292 ));
 sky130_fd_sc_hd__xor2_1 \U$$3695  (.A(\t$6292 ),
    .B(net1321),
    .X(booth_b52_m63));
 sky130_fd_sc_hd__a22o_1 \U$$3696  (.A1(net1529),
    .A2(net477),
    .B1(net1796),
    .B2(net750),
    .X(\t$6293 ));
 sky130_fd_sc_hd__xor2_1 \U$$3697  (.A(\t$6293 ),
    .B(net1321),
    .X(booth_b52_m64));
 sky130_fd_sc_hd__inv_1 \U$$3698  (.A(net1322),
    .Y(\notsign$6294 ));
 sky130_fd_sc_hd__inv_1 \U$$3699  (.A(net1321),
    .Y(\notblock$6295[0] ));
 sky130_fd_sc_hd__xor2_1 \U$$37  (.A(\t$4425 ),
    .B(net1568),
    .X(booth_b0_m15));
 sky130_fd_sc_hd__a22o_1 \U$$370  (.A1(net1724),
    .A2(net533),
    .B1(net1715),
    .B2(net806),
    .X(\t$4594 ));
 sky130_fd_sc_hd__inv_1 \U$$3700  (.A(net50),
    .Y(\notblock$6295[1] ));
 sky130_fd_sc_hd__inv_1 \U$$3701  (.A(net1301),
    .Y(\notblock$6295[2] ));
 sky130_fd_sc_hd__and2_1 \U$$3702  (.A(net1301),
    .B(\notblock$6295[1] ),
    .X(\t$6296 ));
 sky130_fd_sc_hd__a32o_2 \U$$3703  (.A1(\notblock$6295[2] ),
    .A2(net50),
    .A3(net1321),
    .B1(\t$6296 ),
    .B2(\notblock$6295[0] ),
    .X(\sel_0$6297 ));
 sky130_fd_sc_hd__xor2_4 \U$$3704  (.A(net50),
    .B(net1321),
    .X(\sel_1$6298 ));
 sky130_fd_sc_hd__a22o_1 \U$$3705  (.A1(net1797),
    .A2(net472),
    .B1(net1233),
    .B2(net745),
    .X(\t$6299 ));
 sky130_fd_sc_hd__xor2_1 \U$$3706  (.A(\t$6299 ),
    .B(net1304),
    .X(booth_b54_m0));
 sky130_fd_sc_hd__a22o_1 \U$$3707  (.A1(net1233),
    .A2(net475),
    .B1(net1129),
    .B2(net748),
    .X(\t$6300 ));
 sky130_fd_sc_hd__xor2_1 \U$$3708  (.A(\t$6300 ),
    .B(net1304),
    .X(booth_b54_m1));
 sky130_fd_sc_hd__a22o_1 \U$$3709  (.A1(net1129),
    .A2(net472),
    .B1(net1037),
    .B2(net745),
    .X(\t$6301 ));
 sky130_fd_sc_hd__xor2_1 \U$$371  (.A(\t$4594 ),
    .B(net1279),
    .X(booth_b4_m45));
 sky130_fd_sc_hd__xor2_1 \U$$3710  (.A(\t$6301 ),
    .B(net1305),
    .X(booth_b54_m2));
 sky130_fd_sc_hd__a22o_1 \U$$3711  (.A1(net1037),
    .A2(net472),
    .B1(net938),
    .B2(net745),
    .X(\t$6302 ));
 sky130_fd_sc_hd__xor2_1 \U$$3712  (.A(\t$6302 ),
    .B(net1305),
    .X(booth_b54_m3));
 sky130_fd_sc_hd__a22o_1 \U$$3713  (.A1(net938),
    .A2(net472),
    .B1(net1677),
    .B2(net745),
    .X(\t$6303 ));
 sky130_fd_sc_hd__xor2_1 \U$$3714  (.A(\t$6303 ),
    .B(net1305),
    .X(booth_b54_m4));
 sky130_fd_sc_hd__a22o_1 \U$$3715  (.A1(net1674),
    .A2(net468),
    .B1(net1563),
    .B2(net741),
    .X(\t$6304 ));
 sky130_fd_sc_hd__xor2_1 \U$$3716  (.A(\t$6304 ),
    .B(net1300),
    .X(booth_b54_m5));
 sky130_fd_sc_hd__a22o_1 \U$$3717  (.A1(net1563),
    .A2(net468),
    .B1(net1522),
    .B2(net741),
    .X(\t$6305 ));
 sky130_fd_sc_hd__xor2_1 \U$$3718  (.A(\t$6305 ),
    .B(net1300),
    .X(booth_b54_m6));
 sky130_fd_sc_hd__a22o_1 \U$$3719  (.A1(net1522),
    .A2(net471),
    .B1(net1514),
    .B2(net744),
    .X(\t$6306 ));
 sky130_fd_sc_hd__a22o_1 \U$$372  (.A1(net1711),
    .A2(net529),
    .B1(net1703),
    .B2(net802),
    .X(\t$4595 ));
 sky130_fd_sc_hd__xor2_1 \U$$3720  (.A(\t$6306 ),
    .B(net1300),
    .X(booth_b54_m7));
 sky130_fd_sc_hd__a22o_1 \U$$3721  (.A1(net1514),
    .A2(net471),
    .B1(net1507),
    .B2(net744),
    .X(\t$6307 ));
 sky130_fd_sc_hd__xor2_1 \U$$3722  (.A(\t$6307 ),
    .B(net1309),
    .X(booth_b54_m8));
 sky130_fd_sc_hd__a22o_1 \U$$3723  (.A1(net1507),
    .A2(net468),
    .B1(net1498),
    .B2(net741),
    .X(\t$6308 ));
 sky130_fd_sc_hd__xor2_1 \U$$3724  (.A(\t$6308 ),
    .B(net1300),
    .X(booth_b54_m9));
 sky130_fd_sc_hd__a22o_1 \U$$3725  (.A1(net1501),
    .A2(net472),
    .B1(net1226),
    .B2(net745),
    .X(\t$6309 ));
 sky130_fd_sc_hd__xor2_1 \U$$3726  (.A(\t$6309 ),
    .B(net1304),
    .X(booth_b54_m10));
 sky130_fd_sc_hd__a22o_1 \U$$3727  (.A1(net1226),
    .A2(net475),
    .B1(net1217),
    .B2(net748),
    .X(\t$6310 ));
 sky130_fd_sc_hd__xor2_1 \U$$3728  (.A(\t$6310 ),
    .B(net1304),
    .X(booth_b54_m11));
 sky130_fd_sc_hd__a22o_1 \U$$3729  (.A1(net1217),
    .A2(net472),
    .B1(net1208),
    .B2(net745),
    .X(\t$6311 ));
 sky130_fd_sc_hd__xor2_1 \U$$373  (.A(\t$4595 ),
    .B(net1275),
    .X(booth_b4_m46));
 sky130_fd_sc_hd__xor2_1 \U$$3730  (.A(\t$6311 ),
    .B(net1304),
    .X(booth_b54_m12));
 sky130_fd_sc_hd__a22o_1 \U$$3731  (.A1(net1208),
    .A2(net472),
    .B1(net1200),
    .B2(net745),
    .X(\t$6312 ));
 sky130_fd_sc_hd__xor2_1 \U$$3732  (.A(\t$6312 ),
    .B(net1304),
    .X(booth_b54_m13));
 sky130_fd_sc_hd__a22o_1 \U$$3733  (.A1(net1200),
    .A2(net475),
    .B1(net1181),
    .B2(net748),
    .X(\t$6313 ));
 sky130_fd_sc_hd__xor2_1 \U$$3734  (.A(\t$6313 ),
    .B(net1304),
    .X(booth_b54_m14));
 sky130_fd_sc_hd__a22o_1 \U$$3735  (.A1(net1182),
    .A2(net475),
    .B1(net1172),
    .B2(net748),
    .X(\t$6314 ));
 sky130_fd_sc_hd__xor2_1 \U$$3736  (.A(\t$6314 ),
    .B(net1304),
    .X(booth_b54_m15));
 sky130_fd_sc_hd__a22o_1 \U$$3737  (.A1(net1169),
    .A2(net468),
    .B1(net1160),
    .B2(net741),
    .X(\t$6315 ));
 sky130_fd_sc_hd__xor2_1 \U$$3738  (.A(\t$6315 ),
    .B(net1309),
    .X(booth_b54_m16));
 sky130_fd_sc_hd__a22o_1 \U$$3739  (.A1(net1160),
    .A2(net470),
    .B1(net1151),
    .B2(net743),
    .X(\t$6316 ));
 sky130_fd_sc_hd__a22o_1 \U$$374  (.A1(net1706),
    .A2(net533),
    .B1(net1699),
    .B2(net806),
    .X(\t$4596 ));
 sky130_fd_sc_hd__xor2_1 \U$$3740  (.A(\t$6316 ),
    .B(net1301),
    .X(booth_b54_m17));
 sky130_fd_sc_hd__a22o_1 \U$$3741  (.A1(net1151),
    .A2(net468),
    .B1(net1141),
    .B2(net741),
    .X(\t$6317 ));
 sky130_fd_sc_hd__xor2_1 \U$$3742  (.A(\t$6317 ),
    .B(net1300),
    .X(booth_b54_m18));
 sky130_fd_sc_hd__a22o_1 \U$$3743  (.A1(net1141),
    .A2(net468),
    .B1(net1136),
    .B2(net741),
    .X(\t$6318 ));
 sky130_fd_sc_hd__xor2_1 \U$$3744  (.A(\t$6318 ),
    .B(net1300),
    .X(booth_b54_m19));
 sky130_fd_sc_hd__a22o_1 \U$$3745  (.A1(net1136),
    .A2(net468),
    .B1(net1120),
    .B2(net741),
    .X(\t$6319 ));
 sky130_fd_sc_hd__xor2_1 \U$$3746  (.A(\t$6319 ),
    .B(net1300),
    .X(booth_b54_m20));
 sky130_fd_sc_hd__a22o_1 \U$$3747  (.A1(net1120),
    .A2(net468),
    .B1(net1111),
    .B2(net741),
    .X(\t$6320 ));
 sky130_fd_sc_hd__xor2_1 \U$$3748  (.A(\t$6320 ),
    .B(net1300),
    .X(booth_b54_m21));
 sky130_fd_sc_hd__a22o_1 \U$$3749  (.A1(net1111),
    .A2(net468),
    .B1(net1102),
    .B2(net741),
    .X(\t$6321 ));
 sky130_fd_sc_hd__xor2_1 \U$$375  (.A(\t$4596 ),
    .B(net1278),
    .X(booth_b4_m47));
 sky130_fd_sc_hd__xor2_1 \U$$3750  (.A(\t$6321 ),
    .B(net1300),
    .X(booth_b54_m22));
 sky130_fd_sc_hd__a22o_1 \U$$3751  (.A1(net1102),
    .A2(net470),
    .B1(net1094),
    .B2(net743),
    .X(\t$6322 ));
 sky130_fd_sc_hd__xor2_1 \U$$3752  (.A(\t$6322 ),
    .B(net1301),
    .X(booth_b54_m23));
 sky130_fd_sc_hd__a22o_1 \U$$3753  (.A1(net1094),
    .A2(net468),
    .B1(net1086),
    .B2(net741),
    .X(\t$6323 ));
 sky130_fd_sc_hd__xor2_1 \U$$3754  (.A(\t$6323 ),
    .B(net1300),
    .X(booth_b54_m24));
 sky130_fd_sc_hd__a22o_1 \U$$3755  (.A1(net1085),
    .A2(net470),
    .B1(net1076),
    .B2(net743),
    .X(\t$6324 ));
 sky130_fd_sc_hd__xor2_1 \U$$3756  (.A(\t$6324 ),
    .B(net1301),
    .X(booth_b54_m25));
 sky130_fd_sc_hd__a22o_1 \U$$3757  (.A1(net1077),
    .A2(net469),
    .B1(net1068),
    .B2(net742),
    .X(\t$6325 ));
 sky130_fd_sc_hd__xor2_1 \U$$3758  (.A(\t$6325 ),
    .B(net1303),
    .X(booth_b54_m26));
 sky130_fd_sc_hd__a22o_1 \U$$3759  (.A1(net1069),
    .A2(net469),
    .B1(net1061),
    .B2(net742),
    .X(\t$6326 ));
 sky130_fd_sc_hd__a22o_1 \U$$376  (.A1(net1699),
    .A2(net533),
    .B1(net1690),
    .B2(net806),
    .X(\t$4597 ));
 sky130_fd_sc_hd__xor2_1 \U$$3760  (.A(\t$6326 ),
    .B(net1303),
    .X(booth_b54_m27));
 sky130_fd_sc_hd__a22o_1 \U$$3761  (.A1(net1060),
    .A2(net469),
    .B1(net1051),
    .B2(net742),
    .X(\t$6327 ));
 sky130_fd_sc_hd__xor2_1 \U$$3762  (.A(\t$6327 ),
    .B(net1303),
    .X(booth_b54_m28));
 sky130_fd_sc_hd__a22o_1 \U$$3763  (.A1(net1052),
    .A2(net469),
    .B1(net1044),
    .B2(net742),
    .X(\t$6328 ));
 sky130_fd_sc_hd__xor2_1 \U$$3764  (.A(\t$6328 ),
    .B(net1303),
    .X(booth_b54_m29));
 sky130_fd_sc_hd__a22o_1 \U$$3765  (.A1(net1044),
    .A2(net469),
    .B1(net1028),
    .B2(net742),
    .X(\t$6329 ));
 sky130_fd_sc_hd__xor2_1 \U$$3766  (.A(\t$6329 ),
    .B(net1303),
    .X(booth_b54_m30));
 sky130_fd_sc_hd__a22o_1 \U$$3767  (.A1(net1028),
    .A2(net469),
    .B1(net1020),
    .B2(net742),
    .X(\t$6330 ));
 sky130_fd_sc_hd__xor2_1 \U$$3768  (.A(\t$6330 ),
    .B(net1303),
    .X(booth_b54_m31));
 sky130_fd_sc_hd__a22o_1 \U$$3769  (.A1(net1020),
    .A2(net469),
    .B1(net1003),
    .B2(net742),
    .X(\t$6331 ));
 sky130_fd_sc_hd__xor2_1 \U$$377  (.A(\t$4597 ),
    .B(net1278),
    .X(booth_b4_m48));
 sky130_fd_sc_hd__xor2_1 \U$$3770  (.A(\t$6331 ),
    .B(net1303),
    .X(booth_b54_m32));
 sky130_fd_sc_hd__a22o_1 \U$$3771  (.A1(net1003),
    .A2(net469),
    .B1(net995),
    .B2(net742),
    .X(\t$6332 ));
 sky130_fd_sc_hd__xor2_1 \U$$3772  (.A(\t$6332 ),
    .B(net1301),
    .X(booth_b54_m33));
 sky130_fd_sc_hd__a22o_1 \U$$3773  (.A1(net997),
    .A2(net470),
    .B1(net988),
    .B2(net743),
    .X(\t$6333 ));
 sky130_fd_sc_hd__xor2_1 \U$$3774  (.A(\t$6333 ),
    .B(net1301),
    .X(booth_b54_m34));
 sky130_fd_sc_hd__a22o_1 \U$$3775  (.A1(net985),
    .A2(net470),
    .B1(net976),
    .B2(net743),
    .X(\t$6334 ));
 sky130_fd_sc_hd__xor2_1 \U$$3776  (.A(\t$6334 ),
    .B(net1301),
    .X(booth_b54_m35));
 sky130_fd_sc_hd__a22o_1 \U$$3777  (.A1(net979),
    .A2(net473),
    .B1(net970),
    .B2(net746),
    .X(\t$6335 ));
 sky130_fd_sc_hd__xor2_1 \U$$3778  (.A(\t$6335 ),
    .B(net1306),
    .X(booth_b54_m36));
 sky130_fd_sc_hd__a22o_1 \U$$3779  (.A1(net970),
    .A2(net472),
    .B1(net962),
    .B2(net745),
    .X(\t$6336 ));
 sky130_fd_sc_hd__a22o_1 \U$$378  (.A1(net1691),
    .A2(net533),
    .B1(net1682),
    .B2(net806),
    .X(\t$4598 ));
 sky130_fd_sc_hd__xor2_1 \U$$3780  (.A(\t$6336 ),
    .B(net1304),
    .X(booth_b54_m37));
 sky130_fd_sc_hd__a22o_1 \U$$3781  (.A1(net962),
    .A2(net474),
    .B1(net953),
    .B2(net747),
    .X(\t$6337 ));
 sky130_fd_sc_hd__xor2_1 \U$$3782  (.A(\t$6337 ),
    .B(net1307),
    .X(booth_b54_m38));
 sky130_fd_sc_hd__a22o_1 \U$$3783  (.A1(net954),
    .A2(net470),
    .B1(net946),
    .B2(net743),
    .X(\t$6338 ));
 sky130_fd_sc_hd__xor2_1 \U$$3784  (.A(\t$6338 ),
    .B(net1301),
    .X(booth_b54_m39));
 sky130_fd_sc_hd__a22o_1 \U$$3785  (.A1(net946),
    .A2(net472),
    .B1(net930),
    .B2(net745),
    .X(\t$6339 ));
 sky130_fd_sc_hd__xor2_1 \U$$3786  (.A(\t$6339 ),
    .B(net1305),
    .X(booth_b54_m40));
 sky130_fd_sc_hd__a22o_1 \U$$3787  (.A1(net928),
    .A2(net472),
    .B1(net1749),
    .B2(net745),
    .X(\t$6340 ));
 sky130_fd_sc_hd__xor2_1 \U$$3788  (.A(\t$6340 ),
    .B(net1305),
    .X(booth_b54_m41));
 sky130_fd_sc_hd__a22o_1 \U$$3789  (.A1(net1750),
    .A2(net474),
    .B1(net1742),
    .B2(net747),
    .X(\t$6341 ));
 sky130_fd_sc_hd__xor2_1 \U$$379  (.A(\t$4598 ),
    .B(net1280),
    .X(booth_b4_m49));
 sky130_fd_sc_hd__xor2_1 \U$$3790  (.A(\t$6341 ),
    .B(net1307),
    .X(booth_b54_m42));
 sky130_fd_sc_hd__a22o_1 \U$$3791  (.A1(net1742),
    .A2(net474),
    .B1(net1734),
    .B2(net747),
    .X(\t$6342 ));
 sky130_fd_sc_hd__xor2_1 \U$$3792  (.A(\t$6342 ),
    .B(net1307),
    .X(booth_b54_m43));
 sky130_fd_sc_hd__a22o_1 \U$$3793  (.A1(net1734),
    .A2(net475),
    .B1(net1726),
    .B2(net748),
    .X(\t$6343 ));
 sky130_fd_sc_hd__xor2_1 \U$$3794  (.A(\t$6343 ),
    .B(net1307),
    .X(booth_b54_m44));
 sky130_fd_sc_hd__a22o_1 \U$$3795  (.A1(net1726),
    .A2(net474),
    .B1(net1717),
    .B2(net747),
    .X(\t$6344 ));
 sky130_fd_sc_hd__xor2_1 \U$$3796  (.A(\t$6344 ),
    .B(net1307),
    .X(booth_b54_m45));
 sky130_fd_sc_hd__a22o_1 \U$$3797  (.A1(net1718),
    .A2(net474),
    .B1(net1709),
    .B2(net747),
    .X(\t$6345 ));
 sky130_fd_sc_hd__xor2_1 \U$$3798  (.A(\t$6345 ),
    .B(net1307),
    .X(booth_b54_m46));
 sky130_fd_sc_hd__a22o_1 \U$$3799  (.A1(net1709),
    .A2(net474),
    .B1(net1701),
    .B2(net747),
    .X(\t$6346 ));
 sky130_fd_sc_hd__a22o_1 \U$$38  (.A1(net1166),
    .A2(net443),
    .B1(net1157),
    .B2(net685),
    .X(\t$4426 ));
 sky130_fd_sc_hd__a22o_1 \U$$380  (.A1(net1683),
    .A2(net534),
    .B1(net1658),
    .B2(net807),
    .X(\t$4599 ));
 sky130_fd_sc_hd__xor2_1 \U$$3800  (.A(\t$6346 ),
    .B(net1307),
    .X(booth_b54_m47));
 sky130_fd_sc_hd__a22o_1 \U$$3801  (.A1(net1701),
    .A2(net474),
    .B1(net1694),
    .B2(net747),
    .X(\t$6347 ));
 sky130_fd_sc_hd__xor2_1 \U$$3802  (.A(\t$6347 ),
    .B(net1307),
    .X(booth_b54_m48));
 sky130_fd_sc_hd__a22o_1 \U$$3803  (.A1(net1693),
    .A2(net474),
    .B1(net1684),
    .B2(net747),
    .X(\t$6348 ));
 sky130_fd_sc_hd__xor2_1 \U$$3804  (.A(\t$6348 ),
    .B(net1307),
    .X(booth_b54_m49));
 sky130_fd_sc_hd__a22o_1 \U$$3805  (.A1(net1686),
    .A2(net474),
    .B1(net1661),
    .B2(net747),
    .X(\t$6349 ));
 sky130_fd_sc_hd__xor2_1 \U$$3806  (.A(\t$6349 ),
    .B(net1308),
    .X(booth_b54_m50));
 sky130_fd_sc_hd__a22o_1 \U$$3807  (.A1(net1660),
    .A2(net474),
    .B1(net1652),
    .B2(net747),
    .X(\t$6350 ));
 sky130_fd_sc_hd__xor2_1 \U$$3808  (.A(\t$6350 ),
    .B(net1307),
    .X(booth_b54_m51));
 sky130_fd_sc_hd__a22o_1 \U$$3809  (.A1(net1651),
    .A2(net473),
    .B1(net1643),
    .B2(net746),
    .X(\t$6351 ));
 sky130_fd_sc_hd__xor2_1 \U$$381  (.A(\t$4599 ),
    .B(net1280),
    .X(booth_b4_m50));
 sky130_fd_sc_hd__xor2_1 \U$$3810  (.A(\t$6351 ),
    .B(net1306),
    .X(booth_b54_m52));
 sky130_fd_sc_hd__a22o_1 \U$$3811  (.A1(net1643),
    .A2(net470),
    .B1(net1634),
    .B2(net743),
    .X(\t$6352 ));
 sky130_fd_sc_hd__xor2_1 \U$$3812  (.A(\t$6352 ),
    .B(net1301),
    .X(booth_b54_m53));
 sky130_fd_sc_hd__a22o_1 \U$$3813  (.A1(net1634),
    .A2(net473),
    .B1(net1624),
    .B2(net746),
    .X(\t$6353 ));
 sky130_fd_sc_hd__xor2_1 \U$$3814  (.A(\t$6353 ),
    .B(net1306),
    .X(booth_b54_m54));
 sky130_fd_sc_hd__a22o_1 \U$$3815  (.A1(net1624),
    .A2(net473),
    .B1(net1616),
    .B2(net746),
    .X(\t$6354 ));
 sky130_fd_sc_hd__xor2_1 \U$$3816  (.A(\t$6354 ),
    .B(net1306),
    .X(booth_b54_m55));
 sky130_fd_sc_hd__a22o_1 \U$$3817  (.A1(net1616),
    .A2(net473),
    .B1(net1608),
    .B2(net746),
    .X(\t$6355 ));
 sky130_fd_sc_hd__xor2_1 \U$$3818  (.A(\t$6355 ),
    .B(net1306),
    .X(booth_b54_m56));
 sky130_fd_sc_hd__a22o_1 \U$$3819  (.A1(net1608),
    .A2(net473),
    .B1(net1600),
    .B2(net746),
    .X(\t$6356 ));
 sky130_fd_sc_hd__a22o_1 \U$$382  (.A1(net1658),
    .A2(net533),
    .B1(net1650),
    .B2(net806),
    .X(\t$4600 ));
 sky130_fd_sc_hd__xor2_1 \U$$3820  (.A(\t$6356 ),
    .B(net1306),
    .X(booth_b54_m57));
 sky130_fd_sc_hd__a22o_1 \U$$3821  (.A1(net1600),
    .A2(net473),
    .B1(net1591),
    .B2(net746),
    .X(\t$6357 ));
 sky130_fd_sc_hd__xor2_1 \U$$3822  (.A(\t$6357 ),
    .B(net1306),
    .X(booth_b54_m58));
 sky130_fd_sc_hd__a22o_1 \U$$3823  (.A1(net1591),
    .A2(net473),
    .B1(net1583),
    .B2(net746),
    .X(\t$6358 ));
 sky130_fd_sc_hd__xor2_1 \U$$3824  (.A(\t$6358 ),
    .B(net1306),
    .X(booth_b54_m59));
 sky130_fd_sc_hd__a22o_1 \U$$3825  (.A1(net1583),
    .A2(net473),
    .B1(net1556),
    .B2(net746),
    .X(\t$6359 ));
 sky130_fd_sc_hd__xor2_1 \U$$3826  (.A(\t$6359 ),
    .B(net1306),
    .X(booth_b54_m60));
 sky130_fd_sc_hd__a22o_1 \U$$3827  (.A1(net1554),
    .A2(net469),
    .B1(net1545),
    .B2(net742),
    .X(\t$6360 ));
 sky130_fd_sc_hd__xor2_1 \U$$3828  (.A(\t$6360 ),
    .B(net1302),
    .X(booth_b54_m61));
 sky130_fd_sc_hd__a22o_1 \U$$3829  (.A1(net1549),
    .A2(net473),
    .B1(net1541),
    .B2(net746),
    .X(\t$6361 ));
 sky130_fd_sc_hd__xor2_1 \U$$383  (.A(\t$4600 ),
    .B(net1280),
    .X(booth_b4_m51));
 sky130_fd_sc_hd__xor2_1 \U$$3830  (.A(\t$6361 ),
    .B(net1306),
    .X(booth_b54_m62));
 sky130_fd_sc_hd__a22o_1 \U$$3831  (.A1(net1537),
    .A2(net469),
    .B1(net1529),
    .B2(net742),
    .X(\t$6362 ));
 sky130_fd_sc_hd__xor2_1 \U$$3832  (.A(\t$6362 ),
    .B(net1302),
    .X(booth_b54_m63));
 sky130_fd_sc_hd__a22o_1 \U$$3833  (.A1(net1533),
    .A2(net475),
    .B1(net1798),
    .B2(net748),
    .X(\t$6363 ));
 sky130_fd_sc_hd__xor2_1 \U$$3834  (.A(\t$6363 ),
    .B(net1308),
    .X(booth_b54_m64));
 sky130_fd_sc_hd__inv_1 \U$$3835  (.A(net1302),
    .Y(\notsign$6364 ));
 sky130_fd_sc_hd__inv_1 \U$$3836  (.A(net1302),
    .Y(\notblock$6365[0] ));
 sky130_fd_sc_hd__inv_1 \U$$3837  (.A(net52),
    .Y(\notblock$6365[1] ));
 sky130_fd_sc_hd__inv_1 \U$$3838  (.A(net1292),
    .Y(\notblock$6365[2] ));
 sky130_fd_sc_hd__and2_1 \U$$3839  (.A(net1292),
    .B(\notblock$6365[1] ),
    .X(\t$6366 ));
 sky130_fd_sc_hd__a22o_1 \U$$384  (.A1(net1649),
    .A2(net534),
    .B1(net1641),
    .B2(net807),
    .X(\t$4601 ));
 sky130_fd_sc_hd__a32o_4 \U$$3840  (.A1(\notblock$6365[2] ),
    .A2(net52),
    .A3(net1302),
    .B1(\t$6366 ),
    .B2(\notblock$6365[0] ),
    .X(\sel_0$6367 ));
 sky130_fd_sc_hd__xor2_4 \U$$3841  (.A(net52),
    .B(net1302),
    .X(\sel_1$6368 ));
 sky130_fd_sc_hd__a22o_1 \U$$3842  (.A1(net1799),
    .A2(net464),
    .B1(net1233),
    .B2(net737),
    .X(\t$6369 ));
 sky130_fd_sc_hd__xor2_1 \U$$3843  (.A(\t$6369 ),
    .B(net1296),
    .X(booth_b56_m0));
 sky130_fd_sc_hd__a22o_1 \U$$3844  (.A1(net1233),
    .A2(net464),
    .B1(net1129),
    .B2(net737),
    .X(\t$6370 ));
 sky130_fd_sc_hd__xor2_1 \U$$3845  (.A(\t$6370 ),
    .B(net1296),
    .X(booth_b56_m1));
 sky130_fd_sc_hd__a22o_1 \U$$3846  (.A1(net1129),
    .A2(net464),
    .B1(net1037),
    .B2(net737),
    .X(\t$6371 ));
 sky130_fd_sc_hd__xor2_1 \U$$3847  (.A(\t$6371 ),
    .B(net1296),
    .X(booth_b56_m2));
 sky130_fd_sc_hd__a22o_1 \U$$3848  (.A1(net1037),
    .A2(net461),
    .B1(net935),
    .B2(net734),
    .X(\t$6372 ));
 sky130_fd_sc_hd__xor2_1 \U$$3849  (.A(\t$6372 ),
    .B(net1291),
    .X(booth_b56_m3));
 sky130_fd_sc_hd__xor2_1 \U$$385  (.A(\t$4601 ),
    .B(net1280),
    .X(booth_b4_m52));
 sky130_fd_sc_hd__a22o_1 \U$$3850  (.A1(net935),
    .A2(net460),
    .B1(net1674),
    .B2(net733),
    .X(\t$6373 ));
 sky130_fd_sc_hd__xor2_1 \U$$3851  (.A(\t$6373 ),
    .B(net1291),
    .X(booth_b56_m4));
 sky130_fd_sc_hd__a22o_1 \U$$3852  (.A1(net1674),
    .A2(net461),
    .B1(net1563),
    .B2(net734),
    .X(\t$6374 ));
 sky130_fd_sc_hd__xor2_1 \U$$3853  (.A(\t$6374 ),
    .B(net1291),
    .X(booth_b56_m5));
 sky130_fd_sc_hd__a22o_1 \U$$3854  (.A1(net1563),
    .A2(net461),
    .B1(net1522),
    .B2(net734),
    .X(\t$6375 ));
 sky130_fd_sc_hd__xor2_1 \U$$3855  (.A(\t$6375 ),
    .B(net1295),
    .X(booth_b56_m6));
 sky130_fd_sc_hd__a22o_1 \U$$3856  (.A1(net1522),
    .A2(net460),
    .B1(net1518),
    .B2(net733),
    .X(\t$6376 ));
 sky130_fd_sc_hd__xor2_1 \U$$3857  (.A(\t$6376 ),
    .B(net1291),
    .X(booth_b56_m7));
 sky130_fd_sc_hd__a22o_1 \U$$3858  (.A1(net1517),
    .A2(net467),
    .B1(net1510),
    .B2(net740),
    .X(\t$6377 ));
 sky130_fd_sc_hd__xor2_1 \U$$3859  (.A(\t$6377 ),
    .B(net1296),
    .X(booth_b56_m8));
 sky130_fd_sc_hd__a22o_1 \U$$386  (.A1(net1641),
    .A2(net533),
    .B1(net1633),
    .B2(net806),
    .X(\t$4602 ));
 sky130_fd_sc_hd__a22o_1 \U$$3860  (.A1(net1510),
    .A2(net464),
    .B1(net1501),
    .B2(net737),
    .X(\t$6378 ));
 sky130_fd_sc_hd__xor2_1 \U$$3861  (.A(\t$6378 ),
    .B(net1296),
    .X(booth_b56_m9));
 sky130_fd_sc_hd__a22o_1 \U$$3862  (.A1(net1501),
    .A2(net467),
    .B1(net1226),
    .B2(net740),
    .X(\t$6379 ));
 sky130_fd_sc_hd__xor2_1 \U$$3863  (.A(\t$6379 ),
    .B(net1296),
    .X(booth_b56_m10));
 sky130_fd_sc_hd__a22o_1 \U$$3864  (.A1(net1226),
    .A2(net467),
    .B1(net1217),
    .B2(net740),
    .X(\t$6380 ));
 sky130_fd_sc_hd__xor2_1 \U$$3865  (.A(\t$6380 ),
    .B(net1296),
    .X(booth_b56_m11));
 sky130_fd_sc_hd__a22o_1 \U$$3866  (.A1(net1217),
    .A2(net464),
    .B1(net1208),
    .B2(net737),
    .X(\t$6381 ));
 sky130_fd_sc_hd__xor2_1 \U$$3867  (.A(\t$6381 ),
    .B(net1296),
    .X(booth_b56_m12));
 sky130_fd_sc_hd__a22o_1 \U$$3868  (.A1(net1208),
    .A2(net464),
    .B1(net1200),
    .B2(net737),
    .X(\t$6382 ));
 sky130_fd_sc_hd__xor2_1 \U$$3869  (.A(\t$6382 ),
    .B(net1299),
    .X(booth_b56_m13));
 sky130_fd_sc_hd__xor2_1 \U$$387  (.A(\t$4602 ),
    .B(net1280),
    .X(booth_b4_m53));
 sky130_fd_sc_hd__a22o_1 \U$$3870  (.A1(net1197),
    .A2(net460),
    .B1(net1178),
    .B2(net733),
    .X(\t$6383 ));
 sky130_fd_sc_hd__xor2_1 \U$$3871  (.A(\t$6383 ),
    .B(net1295),
    .X(booth_b56_m14));
 sky130_fd_sc_hd__a22o_1 \U$$3872  (.A1(net1178),
    .A2(net461),
    .B1(net1169),
    .B2(net734),
    .X(\t$6384 ));
 sky130_fd_sc_hd__xor2_1 \U$$3873  (.A(\t$6384 ),
    .B(net1295),
    .X(booth_b56_m15));
 sky130_fd_sc_hd__a22o_1 \U$$3874  (.A1(net1168),
    .A2(net460),
    .B1(net1159),
    .B2(net733),
    .X(\t$6385 ));
 sky130_fd_sc_hd__xor2_1 \U$$3875  (.A(\t$6385 ),
    .B(net1291),
    .X(booth_b56_m16));
 sky130_fd_sc_hd__a22o_1 \U$$3876  (.A1(net1159),
    .A2(net460),
    .B1(net1151),
    .B2(net733),
    .X(\t$6386 ));
 sky130_fd_sc_hd__xor2_1 \U$$3877  (.A(\t$6386 ),
    .B(net1291),
    .X(booth_b56_m17));
 sky130_fd_sc_hd__a22o_1 \U$$3878  (.A1(net1151),
    .A2(net460),
    .B1(net1141),
    .B2(net733),
    .X(\t$6387 ));
 sky130_fd_sc_hd__xor2_1 \U$$3879  (.A(\t$6387 ),
    .B(net1291),
    .X(booth_b56_m18));
 sky130_fd_sc_hd__a22o_1 \U$$388  (.A1(net1633),
    .A2(net533),
    .B1(net1623),
    .B2(net806),
    .X(\t$4603 ));
 sky130_fd_sc_hd__a22o_1 \U$$3880  (.A1(net1141),
    .A2(net460),
    .B1(net1136),
    .B2(net733),
    .X(\t$6388 ));
 sky130_fd_sc_hd__xor2_1 \U$$3881  (.A(\t$6388 ),
    .B(net1291),
    .X(booth_b56_m19));
 sky130_fd_sc_hd__a22o_1 \U$$3882  (.A1(net1135),
    .A2(net460),
    .B1(net1119),
    .B2(net733),
    .X(\t$6389 ));
 sky130_fd_sc_hd__xor2_1 \U$$3883  (.A(\t$6389 ),
    .B(net1291),
    .X(booth_b56_m20));
 sky130_fd_sc_hd__a22o_1 \U$$3884  (.A1(net1119),
    .A2(net460),
    .B1(net1111),
    .B2(net733),
    .X(\t$6390 ));
 sky130_fd_sc_hd__xor2_1 \U$$3885  (.A(\t$6390 ),
    .B(net1294),
    .X(booth_b56_m21));
 sky130_fd_sc_hd__a22o_1 \U$$3886  (.A1(net1111),
    .A2(net461),
    .B1(net1102),
    .B2(net734),
    .X(\t$6391 ));
 sky130_fd_sc_hd__xor2_1 \U$$3887  (.A(\t$6391 ),
    .B(net1291),
    .X(booth_b56_m22));
 sky130_fd_sc_hd__a22o_1 \U$$3888  (.A1(net1102),
    .A2(net463),
    .B1(net1094),
    .B2(net736),
    .X(\t$6392 ));
 sky130_fd_sc_hd__xor2_1 \U$$3889  (.A(\t$6392 ),
    .B(net1294),
    .X(booth_b56_m23));
 sky130_fd_sc_hd__xor2_1 \U$$389  (.A(\t$4603 ),
    .B(net1280),
    .X(booth_b4_m54));
 sky130_fd_sc_hd__a22o_1 \U$$3890  (.A1(net1094),
    .A2(net462),
    .B1(net1085),
    .B2(net735),
    .X(\t$6393 ));
 sky130_fd_sc_hd__xor2_1 \U$$3891  (.A(\t$6393 ),
    .B(net1292),
    .X(booth_b56_m24));
 sky130_fd_sc_hd__a22o_1 \U$$3892  (.A1(net1085),
    .A2(net463),
    .B1(net1077),
    .B2(net736),
    .X(\t$6394 ));
 sky130_fd_sc_hd__xor2_1 \U$$3893  (.A(\t$6394 ),
    .B(net1294),
    .X(booth_b56_m25));
 sky130_fd_sc_hd__a22o_1 \U$$3894  (.A1(net1076),
    .A2(net460),
    .B1(net1068),
    .B2(net733),
    .X(\t$6395 ));
 sky130_fd_sc_hd__xor2_1 \U$$3895  (.A(\t$6395 ),
    .B(net1294),
    .X(booth_b56_m26));
 sky130_fd_sc_hd__a22o_1 \U$$3896  (.A1(net1069),
    .A2(net463),
    .B1(net1061),
    .B2(net736),
    .X(\t$6396 ));
 sky130_fd_sc_hd__xor2_1 \U$$3897  (.A(\t$6396 ),
    .B(net1294),
    .X(booth_b56_m27));
 sky130_fd_sc_hd__a22o_1 \U$$3898  (.A1(net1061),
    .A2(net463),
    .B1(net1052),
    .B2(net736),
    .X(\t$6397 ));
 sky130_fd_sc_hd__xor2_1 \U$$3899  (.A(\t$6397 ),
    .B(net1294),
    .X(booth_b56_m28));
 sky130_fd_sc_hd__xor2_1 \U$$39  (.A(\t$4426 ),
    .B(net1568),
    .X(booth_b0_m16));
 sky130_fd_sc_hd__a22o_1 \U$$390  (.A1(net1620),
    .A2(net530),
    .B1(net1612),
    .B2(net803),
    .X(\t$4604 ));
 sky130_fd_sc_hd__a22o_1 \U$$3900  (.A1(net1052),
    .A2(net463),
    .B1(net1044),
    .B2(net736),
    .X(\t$6398 ));
 sky130_fd_sc_hd__xor2_1 \U$$3901  (.A(\t$6398 ),
    .B(net1294),
    .X(booth_b56_m29));
 sky130_fd_sc_hd__a22o_1 \U$$3902  (.A1(net1044),
    .A2(net463),
    .B1(net1028),
    .B2(net736),
    .X(\t$6399 ));
 sky130_fd_sc_hd__xor2_1 \U$$3903  (.A(\t$6399 ),
    .B(net1294),
    .X(booth_b56_m30));
 sky130_fd_sc_hd__a22o_1 \U$$3904  (.A1(net1028),
    .A2(net463),
    .B1(net1020),
    .B2(net736),
    .X(\t$6400 ));
 sky130_fd_sc_hd__xor2_1 \U$$3905  (.A(\t$6400 ),
    .B(net1292),
    .X(booth_b56_m31));
 sky130_fd_sc_hd__a22o_1 \U$$3906  (.A1(net1020),
    .A2(net462),
    .B1(net1003),
    .B2(net735),
    .X(\t$6401 ));
 sky130_fd_sc_hd__xor2_1 \U$$3907  (.A(\t$6401 ),
    .B(net1292),
    .X(booth_b56_m32));
 sky130_fd_sc_hd__a22o_1 \U$$3908  (.A1(net1003),
    .A2(net462),
    .B1(net995),
    .B2(net735),
    .X(\t$6402 ));
 sky130_fd_sc_hd__xor2_1 \U$$3909  (.A(\t$6402 ),
    .B(net1293),
    .X(booth_b56_m33));
 sky130_fd_sc_hd__xor2_1 \U$$391  (.A(\t$4604 ),
    .B(net1276),
    .X(booth_b4_m55));
 sky130_fd_sc_hd__a22o_1 \U$$3910  (.A1(net997),
    .A2(net465),
    .B1(net988),
    .B2(net738),
    .X(\t$6403 ));
 sky130_fd_sc_hd__xor2_1 \U$$3911  (.A(\t$6403 ),
    .B(net1297),
    .X(booth_b56_m34));
 sky130_fd_sc_hd__a22o_1 \U$$3912  (.A1(net988),
    .A2(net464),
    .B1(net979),
    .B2(net737),
    .X(\t$6404 ));
 sky130_fd_sc_hd__xor2_1 \U$$3913  (.A(\t$6404 ),
    .B(net1299),
    .X(booth_b56_m35));
 sky130_fd_sc_hd__a22o_1 \U$$3914  (.A1(net979),
    .A2(net465),
    .B1(net970),
    .B2(net738),
    .X(\t$6405 ));
 sky130_fd_sc_hd__xor2_1 \U$$3915  (.A(\t$6405 ),
    .B(net1297),
    .X(booth_b56_m36));
 sky130_fd_sc_hd__a22o_1 \U$$3916  (.A1(net970),
    .A2(net462),
    .B1(net962),
    .B2(net735),
    .X(\t$6406 ));
 sky130_fd_sc_hd__xor2_1 \U$$3917  (.A(\t$6406 ),
    .B(net1293),
    .X(booth_b56_m37));
 sky130_fd_sc_hd__a22o_1 \U$$3918  (.A1(net962),
    .A2(net464),
    .B1(net954),
    .B2(net737),
    .X(\t$6407 ));
 sky130_fd_sc_hd__xor2_1 \U$$3919  (.A(\t$6407 ),
    .B(net1296),
    .X(booth_b56_m38));
 sky130_fd_sc_hd__a22o_1 \U$$392  (.A1(net1614),
    .A2(net530),
    .B1(net1606),
    .B2(net803),
    .X(\t$4605 ));
 sky130_fd_sc_hd__a22o_1 \U$$3920  (.A1(net953),
    .A2(net464),
    .B1(net947),
    .B2(net737),
    .X(\t$6408 ));
 sky130_fd_sc_hd__xor2_1 \U$$3921  (.A(\t$6408 ),
    .B(net1299),
    .X(booth_b56_m39));
 sky130_fd_sc_hd__a22o_1 \U$$3922  (.A1(net945),
    .A2(net464),
    .B1(net929),
    .B2(net737),
    .X(\t$6409 ));
 sky130_fd_sc_hd__xor2_1 \U$$3923  (.A(\t$6409 ),
    .B(net1299),
    .X(booth_b56_m40));
 sky130_fd_sc_hd__a22o_1 \U$$3924  (.A1(net929),
    .A2(net465),
    .B1(net1750),
    .B2(net738),
    .X(\t$6410 ));
 sky130_fd_sc_hd__xor2_1 \U$$3925  (.A(\t$6410 ),
    .B(net1297),
    .X(booth_b56_m41));
 sky130_fd_sc_hd__a22o_1 \U$$3926  (.A1(net1750),
    .A2(net466),
    .B1(net1742),
    .B2(net739),
    .X(\t$6411 ));
 sky130_fd_sc_hd__xor2_1 \U$$3927  (.A(\t$6411 ),
    .B(net1298),
    .X(booth_b56_m42));
 sky130_fd_sc_hd__a22o_1 \U$$3928  (.A1(net1742),
    .A2(net466),
    .B1(net1734),
    .B2(net739),
    .X(\t$6412 ));
 sky130_fd_sc_hd__xor2_1 \U$$3929  (.A(\t$6412 ),
    .B(net1298),
    .X(booth_b56_m43));
 sky130_fd_sc_hd__xor2_1 \U$$393  (.A(\t$4605 ),
    .B(net1276),
    .X(booth_b4_m56));
 sky130_fd_sc_hd__a22o_1 \U$$3930  (.A1(net1734),
    .A2(net466),
    .B1(net1726),
    .B2(net739),
    .X(\t$6413 ));
 sky130_fd_sc_hd__xor2_1 \U$$3931  (.A(\t$6413 ),
    .B(net1298),
    .X(booth_b56_m44));
 sky130_fd_sc_hd__a22o_1 \U$$3932  (.A1(net1726),
    .A2(net466),
    .B1(net1718),
    .B2(net739),
    .X(\t$6414 ));
 sky130_fd_sc_hd__xor2_1 \U$$3933  (.A(\t$6414 ),
    .B(net1298),
    .X(booth_b56_m45));
 sky130_fd_sc_hd__a22o_1 \U$$3934  (.A1(net1718),
    .A2(net466),
    .B1(net1709),
    .B2(net739),
    .X(\t$6415 ));
 sky130_fd_sc_hd__xor2_1 \U$$3935  (.A(\t$6415 ),
    .B(net1298),
    .X(booth_b56_m46));
 sky130_fd_sc_hd__a22o_1 \U$$3936  (.A1(net1709),
    .A2(net466),
    .B1(net1701),
    .B2(net739),
    .X(\t$6416 ));
 sky130_fd_sc_hd__xor2_1 \U$$3937  (.A(\t$6416 ),
    .B(net1298),
    .X(booth_b56_m47));
 sky130_fd_sc_hd__a22o_1 \U$$3938  (.A1(net1701),
    .A2(net466),
    .B1(net1694),
    .B2(net739),
    .X(\t$6417 ));
 sky130_fd_sc_hd__xor2_1 \U$$3939  (.A(\t$6417 ),
    .B(net1298),
    .X(booth_b56_m48));
 sky130_fd_sc_hd__a22o_1 \U$$394  (.A1(net1604),
    .A2(net529),
    .B1(net1595),
    .B2(net802),
    .X(\t$4606 ));
 sky130_fd_sc_hd__a22o_1 \U$$3940  (.A1(net1693),
    .A2(net466),
    .B1(net1684),
    .B2(net739),
    .X(\t$6418 ));
 sky130_fd_sc_hd__xor2_1 \U$$3941  (.A(\t$6418 ),
    .B(net1298),
    .X(booth_b56_m49));
 sky130_fd_sc_hd__a22o_1 \U$$3942  (.A1(net1684),
    .A2(net465),
    .B1(net1660),
    .B2(net738),
    .X(\t$6419 ));
 sky130_fd_sc_hd__xor2_1 \U$$3943  (.A(\t$6419 ),
    .B(net1297),
    .X(booth_b56_m50));
 sky130_fd_sc_hd__a22o_1 \U$$3944  (.A1(net1659),
    .A2(net462),
    .B1(net1651),
    .B2(net735),
    .X(\t$6420 ));
 sky130_fd_sc_hd__xor2_1 \U$$3945  (.A(\t$6420 ),
    .B(net1293),
    .X(booth_b56_m51));
 sky130_fd_sc_hd__a22o_1 \U$$3946  (.A1(net1651),
    .A2(net462),
    .B1(net1643),
    .B2(net735),
    .X(\t$6421 ));
 sky130_fd_sc_hd__xor2_1 \U$$3947  (.A(\t$6421 ),
    .B(net1293),
    .X(booth_b56_m52));
 sky130_fd_sc_hd__a22o_1 \U$$3948  (.A1(net1643),
    .A2(net462),
    .B1(net1634),
    .B2(net735),
    .X(\t$6422 ));
 sky130_fd_sc_hd__xor2_1 \U$$3949  (.A(\t$6422 ),
    .B(net1293),
    .X(booth_b56_m53));
 sky130_fd_sc_hd__xor2_1 \U$$395  (.A(\t$4606 ),
    .B(net1275),
    .X(booth_b4_m57));
 sky130_fd_sc_hd__a22o_1 \U$$3950  (.A1(net1634),
    .A2(net465),
    .B1(net1624),
    .B2(net738),
    .X(\t$6423 ));
 sky130_fd_sc_hd__xor2_1 \U$$3951  (.A(\t$6423 ),
    .B(net1297),
    .X(booth_b56_m54));
 sky130_fd_sc_hd__a22o_1 \U$$3952  (.A1(net1624),
    .A2(net465),
    .B1(net1616),
    .B2(net738),
    .X(\t$6424 ));
 sky130_fd_sc_hd__xor2_1 \U$$3953  (.A(\t$6424 ),
    .B(net1297),
    .X(booth_b56_m55));
 sky130_fd_sc_hd__a22o_1 \U$$3954  (.A1(net1616),
    .A2(net465),
    .B1(net1608),
    .B2(net738),
    .X(\t$6425 ));
 sky130_fd_sc_hd__xor2_1 \U$$3955  (.A(\t$6425 ),
    .B(net1297),
    .X(booth_b56_m56));
 sky130_fd_sc_hd__a22o_1 \U$$3956  (.A1(net1608),
    .A2(net465),
    .B1(net1600),
    .B2(net738),
    .X(\t$6426 ));
 sky130_fd_sc_hd__xor2_1 \U$$3957  (.A(\t$6426 ),
    .B(net1297),
    .X(booth_b56_m57));
 sky130_fd_sc_hd__a22o_1 \U$$3958  (.A1(net1601),
    .A2(net465),
    .B1(net1591),
    .B2(net738),
    .X(\t$6427 ));
 sky130_fd_sc_hd__xor2_1 \U$$3959  (.A(\t$6427 ),
    .B(net1297),
    .X(booth_b56_m58));
 sky130_fd_sc_hd__a22o_1 \U$$396  (.A1(net1595),
    .A2(net529),
    .B1(net1586),
    .B2(net802),
    .X(\t$4607 ));
 sky130_fd_sc_hd__a22o_1 \U$$3960  (.A1(net1591),
    .A2(net462),
    .B1(net1583),
    .B2(net735),
    .X(\t$6428 ));
 sky130_fd_sc_hd__xor2_1 \U$$3961  (.A(\t$6428 ),
    .B(net1292),
    .X(booth_b56_m59));
 sky130_fd_sc_hd__a22o_1 \U$$3962  (.A1(net1584),
    .A2(net465),
    .B1(net1557),
    .B2(net738),
    .X(\t$6429 ));
 sky130_fd_sc_hd__xor2_1 \U$$3963  (.A(\t$6429 ),
    .B(net1297),
    .X(booth_b56_m60));
 sky130_fd_sc_hd__a22o_1 \U$$3964  (.A1(net1554),
    .A2(net463),
    .B1(net1545),
    .B2(net736),
    .X(\t$6430 ));
 sky130_fd_sc_hd__xor2_1 \U$$3965  (.A(\t$6430 ),
    .B(net1292),
    .X(booth_b56_m61));
 sky130_fd_sc_hd__a22o_1 \U$$3966  (.A1(net1549),
    .A2(net462),
    .B1(net1541),
    .B2(net735),
    .X(\t$6431 ));
 sky130_fd_sc_hd__xor2_1 \U$$3967  (.A(\t$6431 ),
    .B(net1293),
    .X(booth_b56_m62));
 sky130_fd_sc_hd__a22o_1 \U$$3968  (.A1(net1541),
    .A2(net463),
    .B1(net1533),
    .B2(net736),
    .X(\t$6432 ));
 sky130_fd_sc_hd__xor2_1 \U$$3969  (.A(\t$6432 ),
    .B(net1293),
    .X(booth_b56_m63));
 sky130_fd_sc_hd__xor2_1 \U$$397  (.A(\t$4607 ),
    .B(net1275),
    .X(booth_b4_m58));
 sky130_fd_sc_hd__a22o_1 \U$$3970  (.A1(net1529),
    .A2(net462),
    .B1(net1800),
    .B2(net735),
    .X(\t$6433 ));
 sky130_fd_sc_hd__xor2_1 \U$$3971  (.A(\t$6433 ),
    .B(net1293),
    .X(booth_b56_m64));
 sky130_fd_sc_hd__inv_1 \U$$3972  (.A(net1293),
    .Y(\notsign$6434 ));
 sky130_fd_sc_hd__inv_1 \U$$3973  (.A(net1292),
    .Y(\notblock$6435[0] ));
 sky130_fd_sc_hd__inv_1 \U$$3974  (.A(net54),
    .Y(\notblock$6435[1] ));
 sky130_fd_sc_hd__inv_1 \U$$3975  (.A(net1284),
    .Y(\notblock$6435[2] ));
 sky130_fd_sc_hd__and2_1 \U$$3976  (.A(net1284),
    .B(\notblock$6435[1] ),
    .X(\t$6436 ));
 sky130_fd_sc_hd__a32o_1 \U$$3977  (.A1(\notblock$6435[2] ),
    .A2(net54),
    .A3(net1292),
    .B1(\t$6436 ),
    .B2(\notblock$6435[0] ),
    .X(\sel_0$6437 ));
 sky130_fd_sc_hd__xor2_1 \U$$3978  (.A(net54),
    .B(net1292),
    .X(\sel_1$6438 ));
 sky130_fd_sc_hd__a22o_1 \U$$3979  (.A1(net1801),
    .A2(net455),
    .B1(net1233),
    .B2(net728),
    .X(\t$6439 ));
 sky130_fd_sc_hd__a22o_1 \U$$398  (.A1(net1586),
    .A2(net529),
    .B1(net1578),
    .B2(net802),
    .X(\t$4608 ));
 sky130_fd_sc_hd__xor2_1 \U$$3980  (.A(\t$6439 ),
    .B(net1287),
    .X(booth_b58_m0));
 sky130_fd_sc_hd__a22o_1 \U$$3981  (.A1(net1233),
    .A2(net451),
    .B1(net1129),
    .B2(net724),
    .X(\t$6440 ));
 sky130_fd_sc_hd__xor2_1 \U$$3982  (.A(\t$6440 ),
    .B(net1282),
    .X(booth_b58_m1));
 sky130_fd_sc_hd__a22o_1 \U$$3983  (.A1(net1125),
    .A2(net451),
    .B1(net1034),
    .B2(net724),
    .X(\t$6441 ));
 sky130_fd_sc_hd__xor2_1 \U$$3984  (.A(\t$6441 ),
    .B(net1282),
    .X(booth_b58_m2));
 sky130_fd_sc_hd__a22o_1 \U$$3985  (.A1(net1034),
    .A2(net451),
    .B1(net935),
    .B2(net724),
    .X(\t$6442 ));
 sky130_fd_sc_hd__xor2_1 \U$$3986  (.A(\t$6442 ),
    .B(net1282),
    .X(booth_b58_m3));
 sky130_fd_sc_hd__a22o_1 \U$$3987  (.A1(net935),
    .A2(net452),
    .B1(net1674),
    .B2(net725),
    .X(\t$6443 ));
 sky130_fd_sc_hd__xor2_1 \U$$3988  (.A(\t$6443 ),
    .B(net1283),
    .X(booth_b58_m4));
 sky130_fd_sc_hd__a22o_1 \U$$3989  (.A1(net1674),
    .A2(net451),
    .B1(net1563),
    .B2(net724),
    .X(\t$6444 ));
 sky130_fd_sc_hd__xor2_1 \U$$399  (.A(\t$4608 ),
    .B(net1275),
    .X(booth_b4_m59));
 sky130_fd_sc_hd__xor2_1 \U$$3990  (.A(\t$6444 ),
    .B(net1282),
    .X(booth_b58_m5));
 sky130_fd_sc_hd__a22o_1 \U$$3991  (.A1(net1566),
    .A2(net458),
    .B1(net1525),
    .B2(net731),
    .X(\t$6445 ));
 sky130_fd_sc_hd__xor2_1 \U$$3992  (.A(\t$6445 ),
    .B(net1287),
    .X(booth_b58_m6));
 sky130_fd_sc_hd__a22o_1 \U$$3993  (.A1(net1525),
    .A2(net455),
    .B1(net1517),
    .B2(net728),
    .X(\t$6446 ));
 sky130_fd_sc_hd__xor2_1 \U$$3994  (.A(\t$6446 ),
    .B(net1287),
    .X(booth_b58_m7));
 sky130_fd_sc_hd__a22o_1 \U$$3995  (.A1(net1517),
    .A2(net455),
    .B1(net1510),
    .B2(net728),
    .X(\t$6447 ));
 sky130_fd_sc_hd__xor2_1 \U$$3996  (.A(\t$6447 ),
    .B(net1287),
    .X(booth_b58_m8));
 sky130_fd_sc_hd__a22o_1 \U$$3997  (.A1(net1510),
    .A2(net455),
    .B1(net1501),
    .B2(net728),
    .X(\t$6448 ));
 sky130_fd_sc_hd__xor2_1 \U$$3998  (.A(\t$6448 ),
    .B(net1287),
    .X(booth_b58_m9));
 sky130_fd_sc_hd__a22o_1 \U$$3999  (.A1(net1502),
    .A2(net455),
    .B1(net66),
    .B2(net728),
    .X(\t$6449 ));
 sky130_fd_sc_hd__a32o_1 \U$$4  (.A1(\notblock[2] ),
    .A2(net1),
    .A3(net1802),
    .B1(t),
    .B2(\notblock[0] ),
    .X(sel_0));
 sky130_fd_sc_hd__a22o_1 \U$$40  (.A1(net1157),
    .A2(net443),
    .B1(net1147),
    .B2(net685),
    .X(\t$4427 ));
 sky130_fd_sc_hd__a22o_1 \U$$400  (.A1(net1578),
    .A2(net529),
    .B1(net1551),
    .B2(net802),
    .X(\t$4609 ));
 sky130_fd_sc_hd__xor2_1 \U$$4000  (.A(\t$6449 ),
    .B(net1287),
    .X(booth_b58_m10));
 sky130_fd_sc_hd__a22o_1 \U$$4001  (.A1(net66),
    .A2(net458),
    .B1(net1218),
    .B2(net731),
    .X(\t$6450 ));
 sky130_fd_sc_hd__xor2_1 \U$$4002  (.A(\t$6450 ),
    .B(net1287),
    .X(booth_b58_m11));
 sky130_fd_sc_hd__a22o_1 \U$$4003  (.A1(net1215),
    .A2(net452),
    .B1(net1205),
    .B2(net725),
    .X(\t$6451 ));
 sky130_fd_sc_hd__xor2_1 \U$$4004  (.A(\t$6451 ),
    .B(net1283),
    .X(booth_b58_m12));
 sky130_fd_sc_hd__a22o_1 \U$$4005  (.A1(net1205),
    .A2(net452),
    .B1(net1197),
    .B2(net725),
    .X(\t$6452 ));
 sky130_fd_sc_hd__xor2_1 \U$$4006  (.A(\t$6452 ),
    .B(net1283),
    .X(booth_b58_m13));
 sky130_fd_sc_hd__a22o_1 \U$$4007  (.A1(net1196),
    .A2(net451),
    .B1(net1177),
    .B2(net724),
    .X(\t$6453 ));
 sky130_fd_sc_hd__xor2_1 \U$$4008  (.A(\t$6453 ),
    .B(net1282),
    .X(booth_b58_m14));
 sky130_fd_sc_hd__a22o_1 \U$$4009  (.A1(net1177),
    .A2(net451),
    .B1(net1168),
    .B2(net724),
    .X(\t$6454 ));
 sky130_fd_sc_hd__xor2_1 \U$$401  (.A(\t$4609 ),
    .B(net1275),
    .X(booth_b4_m60));
 sky130_fd_sc_hd__xor2_1 \U$$4010  (.A(\t$6454 ),
    .B(net1282),
    .X(booth_b58_m15));
 sky130_fd_sc_hd__a22o_1 \U$$4011  (.A1(net1168),
    .A2(net451),
    .B1(net1159),
    .B2(net724),
    .X(\t$6455 ));
 sky130_fd_sc_hd__xor2_1 \U$$4012  (.A(\t$6455 ),
    .B(net1282),
    .X(booth_b58_m16));
 sky130_fd_sc_hd__a22o_1 \U$$4013  (.A1(net1159),
    .A2(net451),
    .B1(net1152),
    .B2(net724),
    .X(\t$6456 ));
 sky130_fd_sc_hd__xor2_1 \U$$4014  (.A(\t$6456 ),
    .B(net1282),
    .X(booth_b58_m17));
 sky130_fd_sc_hd__a22o_1 \U$$4015  (.A1(net1152),
    .A2(net451),
    .B1(net1141),
    .B2(net724),
    .X(\t$6457 ));
 sky130_fd_sc_hd__xor2_1 \U$$4016  (.A(\t$6457 ),
    .B(net1282),
    .X(booth_b58_m18));
 sky130_fd_sc_hd__a22o_1 \U$$4017  (.A1(net1142),
    .A2(net452),
    .B1(net1135),
    .B2(net725),
    .X(\t$6458 ));
 sky130_fd_sc_hd__xor2_1 \U$$4018  (.A(\t$6458 ),
    .B(net1283),
    .X(booth_b58_m19));
 sky130_fd_sc_hd__a22o_1 \U$$4019  (.A1(net1135),
    .A2(net451),
    .B1(net1119),
    .B2(net724),
    .X(\t$6459 ));
 sky130_fd_sc_hd__a22o_1 \U$$402  (.A1(net1555),
    .A2(net533),
    .B1(net1547),
    .B2(net806),
    .X(\t$4610 ));
 sky130_fd_sc_hd__xor2_1 \U$$4020  (.A(\t$6459 ),
    .B(net1282),
    .X(booth_b58_m20));
 sky130_fd_sc_hd__a22o_1 \U$$4021  (.A1(net1119),
    .A2(net454),
    .B1(net1112),
    .B2(net727),
    .X(\t$6460 ));
 sky130_fd_sc_hd__xor2_1 \U$$4022  (.A(\t$6460 ),
    .B(net1286),
    .X(booth_b58_m21));
 sky130_fd_sc_hd__a22o_1 \U$$4023  (.A1(net1112),
    .A2(net453),
    .B1(net1103),
    .B2(net726),
    .X(\t$6461 ));
 sky130_fd_sc_hd__xor2_1 \U$$4024  (.A(\t$6461 ),
    .B(net1285),
    .X(booth_b58_m22));
 sky130_fd_sc_hd__a22o_1 \U$$4025  (.A1(net1103),
    .A2(net454),
    .B1(net1094),
    .B2(net727),
    .X(\t$6462 ));
 sky130_fd_sc_hd__xor2_1 \U$$4026  (.A(\t$6462 ),
    .B(net1286),
    .X(booth_b58_m23));
 sky130_fd_sc_hd__a22o_1 \U$$4027  (.A1(net1095),
    .A2(net454),
    .B1(net1085),
    .B2(net727),
    .X(\t$6463 ));
 sky130_fd_sc_hd__xor2_1 \U$$4028  (.A(\t$6463 ),
    .B(net1286),
    .X(booth_b58_m24));
 sky130_fd_sc_hd__a22o_1 \U$$4029  (.A1(net1085),
    .A2(net454),
    .B1(net1077),
    .B2(net727),
    .X(\t$6464 ));
 sky130_fd_sc_hd__xor2_1 \U$$403  (.A(\t$4610 ),
    .B(net1280),
    .X(booth_b4_m61));
 sky130_fd_sc_hd__xor2_1 \U$$4030  (.A(\t$6464 ),
    .B(net1286),
    .X(booth_b58_m25));
 sky130_fd_sc_hd__a22o_1 \U$$4031  (.A1(net1077),
    .A2(net454),
    .B1(net1069),
    .B2(net727),
    .X(\t$6465 ));
 sky130_fd_sc_hd__xor2_1 \U$$4032  (.A(\t$6465 ),
    .B(net1286),
    .X(booth_b58_m26));
 sky130_fd_sc_hd__a22o_1 \U$$4033  (.A1(net1069),
    .A2(net454),
    .B1(net1061),
    .B2(net727),
    .X(\t$6466 ));
 sky130_fd_sc_hd__xor2_1 \U$$4034  (.A(\t$6466 ),
    .B(net1286),
    .X(booth_b58_m27));
 sky130_fd_sc_hd__a22o_1 \U$$4035  (.A1(net1061),
    .A2(net454),
    .B1(net1052),
    .B2(net727),
    .X(\t$6467 ));
 sky130_fd_sc_hd__xor2_1 \U$$4036  (.A(\t$6467 ),
    .B(net1286),
    .X(booth_b58_m28));
 sky130_fd_sc_hd__a22o_1 \U$$4037  (.A1(net1052),
    .A2(net454),
    .B1(net1044),
    .B2(net727),
    .X(\t$6468 ));
 sky130_fd_sc_hd__xor2_1 \U$$4038  (.A(\t$6468 ),
    .B(net1286),
    .X(booth_b58_m29));
 sky130_fd_sc_hd__a22o_1 \U$$4039  (.A1(net1045),
    .A2(net453),
    .B1(net1028),
    .B2(net726),
    .X(\t$6469 ));
 sky130_fd_sc_hd__a22o_1 \U$$404  (.A1(net1547),
    .A2(net533),
    .B1(net1539),
    .B2(net806),
    .X(\t$4611 ));
 sky130_fd_sc_hd__xor2_1 \U$$4040  (.A(\t$6469 ),
    .B(net1284),
    .X(booth_b58_m30));
 sky130_fd_sc_hd__a22o_1 \U$$4041  (.A1(net1028),
    .A2(net453),
    .B1(net1020),
    .B2(net726),
    .X(\t$6470 ));
 sky130_fd_sc_hd__xor2_1 \U$$4042  (.A(\t$6470 ),
    .B(net1285),
    .X(booth_b58_m31));
 sky130_fd_sc_hd__a22o_1 \U$$4043  (.A1(net1021),
    .A2(net456),
    .B1(net1004),
    .B2(net729),
    .X(\t$6471 ));
 sky130_fd_sc_hd__xor2_1 \U$$4044  (.A(\t$6471 ),
    .B(net1288),
    .X(booth_b58_m32));
 sky130_fd_sc_hd__a22o_1 \U$$4045  (.A1(net1004),
    .A2(net455),
    .B1(net996),
    .B2(net728),
    .X(\t$6472 ));
 sky130_fd_sc_hd__xor2_1 \U$$4046  (.A(\t$6472 ),
    .B(net1287),
    .X(booth_b58_m33));
 sky130_fd_sc_hd__a22o_1 \U$$4047  (.A1(net996),
    .A2(net455),
    .B1(net988),
    .B2(net728),
    .X(\t$6473 ));
 sky130_fd_sc_hd__xor2_1 \U$$4048  (.A(\t$6473 ),
    .B(net1289),
    .X(booth_b58_m34));
 sky130_fd_sc_hd__a22o_1 \U$$4049  (.A1(net988),
    .A2(net452),
    .B1(net979),
    .B2(net725),
    .X(\t$6474 ));
 sky130_fd_sc_hd__xor2_1 \U$$405  (.A(\t$4611 ),
    .B(net1280),
    .X(booth_b4_m62));
 sky130_fd_sc_hd__xor2_1 \U$$4050  (.A(\t$6474 ),
    .B(net1283),
    .X(booth_b58_m35));
 sky130_fd_sc_hd__a22o_1 \U$$4051  (.A1(net979),
    .A2(net455),
    .B1(net970),
    .B2(net728),
    .X(\t$6475 ));
 sky130_fd_sc_hd__xor2_1 \U$$4052  (.A(\t$6475 ),
    .B(net1287),
    .X(booth_b58_m36));
 sky130_fd_sc_hd__a22o_1 \U$$4053  (.A1(net970),
    .A2(net455),
    .B1(net962),
    .B2(net728),
    .X(\t$6476 ));
 sky130_fd_sc_hd__xor2_1 \U$$4054  (.A(\t$6476 ),
    .B(net1290),
    .X(booth_b58_m37));
 sky130_fd_sc_hd__a22o_1 \U$$4055  (.A1(net962),
    .A2(net455),
    .B1(net953),
    .B2(net728),
    .X(\t$6477 ));
 sky130_fd_sc_hd__xor2_1 \U$$4056  (.A(\t$6477 ),
    .B(net1290),
    .X(booth_b58_m38));
 sky130_fd_sc_hd__a22o_1 \U$$4057  (.A1(net953),
    .A2(net457),
    .B1(net945),
    .B2(net730),
    .X(\t$6478 ));
 sky130_fd_sc_hd__xor2_1 \U$$4058  (.A(\t$6478 ),
    .B(net1289),
    .X(booth_b58_m39));
 sky130_fd_sc_hd__a22o_1 \U$$4059  (.A1(net945),
    .A2(net457),
    .B1(net929),
    .B2(net730),
    .X(\t$6479 ));
 sky130_fd_sc_hd__a22o_1 \U$$406  (.A1(net1539),
    .A2(net534),
    .B1(net1531),
    .B2(net807),
    .X(\t$4612 ));
 sky130_fd_sc_hd__xor2_1 \U$$4060  (.A(\t$6479 ),
    .B(net1289),
    .X(booth_b58_m40));
 sky130_fd_sc_hd__a22o_1 \U$$4061  (.A1(net929),
    .A2(net457),
    .B1(net1750),
    .B2(net730),
    .X(\t$6480 ));
 sky130_fd_sc_hd__xor2_1 \U$$4062  (.A(\t$6480 ),
    .B(net1289),
    .X(booth_b58_m41));
 sky130_fd_sc_hd__a22o_1 \U$$4063  (.A1(net1750),
    .A2(net457),
    .B1(net1742),
    .B2(net730),
    .X(\t$6481 ));
 sky130_fd_sc_hd__xor2_1 \U$$4064  (.A(\t$6481 ),
    .B(net1289),
    .X(booth_b58_m42));
 sky130_fd_sc_hd__a22o_1 \U$$4065  (.A1(net1742),
    .A2(net457),
    .B1(net1734),
    .B2(net730),
    .X(\t$6482 ));
 sky130_fd_sc_hd__xor2_1 \U$$4066  (.A(\t$6482 ),
    .B(net1289),
    .X(booth_b58_m43));
 sky130_fd_sc_hd__a22o_1 \U$$4067  (.A1(net1736),
    .A2(net457),
    .B1(net1728),
    .B2(net730),
    .X(\t$6483 ));
 sky130_fd_sc_hd__xor2_1 \U$$4068  (.A(\t$6483 ),
    .B(net1289),
    .X(booth_b58_m44));
 sky130_fd_sc_hd__a22o_1 \U$$4069  (.A1(net1728),
    .A2(net457),
    .B1(net1718),
    .B2(net730),
    .X(\t$6484 ));
 sky130_fd_sc_hd__xor2_1 \U$$407  (.A(\t$4612 ),
    .B(net1281),
    .X(booth_b4_m63));
 sky130_fd_sc_hd__xor2_1 \U$$4070  (.A(\t$6484 ),
    .B(net1289),
    .X(booth_b58_m45));
 sky130_fd_sc_hd__a22o_1 \U$$4071  (.A1(net1718),
    .A2(net457),
    .B1(net1709),
    .B2(net730),
    .X(\t$6485 ));
 sky130_fd_sc_hd__xor2_1 \U$$4072  (.A(\t$6485 ),
    .B(net1289),
    .X(booth_b58_m46));
 sky130_fd_sc_hd__a22o_1 \U$$4073  (.A1(net1708),
    .A2(net456),
    .B1(net1700),
    .B2(net729),
    .X(\t$6486 ));
 sky130_fd_sc_hd__xor2_1 \U$$4074  (.A(\t$6486 ),
    .B(net1289),
    .X(booth_b58_m47));
 sky130_fd_sc_hd__a22o_1 \U$$4075  (.A1(net1700),
    .A2(net456),
    .B1(net1693),
    .B2(net729),
    .X(\t$6487 ));
 sky130_fd_sc_hd__xor2_1 \U$$4076  (.A(\t$6487 ),
    .B(net1288),
    .X(booth_b58_m48));
 sky130_fd_sc_hd__a22o_1 \U$$4077  (.A1(net1692),
    .A2(net453),
    .B1(net1685),
    .B2(net726),
    .X(\t$6488 ));
 sky130_fd_sc_hd__xor2_1 \U$$4078  (.A(\t$6488 ),
    .B(net1285),
    .X(booth_b58_m49));
 sky130_fd_sc_hd__a22o_1 \U$$4079  (.A1(net1685),
    .A2(net453),
    .B1(net1659),
    .B2(net726),
    .X(\t$6489 ));
 sky130_fd_sc_hd__a22o_1 \U$$408  (.A1(net1531),
    .A2(net533),
    .B1(net1803),
    .B2(net806),
    .X(\t$4613 ));
 sky130_fd_sc_hd__xor2_1 \U$$4080  (.A(\t$6489 ),
    .B(net1285),
    .X(booth_b58_m50));
 sky130_fd_sc_hd__a22o_1 \U$$4081  (.A1(net1659),
    .A2(net453),
    .B1(net1651),
    .B2(net726),
    .X(\t$6490 ));
 sky130_fd_sc_hd__xor2_1 \U$$4082  (.A(\t$6490 ),
    .B(net1285),
    .X(booth_b58_m51));
 sky130_fd_sc_hd__a22o_1 \U$$4083  (.A1(net1651),
    .A2(net456),
    .B1(net1643),
    .B2(net729),
    .X(\t$6491 ));
 sky130_fd_sc_hd__xor2_1 \U$$4084  (.A(\t$6491 ),
    .B(net1288),
    .X(booth_b58_m52));
 sky130_fd_sc_hd__a22o_1 \U$$4085  (.A1(net1643),
    .A2(net456),
    .B1(net1634),
    .B2(net729),
    .X(\t$6492 ));
 sky130_fd_sc_hd__xor2_1 \U$$4086  (.A(\t$6492 ),
    .B(net1288),
    .X(booth_b58_m53));
 sky130_fd_sc_hd__a22o_1 \U$$4087  (.A1(net1634),
    .A2(net456),
    .B1(net1624),
    .B2(net729),
    .X(\t$6493 ));
 sky130_fd_sc_hd__xor2_1 \U$$4088  (.A(\t$6493 ),
    .B(net1288),
    .X(booth_b58_m54));
 sky130_fd_sc_hd__a22o_1 \U$$4089  (.A1(net1625),
    .A2(net456),
    .B1(net1616),
    .B2(net729),
    .X(\t$6494 ));
 sky130_fd_sc_hd__xor2_1 \U$$409  (.A(\t$4613 ),
    .B(net1280),
    .X(booth_b4_m64));
 sky130_fd_sc_hd__xor2_1 \U$$4090  (.A(\t$6494 ),
    .B(net1288),
    .X(booth_b58_m55));
 sky130_fd_sc_hd__a22o_1 \U$$4091  (.A1(net1617),
    .A2(net456),
    .B1(net1610),
    .B2(net729),
    .X(\t$6495 ));
 sky130_fd_sc_hd__xor2_1 \U$$4092  (.A(\t$6495 ),
    .B(net1288),
    .X(booth_b58_m56));
 sky130_fd_sc_hd__a22o_1 \U$$4093  (.A1(net1610),
    .A2(net456),
    .B1(net1601),
    .B2(net729),
    .X(\t$6496 ));
 sky130_fd_sc_hd__xor2_1 \U$$4094  (.A(\t$6496 ),
    .B(net1288),
    .X(booth_b58_m57));
 sky130_fd_sc_hd__a22o_1 \U$$4095  (.A1(net1601),
    .A2(net456),
    .B1(net1592),
    .B2(net729),
    .X(\t$6497 ));
 sky130_fd_sc_hd__xor2_1 \U$$4096  (.A(\t$6497 ),
    .B(net1288),
    .X(booth_b58_m58));
 sky130_fd_sc_hd__a22o_1 \U$$4097  (.A1(net1589),
    .A2(net453),
    .B1(net1580),
    .B2(net726),
    .X(\t$6498 ));
 sky130_fd_sc_hd__xor2_1 \U$$4098  (.A(\t$6498 ),
    .B(net1284),
    .X(booth_b58_m59));
 sky130_fd_sc_hd__a22o_1 \U$$4099  (.A1(net1584),
    .A2(net459),
    .B1(net1557),
    .B2(net732),
    .X(\t$6499 ));
 sky130_fd_sc_hd__xor2_1 \U$$41  (.A(\t$4427 ),
    .B(net1569),
    .X(booth_b0_m17));
 sky130_fd_sc_hd__inv_1 \U$$410  (.A(net1280),
    .Y(\notsign$4614 ));
 sky130_fd_sc_hd__xor2_1 \U$$4100  (.A(\t$6499 ),
    .B(net1284),
    .X(booth_b58_m60));
 sky130_fd_sc_hd__a22o_1 \U$$4101  (.A1(net1557),
    .A2(net453),
    .B1(net1549),
    .B2(net726),
    .X(\t$6500 ));
 sky130_fd_sc_hd__xor2_1 \U$$4102  (.A(\t$6500 ),
    .B(net1288),
    .X(booth_b58_m61));
 sky130_fd_sc_hd__a22o_1 \U$$4103  (.A1(net1548),
    .A2(net453),
    .B1(net1540),
    .B2(net726),
    .X(\t$6501 ));
 sky130_fd_sc_hd__xor2_1 \U$$4104  (.A(\t$6501 ),
    .B(net1285),
    .X(booth_b58_m62));
 sky130_fd_sc_hd__a22o_1 \U$$4105  (.A1(net1541),
    .A2(net454),
    .B1(net1533),
    .B2(net727),
    .X(\t$6502 ));
 sky130_fd_sc_hd__xor2_1 \U$$4106  (.A(\t$6502 ),
    .B(net1285),
    .X(booth_b58_m63));
 sky130_fd_sc_hd__a22o_1 \U$$4107  (.A1(net1529),
    .A2(net453),
    .B1(net1804),
    .B2(net726),
    .X(\t$6503 ));
 sky130_fd_sc_hd__xor2_1 \U$$4108  (.A(\t$6503 ),
    .B(net1284),
    .X(booth_b58_m64));
 sky130_fd_sc_hd__inv_1 \U$$4109  (.A(net1284),
    .Y(\notsign$6504 ));
 sky130_fd_sc_hd__inv_1 \U$$411  (.A(net1275),
    .Y(\notblock$4615[0] ));
 sky130_fd_sc_hd__inv_1 \U$$4110  (.A(net1284),
    .Y(\notblock$6505[0] ));
 sky130_fd_sc_hd__inv_1 \U$$4111  (.A(net57),
    .Y(\notblock$6505[1] ));
 sky130_fd_sc_hd__inv_1 \U$$4112  (.A(net1265),
    .Y(\notblock$6505[2] ));
 sky130_fd_sc_hd__and2_1 \U$$4113  (.A(net1265),
    .B(\notblock$6505[1] ),
    .X(\t$6506 ));
 sky130_fd_sc_hd__a32o_1 \U$$4114  (.A1(\notblock$6505[2] ),
    .A2(net57),
    .A3(net1284),
    .B1(\t$6506 ),
    .B2(\notblock$6505[0] ),
    .X(\sel_0$6507 ));
 sky130_fd_sc_hd__xor2_1 \U$$4115  (.A(net57),
    .B(net1284),
    .X(\sel_1$6508 ));
 sky130_fd_sc_hd__a22o_1 \U$$4116  (.A1(net1805),
    .A2(net434),
    .B1(net1229),
    .B2(net716),
    .X(\t$6509 ));
 sky130_fd_sc_hd__xor2_1 \U$$4117  (.A(\t$6509 ),
    .B(net1263),
    .X(booth_b60_m0));
 sky130_fd_sc_hd__a22o_1 \U$$4118  (.A1(net1229),
    .A2(net434),
    .B1(net1125),
    .B2(net716),
    .X(\t$6510 ));
 sky130_fd_sc_hd__xor2_1 \U$$4119  (.A(\t$6510 ),
    .B(net1263),
    .X(booth_b60_m1));
 sky130_fd_sc_hd__inv_1 \U$$412  (.A(net61),
    .Y(\notblock$4615[1] ));
 sky130_fd_sc_hd__a22o_1 \U$$4120  (.A1(net1125),
    .A2(net437),
    .B1(net1034),
    .B2(net719),
    .X(\t$6511 ));
 sky130_fd_sc_hd__xor2_1 \U$$4121  (.A(\t$6511 ),
    .B(net1264),
    .X(booth_b60_m2));
 sky130_fd_sc_hd__a22o_1 \U$$4122  (.A1(net87),
    .A2(net434),
    .B1(net98),
    .B2(net716),
    .X(\t$6512 ));
 sky130_fd_sc_hd__xor2_1 \U$$4123  (.A(\t$6512 ),
    .B(net1264),
    .X(booth_b60_m3));
 sky130_fd_sc_hd__a22o_1 \U$$4124  (.A1(net938),
    .A2(net438),
    .B1(net1677),
    .B2(net720),
    .X(\t$6513 ));
 sky130_fd_sc_hd__xor2_1 \U$$4125  (.A(\t$6513 ),
    .B(net1269),
    .X(booth_b60_m4));
 sky130_fd_sc_hd__a22o_1 \U$$4126  (.A1(net1677),
    .A2(net438),
    .B1(net1566),
    .B2(net720),
    .X(\t$6514 ));
 sky130_fd_sc_hd__xor2_1 \U$$4127  (.A(\t$6514 ),
    .B(net1269),
    .X(booth_b60_m5));
 sky130_fd_sc_hd__a22o_1 \U$$4128  (.A1(net1567),
    .A2(net438),
    .B1(net1525),
    .B2(net720),
    .X(\t$6515 ));
 sky130_fd_sc_hd__xor2_1 \U$$4129  (.A(\t$6515 ),
    .B(net1269),
    .X(booth_b60_m6));
 sky130_fd_sc_hd__inv_1 \U$$413  (.A(net1246),
    .Y(\notblock$4615[2] ));
 sky130_fd_sc_hd__a22o_1 \U$$4130  (.A1(net1525),
    .A2(net438),
    .B1(net1517),
    .B2(net720),
    .X(\t$6516 ));
 sky130_fd_sc_hd__xor2_1 \U$$4131  (.A(\t$6516 ),
    .B(net1269),
    .X(booth_b60_m7));
 sky130_fd_sc_hd__a22o_1 \U$$4132  (.A1(net1517),
    .A2(net438),
    .B1(net127),
    .B2(net720),
    .X(\t$6517 ));
 sky130_fd_sc_hd__xor2_1 \U$$4133  (.A(\t$6517 ),
    .B(net1269),
    .X(booth_b60_m8));
 sky130_fd_sc_hd__a22o_1 \U$$4134  (.A1(net127),
    .A2(net438),
    .B1(net1502),
    .B2(net720),
    .X(\t$6518 ));
 sky130_fd_sc_hd__xor2_1 \U$$4135  (.A(\t$6518 ),
    .B(net1269),
    .X(booth_b60_m9));
 sky130_fd_sc_hd__a22o_1 \U$$4136  (.A1(net1498),
    .A2(net437),
    .B1(net1223),
    .B2(net719),
    .X(\t$6519 ));
 sky130_fd_sc_hd__xor2_1 \U$$4137  (.A(\t$6519 ),
    .B(net1264),
    .X(booth_b60_m10));
 sky130_fd_sc_hd__a22o_1 \U$$4138  (.A1(net1223),
    .A2(net434),
    .B1(net1215),
    .B2(net716),
    .X(\t$6520 ));
 sky130_fd_sc_hd__xor2_1 \U$$4139  (.A(\t$6520 ),
    .B(net1264),
    .X(booth_b60_m11));
 sky130_fd_sc_hd__and2_1 \U$$414  (.A(net1246),
    .B(\notblock$4615[1] ),
    .X(\t$4616 ));
 sky130_fd_sc_hd__a22o_1 \U$$4140  (.A1(net1214),
    .A2(net434),
    .B1(net1205),
    .B2(net716),
    .X(\t$6521 ));
 sky130_fd_sc_hd__xor2_1 \U$$4141  (.A(\t$6521 ),
    .B(net1263),
    .X(booth_b60_m12));
 sky130_fd_sc_hd__a22o_1 \U$$4142  (.A1(net1205),
    .A2(net434),
    .B1(net1196),
    .B2(net716),
    .X(\t$6522 ));
 sky130_fd_sc_hd__xor2_1 \U$$4143  (.A(\t$6522 ),
    .B(net1263),
    .X(booth_b60_m13));
 sky130_fd_sc_hd__a22o_1 \U$$4144  (.A1(net1196),
    .A2(net434),
    .B1(net1177),
    .B2(net716),
    .X(\t$6523 ));
 sky130_fd_sc_hd__xor2_1 \U$$4145  (.A(\t$6523 ),
    .B(net1263),
    .X(booth_b60_m14));
 sky130_fd_sc_hd__a22o_1 \U$$4146  (.A1(net1177),
    .A2(net434),
    .B1(net1168),
    .B2(net716),
    .X(\t$6524 ));
 sky130_fd_sc_hd__xor2_1 \U$$4147  (.A(\t$6524 ),
    .B(net1263),
    .X(booth_b60_m15));
 sky130_fd_sc_hd__a22o_1 \U$$4148  (.A1(net1168),
    .A2(net434),
    .B1(net1159),
    .B2(net716),
    .X(\t$6525 ));
 sky130_fd_sc_hd__xor2_1 \U$$4149  (.A(\t$6525 ),
    .B(net1263),
    .X(booth_b60_m16));
 sky130_fd_sc_hd__a32o_1 \U$$415  (.A1(\notblock$4615[2] ),
    .A2(net61),
    .A3(net1275),
    .B1(\t$4616 ),
    .B2(\notblock$4615[0] ),
    .X(\sel_0$4617 ));
 sky130_fd_sc_hd__a22o_1 \U$$4150  (.A1(net1160),
    .A2(net436),
    .B1(net1152),
    .B2(net718),
    .X(\t$6526 ));
 sky130_fd_sc_hd__xor2_1 \U$$4151  (.A(\t$6526 ),
    .B(net1267),
    .X(booth_b60_m17));
 sky130_fd_sc_hd__a22o_1 \U$$4152  (.A1(net1152),
    .A2(net434),
    .B1(net1142),
    .B2(net716),
    .X(\t$6527 ));
 sky130_fd_sc_hd__xor2_1 \U$$4153  (.A(\t$6527 ),
    .B(net1263),
    .X(booth_b60_m18));
 sky130_fd_sc_hd__a22o_1 \U$$4154  (.A1(net1142),
    .A2(net436),
    .B1(net1135),
    .B2(net718),
    .X(\t$6528 ));
 sky130_fd_sc_hd__xor2_1 \U$$4155  (.A(\t$6528 ),
    .B(net1267),
    .X(booth_b60_m19));
 sky130_fd_sc_hd__a22o_1 \U$$4156  (.A1(net1136),
    .A2(net435),
    .B1(net1120),
    .B2(net717),
    .X(\t$6529 ));
 sky130_fd_sc_hd__xor2_1 \U$$4157  (.A(\t$6529 ),
    .B(net1267),
    .X(booth_b60_m20));
 sky130_fd_sc_hd__a22o_1 \U$$4158  (.A1(net1119),
    .A2(net436),
    .B1(net1112),
    .B2(net718),
    .X(\t$6530 ));
 sky130_fd_sc_hd__xor2_1 \U$$4159  (.A(\t$6530 ),
    .B(net1263),
    .X(booth_b60_m21));
 sky130_fd_sc_hd__xor2_1 \U$$416  (.A(net61),
    .B(net1275),
    .X(\sel_1$4618 ));
 sky130_fd_sc_hd__a22o_1 \U$$4160  (.A1(net1112),
    .A2(net436),
    .B1(net1103),
    .B2(net718),
    .X(\t$6531 ));
 sky130_fd_sc_hd__xor2_1 \U$$4161  (.A(\t$6531 ),
    .B(net1268),
    .X(booth_b60_m22));
 sky130_fd_sc_hd__a22o_1 \U$$4162  (.A1(net1103),
    .A2(net436),
    .B1(net1095),
    .B2(net718),
    .X(\t$6532 ));
 sky130_fd_sc_hd__xor2_1 \U$$4163  (.A(\t$6532 ),
    .B(net1268),
    .X(booth_b60_m23));
 sky130_fd_sc_hd__a22o_1 \U$$4164  (.A1(net1095),
    .A2(net436),
    .B1(net1085),
    .B2(net718),
    .X(\t$6533 ));
 sky130_fd_sc_hd__xor2_1 \U$$4165  (.A(\t$6533 ),
    .B(net1268),
    .X(booth_b60_m24));
 sky130_fd_sc_hd__a22o_1 \U$$4166  (.A1(net1085),
    .A2(net436),
    .B1(net1077),
    .B2(net718),
    .X(\t$6534 ));
 sky130_fd_sc_hd__xor2_1 \U$$4167  (.A(\t$6534 ),
    .B(net1268),
    .X(booth_b60_m25));
 sky130_fd_sc_hd__a22o_1 \U$$4168  (.A1(net1077),
    .A2(net436),
    .B1(net1069),
    .B2(net718),
    .X(\t$6535 ));
 sky130_fd_sc_hd__xor2_1 \U$$4169  (.A(\t$6535 ),
    .B(net1268),
    .X(booth_b60_m26));
 sky130_fd_sc_hd__a22o_1 \U$$417  (.A1(net1806),
    .A2(net429),
    .B1(net1231),
    .B2(net711),
    .X(\t$4619 ));
 sky130_fd_sc_hd__a22o_1 \U$$4170  (.A1(net1069),
    .A2(net435),
    .B1(net1061),
    .B2(net717),
    .X(\t$6536 ));
 sky130_fd_sc_hd__xor2_1 \U$$4171  (.A(\t$6536 ),
    .B(net1266),
    .X(booth_b60_m27));
 sky130_fd_sc_hd__a22o_1 \U$$4172  (.A1(net1062),
    .A2(net435),
    .B1(net1053),
    .B2(net717),
    .X(\t$6537 ));
 sky130_fd_sc_hd__xor2_1 \U$$4173  (.A(\t$6537 ),
    .B(net1265),
    .X(booth_b60_m28));
 sky130_fd_sc_hd__a22o_1 \U$$4174  (.A1(net1053),
    .A2(net437),
    .B1(net1045),
    .B2(net719),
    .X(\t$6538 ));
 sky130_fd_sc_hd__xor2_1 \U$$4175  (.A(\t$6538 ),
    .B(net1264),
    .X(booth_b60_m29));
 sky130_fd_sc_hd__a22o_1 \U$$4176  (.A1(net1045),
    .A2(net439),
    .B1(net1029),
    .B2(net721),
    .X(\t$6539 ));
 sky130_fd_sc_hd__xor2_1 \U$$4177  (.A(\t$6539 ),
    .B(net1270),
    .X(booth_b60_m30));
 sky130_fd_sc_hd__a22o_1 \U$$4178  (.A1(net1029),
    .A2(net438),
    .B1(net1021),
    .B2(net720),
    .X(\t$6540 ));
 sky130_fd_sc_hd__xor2_1 \U$$4179  (.A(\t$6540 ),
    .B(net1269),
    .X(booth_b60_m31));
 sky130_fd_sc_hd__xor2_1 \U$$418  (.A(\t$4619 ),
    .B(net1248),
    .X(booth_b6_m0));
 sky130_fd_sc_hd__a22o_1 \U$$4180  (.A1(net1021),
    .A2(net441),
    .B1(net1004),
    .B2(net723),
    .X(\t$6541 ));
 sky130_fd_sc_hd__xor2_1 \U$$4181  (.A(\t$6541 ),
    .B(net1269),
    .X(booth_b60_m32));
 sky130_fd_sc_hd__a22o_1 \U$$4182  (.A1(net1004),
    .A2(net437),
    .B1(net996),
    .B2(net719),
    .X(\t$6542 ));
 sky130_fd_sc_hd__xor2_1 \U$$4183  (.A(\t$6542 ),
    .B(net1272),
    .X(booth_b60_m33));
 sky130_fd_sc_hd__a22o_1 \U$$4184  (.A1(net996),
    .A2(net441),
    .B1(net988),
    .B2(net723),
    .X(\t$6543 ));
 sky130_fd_sc_hd__xor2_1 \U$$4185  (.A(\t$6543 ),
    .B(net1272),
    .X(booth_b60_m34));
 sky130_fd_sc_hd__a22o_1 \U$$4186  (.A1(net988),
    .A2(net438),
    .B1(net979),
    .B2(net720),
    .X(\t$6544 ));
 sky130_fd_sc_hd__xor2_1 \U$$4187  (.A(\t$6544 ),
    .B(net1269),
    .X(booth_b60_m35));
 sky130_fd_sc_hd__a22o_1 \U$$4188  (.A1(net979),
    .A2(net438),
    .B1(net970),
    .B2(net720),
    .X(\t$6545 ));
 sky130_fd_sc_hd__xor2_1 \U$$4189  (.A(\t$6545 ),
    .B(net1269),
    .X(booth_b60_m36));
 sky130_fd_sc_hd__a22o_1 \U$$419  (.A1(net1231),
    .A2(net429),
    .B1(net1127),
    .B2(net711),
    .X(\t$4620 ));
 sky130_fd_sc_hd__a22o_1 \U$$4190  (.A1(net971),
    .A2(net438),
    .B1(net962),
    .B2(net720),
    .X(\t$6546 ));
 sky130_fd_sc_hd__xor2_1 \U$$4191  (.A(\t$6546 ),
    .B(net1272),
    .X(booth_b60_m37));
 sky130_fd_sc_hd__a22o_1 \U$$4192  (.A1(net962),
    .A2(net440),
    .B1(net953),
    .B2(net722),
    .X(\t$6547 ));
 sky130_fd_sc_hd__xor2_1 \U$$4193  (.A(\t$6547 ),
    .B(net1271),
    .X(booth_b60_m38));
 sky130_fd_sc_hd__a22o_1 \U$$4194  (.A1(net953),
    .A2(net440),
    .B1(net945),
    .B2(net722),
    .X(\t$6548 ));
 sky130_fd_sc_hd__xor2_1 \U$$4195  (.A(\t$6548 ),
    .B(net1271),
    .X(booth_b60_m39));
 sky130_fd_sc_hd__a22o_1 \U$$4196  (.A1(net945),
    .A2(net440),
    .B1(net929),
    .B2(net722),
    .X(\t$6549 ));
 sky130_fd_sc_hd__xor2_1 \U$$4197  (.A(\t$6549 ),
    .B(net1271),
    .X(booth_b60_m40));
 sky130_fd_sc_hd__a22o_1 \U$$4198  (.A1(net929),
    .A2(net440),
    .B1(net1750),
    .B2(net722),
    .X(\t$6550 ));
 sky130_fd_sc_hd__xor2_1 \U$$4199  (.A(\t$6550 ),
    .B(net1271),
    .X(booth_b60_m41));
 sky130_fd_sc_hd__a22o_1 \U$$42  (.A1(net1147),
    .A2(net442),
    .B1(net1139),
    .B2(net684),
    .X(\t$4428 ));
 sky130_fd_sc_hd__xor2_1 \U$$420  (.A(\t$4620 ),
    .B(net1248),
    .X(booth_b6_m1));
 sky130_fd_sc_hd__a22o_1 \U$$4200  (.A1(net1750),
    .A2(net440),
    .B1(net1743),
    .B2(net722),
    .X(\t$6551 ));
 sky130_fd_sc_hd__xor2_1 \U$$4201  (.A(\t$6551 ),
    .B(net1271),
    .X(booth_b60_m42));
 sky130_fd_sc_hd__a22o_1 \U$$4202  (.A1(net1743),
    .A2(net440),
    .B1(net1735),
    .B2(net722),
    .X(\t$6552 ));
 sky130_fd_sc_hd__xor2_1 \U$$4203  (.A(\t$6552 ),
    .B(net1271),
    .X(booth_b60_m43));
 sky130_fd_sc_hd__a22o_1 \U$$4204  (.A1(net1735),
    .A2(net440),
    .B1(net1727),
    .B2(net722),
    .X(\t$6553 ));
 sky130_fd_sc_hd__xor2_1 \U$$4205  (.A(\t$6553 ),
    .B(net1271),
    .X(booth_b60_m44));
 sky130_fd_sc_hd__a22o_1 \U$$4206  (.A1(net1726),
    .A2(net440),
    .B1(net1717),
    .B2(net722),
    .X(\t$6554 ));
 sky130_fd_sc_hd__xor2_1 \U$$4207  (.A(\t$6554 ),
    .B(net1271),
    .X(booth_b60_m45));
 sky130_fd_sc_hd__a22o_1 \U$$4208  (.A1(net1717),
    .A2(net439),
    .B1(net1708),
    .B2(net721),
    .X(\t$6555 ));
 sky130_fd_sc_hd__xor2_1 \U$$4209  (.A(\t$6555 ),
    .B(net1270),
    .X(booth_b60_m46));
 sky130_fd_sc_hd__a22o_1 \U$$421  (.A1(net1127),
    .A2(net430),
    .B1(net1035),
    .B2(net712),
    .X(\t$4621 ));
 sky130_fd_sc_hd__a22o_1 \U$$4210  (.A1(net1710),
    .A2(net439),
    .B1(net1702),
    .B2(net721),
    .X(\t$6556 ));
 sky130_fd_sc_hd__xor2_1 \U$$4211  (.A(\t$6556 ),
    .B(net1270),
    .X(booth_b60_m47));
 sky130_fd_sc_hd__a22o_1 \U$$4212  (.A1(net1702),
    .A2(net435),
    .B1(net1692),
    .B2(net717),
    .X(\t$6557 ));
 sky130_fd_sc_hd__xor2_1 \U$$4213  (.A(\t$6557 ),
    .B(net1267),
    .X(booth_b60_m48));
 sky130_fd_sc_hd__a22o_1 \U$$4214  (.A1(net1692),
    .A2(net435),
    .B1(net1685),
    .B2(net717),
    .X(\t$6558 ));
 sky130_fd_sc_hd__xor2_1 \U$$4215  (.A(\t$6558 ),
    .B(net1267),
    .X(booth_b60_m49));
 sky130_fd_sc_hd__a22o_1 \U$$4216  (.A1(net1685),
    .A2(net440),
    .B1(net1659),
    .B2(net722),
    .X(\t$6559 ));
 sky130_fd_sc_hd__xor2_1 \U$$4217  (.A(\t$6559 ),
    .B(net1270),
    .X(booth_b60_m50));
 sky130_fd_sc_hd__a22o_1 \U$$4218  (.A1(net1659),
    .A2(net439),
    .B1(net1651),
    .B2(net721),
    .X(\t$6560 ));
 sky130_fd_sc_hd__xor2_1 \U$$4219  (.A(\t$6560 ),
    .B(net1270),
    .X(booth_b60_m51));
 sky130_fd_sc_hd__xor2_1 \U$$422  (.A(\t$4621 ),
    .B(net1248),
    .X(booth_b6_m2));
 sky130_fd_sc_hd__a22o_1 \U$$4220  (.A1(net1651),
    .A2(net439),
    .B1(net1643),
    .B2(net721),
    .X(\t$6561 ));
 sky130_fd_sc_hd__xor2_1 \U$$4221  (.A(\t$6561 ),
    .B(net1270),
    .X(booth_b60_m52));
 sky130_fd_sc_hd__a22o_1 \U$$4222  (.A1(net1643),
    .A2(net439),
    .B1(net1634),
    .B2(net721),
    .X(\t$6562 ));
 sky130_fd_sc_hd__xor2_1 \U$$4223  (.A(\t$6562 ),
    .B(net1270),
    .X(booth_b60_m53));
 sky130_fd_sc_hd__a22o_1 \U$$4224  (.A1(net1636),
    .A2(net439),
    .B1(net1625),
    .B2(net721),
    .X(\t$6563 ));
 sky130_fd_sc_hd__xor2_1 \U$$4225  (.A(\t$6563 ),
    .B(net1270),
    .X(booth_b60_m54));
 sky130_fd_sc_hd__a22o_1 \U$$4226  (.A1(net1625),
    .A2(net439),
    .B1(net1617),
    .B2(net721),
    .X(\t$6564 ));
 sky130_fd_sc_hd__xor2_1 \U$$4227  (.A(\t$6564 ),
    .B(net1270),
    .X(booth_b60_m55));
 sky130_fd_sc_hd__a22o_1 \U$$4228  (.A1(net1619),
    .A2(net439),
    .B1(net1610),
    .B2(net721),
    .X(\t$6565 ));
 sky130_fd_sc_hd__xor2_1 \U$$4229  (.A(\t$6565 ),
    .B(net1270),
    .X(booth_b60_m56));
 sky130_fd_sc_hd__a22o_1 \U$$423  (.A1(net1035),
    .A2(net430),
    .B1(net937),
    .B2(net712),
    .X(\t$4622 ));
 sky130_fd_sc_hd__a22o_1 \U$$4230  (.A1(net1606),
    .A2(net435),
    .B1(net1598),
    .B2(net717),
    .X(\t$6566 ));
 sky130_fd_sc_hd__xor2_1 \U$$4231  (.A(\t$6566 ),
    .B(net1265),
    .X(booth_b60_m57));
 sky130_fd_sc_hd__a22o_1 \U$$4232  (.A1(net1601),
    .A2(net435),
    .B1(net1592),
    .B2(net717),
    .X(\t$6567 ));
 sky130_fd_sc_hd__xor2_1 \U$$4233  (.A(\t$6567 ),
    .B(net1265),
    .X(booth_b60_m58));
 sky130_fd_sc_hd__a22o_1 \U$$4234  (.A1(net1589),
    .A2(net435),
    .B1(net1580),
    .B2(net717),
    .X(\t$6568 ));
 sky130_fd_sc_hd__xor2_1 \U$$4235  (.A(\t$6568 ),
    .B(net1265),
    .X(booth_b60_m59));
 sky130_fd_sc_hd__a22o_1 \U$$4236  (.A1(net1580),
    .A2(net436),
    .B1(net1554),
    .B2(net718),
    .X(\t$6569 ));
 sky130_fd_sc_hd__xor2_1 \U$$4237  (.A(\t$6569 ),
    .B(net1265),
    .X(booth_b60_m60));
 sky130_fd_sc_hd__a22o_1 \U$$4238  (.A1(net1554),
    .A2(net437),
    .B1(net1545),
    .B2(net719),
    .X(\t$6570 ));
 sky130_fd_sc_hd__xor2_1 \U$$4239  (.A(\t$6570 ),
    .B(net1265),
    .X(booth_b60_m61));
 sky130_fd_sc_hd__xor2_1 \U$$424  (.A(\t$4622 ),
    .B(net1248),
    .X(booth_b6_m3));
 sky130_fd_sc_hd__a22o_1 \U$$4240  (.A1(net1549),
    .A2(net439),
    .B1(net1541),
    .B2(net721),
    .X(\t$6571 ));
 sky130_fd_sc_hd__xor2_1 \U$$4241  (.A(\t$6571 ),
    .B(net1271),
    .X(booth_b60_m62));
 sky130_fd_sc_hd__a22o_1 \U$$4242  (.A1(net1537),
    .A2(net435),
    .B1(net1529),
    .B2(net717),
    .X(\t$6572 ));
 sky130_fd_sc_hd__xor2_1 \U$$4243  (.A(\t$6572 ),
    .B(net1266),
    .X(booth_b60_m63));
 sky130_fd_sc_hd__a22o_1 \U$$4244  (.A1(net1529),
    .A2(net435),
    .B1(net1807),
    .B2(net717),
    .X(\t$6573 ));
 sky130_fd_sc_hd__xor2_1 \U$$4245  (.A(\t$6573 ),
    .B(net1265),
    .X(booth_b60_m64));
 sky130_fd_sc_hd__inv_1 \U$$4246  (.A(net1268),
    .Y(\notsign$6574 ));
 sky130_fd_sc_hd__inv_1 \U$$4247  (.A(net1265),
    .Y(\notblock$6575[0] ));
 sky130_fd_sc_hd__inv_1 \U$$4248  (.A(net59),
    .Y(\notblock$6575[1] ));
 sky130_fd_sc_hd__inv_1 \U$$4249  (.A(net1256),
    .Y(\notblock$6575[2] ));
 sky130_fd_sc_hd__a22o_1 \U$$425  (.A1(net936),
    .A2(net430),
    .B1(net1676),
    .B2(net712),
    .X(\t$4623 ));
 sky130_fd_sc_hd__and2_1 \U$$4250  (.A(net1256),
    .B(\notblock$6575[1] ),
    .X(\t$6576 ));
 sky130_fd_sc_hd__a32o_1 \U$$4251  (.A1(\notblock$6575[2] ),
    .A2(net59),
    .A3(net1266),
    .B1(\t$6576 ),
    .B2(\notblock$6575[0] ),
    .X(\sel_0$6577 ));
 sky130_fd_sc_hd__xor2_2 \U$$4252  (.A(net59),
    .B(net1266),
    .X(\sel_1$6578 ));
 sky130_fd_sc_hd__a22o_1 \U$$4253  (.A1(net1808),
    .A2(net421),
    .B1(net1233),
    .B2(net703),
    .X(\t$6579 ));
 sky130_fd_sc_hd__xor2_1 \U$$4254  (.A(\t$6579 ),
    .B(net1254),
    .X(booth_b62_m0));
 sky130_fd_sc_hd__a22o_1 \U$$4255  (.A1(net1234),
    .A2(net421),
    .B1(net1125),
    .B2(net703),
    .X(\t$6580 ));
 sky130_fd_sc_hd__xor2_1 \U$$4256  (.A(\t$6580 ),
    .B(net1254),
    .X(booth_b62_m1));
 sky130_fd_sc_hd__a22o_1 \U$$4257  (.A1(net1129),
    .A2(net422),
    .B1(net1037),
    .B2(net704),
    .X(\t$6581 ));
 sky130_fd_sc_hd__xor2_1 \U$$4258  (.A(\t$6581 ),
    .B(net1259),
    .X(booth_b62_m2));
 sky130_fd_sc_hd__a22o_1 \U$$4259  (.A1(net1037),
    .A2(net422),
    .B1(net938),
    .B2(net704),
    .X(\t$6582 ));
 sky130_fd_sc_hd__xor2_1 \U$$426  (.A(\t$4623 ),
    .B(net1248),
    .X(booth_b6_m4));
 sky130_fd_sc_hd__xor2_1 \U$$4260  (.A(\t$6582 ),
    .B(net1259),
    .X(booth_b62_m3));
 sky130_fd_sc_hd__a22o_1 \U$$4261  (.A1(net939),
    .A2(net422),
    .B1(net1678),
    .B2(net704),
    .X(\t$6583 ));
 sky130_fd_sc_hd__xor2_1 \U$$4262  (.A(\t$6583 ),
    .B(net1259),
    .X(booth_b62_m4));
 sky130_fd_sc_hd__a22o_1 \U$$4263  (.A1(net1678),
    .A2(net422),
    .B1(net1567),
    .B2(net704),
    .X(\t$6584 ));
 sky130_fd_sc_hd__xor2_1 \U$$4264  (.A(\t$6584 ),
    .B(net1259),
    .X(booth_b62_m5));
 sky130_fd_sc_hd__a22o_1 \U$$4265  (.A1(net1567),
    .A2(net422),
    .B1(net1526),
    .B2(net704),
    .X(\t$6585 ));
 sky130_fd_sc_hd__xor2_1 \U$$4266  (.A(\t$6585 ),
    .B(net1259),
    .X(booth_b62_m6));
 sky130_fd_sc_hd__a22o_1 \U$$4267  (.A1(net1526),
    .A2(net422),
    .B1(net1518),
    .B2(net704),
    .X(\t$6586 ));
 sky130_fd_sc_hd__xor2_1 \U$$4268  (.A(\t$6586 ),
    .B(net1259),
    .X(booth_b62_m7));
 sky130_fd_sc_hd__a22o_1 \U$$4269  (.A1(net1518),
    .A2(net421),
    .B1(net1507),
    .B2(net703),
    .X(\t$6587 ));
 sky130_fd_sc_hd__a22o_1 \U$$427  (.A1(net1676),
    .A2(net430),
    .B1(net1564),
    .B2(net712),
    .X(\t$4624 ));
 sky130_fd_sc_hd__xor2_1 \U$$4270  (.A(\t$6587 ),
    .B(net1254),
    .X(booth_b62_m8));
 sky130_fd_sc_hd__a22o_1 \U$$4271  (.A1(net1507),
    .A2(net418),
    .B1(net1498),
    .B2(net700),
    .X(\t$6588 ));
 sky130_fd_sc_hd__xor2_1 \U$$4272  (.A(\t$6588 ),
    .B(net1258),
    .X(booth_b62_m9));
 sky130_fd_sc_hd__a22o_1 \U$$4273  (.A1(net1502),
    .A2(net418),
    .B1(net1222),
    .B2(net700),
    .X(\t$6589 ));
 sky130_fd_sc_hd__xor2_1 \U$$4274  (.A(\t$6589 ),
    .B(net1254),
    .X(booth_b62_m10));
 sky130_fd_sc_hd__a22o_1 \U$$4275  (.A1(net1222),
    .A2(net418),
    .B1(net1214),
    .B2(net700),
    .X(\t$6590 ));
 sky130_fd_sc_hd__xor2_1 \U$$4276  (.A(\t$6590 ),
    .B(net1254),
    .X(booth_b62_m11));
 sky130_fd_sc_hd__a22o_1 \U$$4277  (.A1(net1214),
    .A2(net418),
    .B1(net1205),
    .B2(net700),
    .X(\t$6591 ));
 sky130_fd_sc_hd__xor2_1 \U$$4278  (.A(\t$6591 ),
    .B(net1254),
    .X(booth_b62_m12));
 sky130_fd_sc_hd__a22o_1 \U$$4279  (.A1(net1205),
    .A2(net418),
    .B1(net1196),
    .B2(net700),
    .X(\t$6592 ));
 sky130_fd_sc_hd__xor2_1 \U$$428  (.A(\t$4624 ),
    .B(net1248),
    .X(booth_b6_m5));
 sky130_fd_sc_hd__xor2_1 \U$$4280  (.A(\t$6592 ),
    .B(net1254),
    .X(booth_b62_m13));
 sky130_fd_sc_hd__a22o_1 \U$$4281  (.A1(net1196),
    .A2(net418),
    .B1(net1177),
    .B2(net700),
    .X(\t$6593 ));
 sky130_fd_sc_hd__xor2_1 \U$$4282  (.A(\t$6593 ),
    .B(net1254),
    .X(booth_b62_m14));
 sky130_fd_sc_hd__a22o_1 \U$$4283  (.A1(net1178),
    .A2(net421),
    .B1(net1169),
    .B2(net703),
    .X(\t$6594 ));
 sky130_fd_sc_hd__xor2_1 \U$$4284  (.A(\t$6594 ),
    .B(net1258),
    .X(booth_b62_m15));
 sky130_fd_sc_hd__a22o_1 \U$$4285  (.A1(net1169),
    .A2(net418),
    .B1(net1160),
    .B2(net700),
    .X(\t$6595 ));
 sky130_fd_sc_hd__xor2_1 \U$$4286  (.A(\t$6595 ),
    .B(net1258),
    .X(booth_b62_m16));
 sky130_fd_sc_hd__a22o_1 \U$$4287  (.A1(net1159),
    .A2(net418),
    .B1(net1152),
    .B2(net700),
    .X(\t$6596 ));
 sky130_fd_sc_hd__xor2_1 \U$$4288  (.A(\t$6596 ),
    .B(net1254),
    .X(booth_b62_m17));
 sky130_fd_sc_hd__a22o_1 \U$$4289  (.A1(net1152),
    .A2(net420),
    .B1(net1142),
    .B2(net702),
    .X(\t$6597 ));
 sky130_fd_sc_hd__a22o_1 \U$$429  (.A1(net1564),
    .A2(net429),
    .B1(net1523),
    .B2(net711),
    .X(\t$4625 ));
 sky130_fd_sc_hd__xor2_1 \U$$4290  (.A(\t$6597 ),
    .B(net1256),
    .X(booth_b62_m18));
 sky130_fd_sc_hd__a22o_1 \U$$4291  (.A1(net1141),
    .A2(net418),
    .B1(net1135),
    .B2(net700),
    .X(\t$6598 ));
 sky130_fd_sc_hd__xor2_1 \U$$4292  (.A(\t$6598 ),
    .B(net1255),
    .X(booth_b62_m19));
 sky130_fd_sc_hd__a22o_1 \U$$4293  (.A1(net1135),
    .A2(net419),
    .B1(net1119),
    .B2(net701),
    .X(\t$6599 ));
 sky130_fd_sc_hd__xor2_1 \U$$4294  (.A(\t$6599 ),
    .B(net1255),
    .X(booth_b62_m20));
 sky130_fd_sc_hd__a22o_1 \U$$4295  (.A1(net1119),
    .A2(net419),
    .B1(net1112),
    .B2(net701),
    .X(\t$6600 ));
 sky130_fd_sc_hd__xor2_1 \U$$4296  (.A(\t$6600 ),
    .B(net1255),
    .X(booth_b62_m21));
 sky130_fd_sc_hd__a22o_1 \U$$4297  (.A1(net1112),
    .A2(net419),
    .B1(net1103),
    .B2(net701),
    .X(\t$6601 ));
 sky130_fd_sc_hd__xor2_1 \U$$4298  (.A(\t$6601 ),
    .B(net1255),
    .X(booth_b62_m22));
 sky130_fd_sc_hd__a22o_1 \U$$4299  (.A1(net1103),
    .A2(net419),
    .B1(net1095),
    .B2(net701),
    .X(\t$6602 ));
 sky130_fd_sc_hd__xor2_1 \U$$43  (.A(\t$4428 ),
    .B(net1569),
    .X(booth_b0_m18));
 sky130_fd_sc_hd__xor2_1 \U$$430  (.A(\t$4625 ),
    .B(net1248),
    .X(booth_b6_m6));
 sky130_fd_sc_hd__xor2_1 \U$$4300  (.A(\t$6602 ),
    .B(net1255),
    .X(booth_b62_m23));
 sky130_fd_sc_hd__a22o_1 \U$$4301  (.A1(net1095),
    .A2(net420),
    .B1(net1085),
    .B2(net702),
    .X(\t$6603 ));
 sky130_fd_sc_hd__xor2_1 \U$$4302  (.A(\t$6603 ),
    .B(net1256),
    .X(booth_b62_m24));
 sky130_fd_sc_hd__a22o_1 \U$$4303  (.A1(net1085),
    .A2(net420),
    .B1(net1077),
    .B2(net702),
    .X(\t$6604 ));
 sky130_fd_sc_hd__xor2_1 \U$$4304  (.A(\t$6604 ),
    .B(net1256),
    .X(booth_b62_m25));
 sky130_fd_sc_hd__a22o_1 \U$$4305  (.A1(net1077),
    .A2(net419),
    .B1(net1069),
    .B2(net701),
    .X(\t$6605 ));
 sky130_fd_sc_hd__xor2_1 \U$$4306  (.A(\t$6605 ),
    .B(net1256),
    .X(booth_b62_m26));
 sky130_fd_sc_hd__a22o_1 \U$$4307  (.A1(net1070),
    .A2(net418),
    .B1(net1062),
    .B2(net700),
    .X(\t$6606 ));
 sky130_fd_sc_hd__xor2_1 \U$$4308  (.A(\t$6606 ),
    .B(net1258),
    .X(booth_b62_m27));
 sky130_fd_sc_hd__a22o_1 \U$$4309  (.A1(net1062),
    .A2(net422),
    .B1(net1053),
    .B2(net704),
    .X(\t$6607 ));
 sky130_fd_sc_hd__a22o_1 \U$$431  (.A1(net1523),
    .A2(net429),
    .B1(net1515),
    .B2(net711),
    .X(\t$4626 ));
 sky130_fd_sc_hd__xor2_1 \U$$4310  (.A(\t$6607 ),
    .B(net1260),
    .X(booth_b62_m28));
 sky130_fd_sc_hd__a22o_1 \U$$4311  (.A1(net1053),
    .A2(net422),
    .B1(net1045),
    .B2(net704),
    .X(\t$6608 ));
 sky130_fd_sc_hd__xor2_1 \U$$4312  (.A(\t$6608 ),
    .B(net1259),
    .X(booth_b62_m29));
 sky130_fd_sc_hd__a22o_1 \U$$4313  (.A1(net1045),
    .A2(net425),
    .B1(net1029),
    .B2(net707),
    .X(\t$6609 ));
 sky130_fd_sc_hd__xor2_1 \U$$4314  (.A(\t$6609 ),
    .B(net1259),
    .X(booth_b62_m30));
 sky130_fd_sc_hd__a22o_1 \U$$4315  (.A1(net1029),
    .A2(net422),
    .B1(net1021),
    .B2(net704),
    .X(\t$6610 ));
 sky130_fd_sc_hd__xor2_1 \U$$4316  (.A(\t$6610 ),
    .B(net1259),
    .X(booth_b62_m31));
 sky130_fd_sc_hd__a22o_1 \U$$4317  (.A1(net1021),
    .A2(net422),
    .B1(net1004),
    .B2(net704),
    .X(\t$6611 ));
 sky130_fd_sc_hd__xor2_1 \U$$4318  (.A(\t$6611 ),
    .B(net1259),
    .X(booth_b62_m32));
 sky130_fd_sc_hd__a22o_1 \U$$4319  (.A1(net1004),
    .A2(net425),
    .B1(net996),
    .B2(net707),
    .X(\t$6612 ));
 sky130_fd_sc_hd__xor2_1 \U$$432  (.A(\t$4626 ),
    .B(net1248),
    .X(booth_b6_m7));
 sky130_fd_sc_hd__xor2_1 \U$$4320  (.A(\t$6612 ),
    .B(net1262),
    .X(booth_b62_m33));
 sky130_fd_sc_hd__a22o_1 \U$$4321  (.A1(net996),
    .A2(net425),
    .B1(net989),
    .B2(net707),
    .X(\t$6613 ));
 sky130_fd_sc_hd__xor2_1 \U$$4322  (.A(\t$6613 ),
    .B(net1262),
    .X(booth_b62_m34));
 sky130_fd_sc_hd__a22o_1 \U$$4323  (.A1(net989),
    .A2(net423),
    .B1(net980),
    .B2(net705),
    .X(\t$6614 ));
 sky130_fd_sc_hd__xor2_1 \U$$4324  (.A(\t$6614 ),
    .B(net1261),
    .X(booth_b62_m35));
 sky130_fd_sc_hd__a22o_1 \U$$4325  (.A1(net980),
    .A2(net424),
    .B1(net971),
    .B2(net706),
    .X(\t$6615 ));
 sky130_fd_sc_hd__xor2_1 \U$$4326  (.A(\t$6615 ),
    .B(net1261),
    .X(booth_b62_m36));
 sky130_fd_sc_hd__a22o_1 \U$$4327  (.A1(net971),
    .A2(net424),
    .B1(net963),
    .B2(net706),
    .X(\t$6616 ));
 sky130_fd_sc_hd__xor2_1 \U$$4328  (.A(\t$6616 ),
    .B(net1261),
    .X(booth_b62_m37));
 sky130_fd_sc_hd__a22o_1 \U$$4329  (.A1(net963),
    .A2(net424),
    .B1(net953),
    .B2(net706),
    .X(\t$6617 ));
 sky130_fd_sc_hd__a22o_1 \U$$433  (.A1(net1513),
    .A2(net431),
    .B1(net1505),
    .B2(net713),
    .X(\t$4627 ));
 sky130_fd_sc_hd__xor2_1 \U$$4330  (.A(\t$6617 ),
    .B(net1261),
    .X(booth_b62_m38));
 sky130_fd_sc_hd__a22o_1 \U$$4331  (.A1(net953),
    .A2(net424),
    .B1(net945),
    .B2(net706),
    .X(\t$6618 ));
 sky130_fd_sc_hd__xor2_1 \U$$4332  (.A(\t$6618 ),
    .B(net1261),
    .X(booth_b62_m39));
 sky130_fd_sc_hd__a22o_1 \U$$4333  (.A1(net945),
    .A2(net424),
    .B1(net929),
    .B2(net706),
    .X(\t$6619 ));
 sky130_fd_sc_hd__xor2_1 \U$$4334  (.A(\t$6619 ),
    .B(net1261),
    .X(booth_b62_m40));
 sky130_fd_sc_hd__a22o_1 \U$$4335  (.A1(net929),
    .A2(net423),
    .B1(net1750),
    .B2(net705),
    .X(\t$6620 ));
 sky130_fd_sc_hd__xor2_1 \U$$4336  (.A(\t$6620 ),
    .B(net1261),
    .X(booth_b62_m41));
 sky130_fd_sc_hd__a22o_1 \U$$4337  (.A1(net1751),
    .A2(net424),
    .B1(net1743),
    .B2(net706),
    .X(\t$6621 ));
 sky130_fd_sc_hd__xor2_1 \U$$4338  (.A(\t$6621 ),
    .B(net1262),
    .X(booth_b62_m42));
 sky130_fd_sc_hd__a22o_1 \U$$4339  (.A1(net1742),
    .A2(net424),
    .B1(net1734),
    .B2(net706),
    .X(\t$6622 ));
 sky130_fd_sc_hd__xor2_1 \U$$434  (.A(\t$4627 ),
    .B(net1250),
    .X(booth_b6_m8));
 sky130_fd_sc_hd__xor2_1 \U$$4340  (.A(\t$6622 ),
    .B(net1262),
    .X(booth_b62_m43));
 sky130_fd_sc_hd__a22o_1 \U$$4341  (.A1(net1731),
    .A2(net419),
    .B1(net1722),
    .B2(net701),
    .X(\t$6623 ));
 sky130_fd_sc_hd__xor2_1 \U$$4342  (.A(\t$6623 ),
    .B(net1255),
    .X(booth_b62_m44));
 sky130_fd_sc_hd__a22o_1 \U$$4343  (.A1(net1727),
    .A2(net423),
    .B1(net1719),
    .B2(net705),
    .X(\t$6624 ));
 sky130_fd_sc_hd__xor2_1 \U$$4344  (.A(\t$6624 ),
    .B(net1260),
    .X(booth_b62_m45));
 sky130_fd_sc_hd__a22o_1 \U$$4345  (.A1(net1719),
    .A2(net420),
    .B1(net1710),
    .B2(net702),
    .X(\t$6625 ));
 sky130_fd_sc_hd__xor2_1 \U$$4346  (.A(\t$6625 ),
    .B(net1256),
    .X(booth_b62_m46));
 sky130_fd_sc_hd__a22o_1 \U$$4347  (.A1(net1710),
    .A2(net423),
    .B1(net1702),
    .B2(net705),
    .X(\t$6626 ));
 sky130_fd_sc_hd__xor2_1 \U$$4348  (.A(\t$6626 ),
    .B(net1260),
    .X(booth_b62_m47));
 sky130_fd_sc_hd__a22o_1 \U$$4349  (.A1(net1702),
    .A2(net420),
    .B1(net1692),
    .B2(net702),
    .X(\t$6627 ));
 sky130_fd_sc_hd__a22o_1 \U$$435  (.A1(net1505),
    .A2(net431),
    .B1(net1496),
    .B2(net713),
    .X(\t$4628 ));
 sky130_fd_sc_hd__xor2_1 \U$$4350  (.A(\t$6627 ),
    .B(net1256),
    .X(booth_b62_m48));
 sky130_fd_sc_hd__a22o_1 \U$$4351  (.A1(net1692),
    .A2(net423),
    .B1(net1685),
    .B2(net705),
    .X(\t$6628 ));
 sky130_fd_sc_hd__xor2_1 \U$$4352  (.A(\t$6628 ),
    .B(net1260),
    .X(booth_b62_m49));
 sky130_fd_sc_hd__a22o_1 \U$$4353  (.A1(net1680),
    .A2(net419),
    .B1(net1655),
    .B2(net701),
    .X(\t$6629 ));
 sky130_fd_sc_hd__xor2_1 \U$$4354  (.A(\t$6629 ),
    .B(net1255),
    .X(booth_b62_m50));
 sky130_fd_sc_hd__a22o_1 \U$$4355  (.A1(net1659),
    .A2(net423),
    .B1(net1651),
    .B2(net705),
    .X(\t$6630 ));
 sky130_fd_sc_hd__xor2_1 \U$$4356  (.A(\t$6630 ),
    .B(net1260),
    .X(booth_b62_m51));
 sky130_fd_sc_hd__a22o_1 \U$$4357  (.A1(net1653),
    .A2(net423),
    .B1(net1645),
    .B2(net705),
    .X(\t$6631 ));
 sky130_fd_sc_hd__xor2_1 \U$$4358  (.A(\t$6631 ),
    .B(net1260),
    .X(booth_b62_m52));
 sky130_fd_sc_hd__a22o_1 \U$$4359  (.A1(net1645),
    .A2(net423),
    .B1(net1636),
    .B2(net705),
    .X(\t$6632 ));
 sky130_fd_sc_hd__xor2_1 \U$$436  (.A(\t$4628 ),
    .B(net1250),
    .X(booth_b6_m9));
 sky130_fd_sc_hd__xor2_1 \U$$4360  (.A(\t$6632 ),
    .B(net1260),
    .X(booth_b62_m53));
 sky130_fd_sc_hd__a22o_1 \U$$4361  (.A1(net1636),
    .A2(net424),
    .B1(net1625),
    .B2(net706),
    .X(\t$6633 ));
 sky130_fd_sc_hd__xor2_1 \U$$4362  (.A(\t$6633 ),
    .B(net1262),
    .X(booth_b62_m54));
 sky130_fd_sc_hd__a22o_1 \U$$4363  (.A1(net1628),
    .A2(net420),
    .B1(net1617),
    .B2(net702),
    .X(\t$6634 ));
 sky130_fd_sc_hd__xor2_1 \U$$4364  (.A(\t$6634 ),
    .B(net1256),
    .X(booth_b62_m55));
 sky130_fd_sc_hd__a22o_1 \U$$4365  (.A1(net1617),
    .A2(net420),
    .B1(net1610),
    .B2(net702),
    .X(\t$6635 ));
 sky130_fd_sc_hd__xor2_1 \U$$4366  (.A(\t$6635 ),
    .B(net1260),
    .X(booth_b62_m56));
 sky130_fd_sc_hd__a22o_1 \U$$4367  (.A1(net1610),
    .A2(net423),
    .B1(net1601),
    .B2(net705),
    .X(\t$6636 ));
 sky130_fd_sc_hd__xor2_1 \U$$4368  (.A(\t$6636 ),
    .B(net1261),
    .X(booth_b62_m57));
 sky130_fd_sc_hd__a22o_1 \U$$4369  (.A1(net1598),
    .A2(net420),
    .B1(net1589),
    .B2(net702),
    .X(\t$6637 ));
 sky130_fd_sc_hd__a22o_1 \U$$437  (.A1(net1496),
    .A2(net427),
    .B1(net1221),
    .B2(net709),
    .X(\t$4629 ));
 sky130_fd_sc_hd__xor2_1 \U$$4370  (.A(\t$6637 ),
    .B(net1257),
    .X(booth_b62_m58));
 sky130_fd_sc_hd__a22o_1 \U$$4371  (.A1(net1588),
    .A2(net419),
    .B1(net1579),
    .B2(net701),
    .X(\t$6638 ));
 sky130_fd_sc_hd__xor2_1 \U$$4372  (.A(\t$6638 ),
    .B(net1255),
    .X(booth_b62_m59));
 sky130_fd_sc_hd__a22o_1 \U$$4373  (.A1(net1584),
    .A2(net423),
    .B1(net1557),
    .B2(net705),
    .X(\t$6639 ));
 sky130_fd_sc_hd__xor2_1 \U$$4374  (.A(\t$6639 ),
    .B(net1261),
    .X(booth_b62_m60));
 sky130_fd_sc_hd__a22o_1 \U$$4375  (.A1(net1554),
    .A2(net420),
    .B1(net1545),
    .B2(net702),
    .X(\t$6640 ));
 sky130_fd_sc_hd__xor2_1 \U$$4376  (.A(\t$6640 ),
    .B(net1257),
    .X(booth_b62_m61));
 sky130_fd_sc_hd__a22o_1 \U$$4377  (.A1(net1545),
    .A2(net420),
    .B1(net1537),
    .B2(net702),
    .X(\t$6641 ));
 sky130_fd_sc_hd__xor2_1 \U$$4378  (.A(\t$6641 ),
    .B(net1257),
    .X(booth_b62_m62));
 sky130_fd_sc_hd__a22o_1 \U$$4379  (.A1(net1536),
    .A2(net419),
    .B1(net1528),
    .B2(net701),
    .X(\t$6642 ));
 sky130_fd_sc_hd__xor2_1 \U$$438  (.A(\t$4629 ),
    .B(net1245),
    .X(booth_b6_m10));
 sky130_fd_sc_hd__xor2_1 \U$$4380  (.A(\t$6642 ),
    .B(net1255),
    .X(booth_b62_m63));
 sky130_fd_sc_hd__a22o_1 \U$$4381  (.A1(net1528),
    .A2(net419),
    .B1(net1809),
    .B2(net701),
    .X(\t$6643 ));
 sky130_fd_sc_hd__xor2_1 \U$$4382  (.A(\t$6643 ),
    .B(net1255),
    .X(booth_b62_m64));
 sky130_fd_sc_hd__inv_1 \U$$4383  (.A(net1257),
    .Y(\notsign$6644 ));
 sky130_fd_sc_hd__inv_1 \U$$4384  (.A(net1260),
    .Y(\notblock$6645[0] ));
 sky130_fd_sc_hd__inv_1 \U$$4385  (.A(net1810),
    .Y(\notblock$6645[1] ));
 sky130_fd_sc_hd__inv_1 \U$$4386  (.A(net1811),
    .Y(\notblock$6645[2] ));
 sky130_fd_sc_hd__and2_1 \U$$4387  (.A(net1812),
    .B(\notblock$6645[1] ),
    .X(\t$6646 ));
 sky130_fd_sc_hd__a32o_1 \U$$4388  (.A1(\notblock$6645[2] ),
    .A2(net1813),
    .A3(net1260),
    .B1(\t$6646 ),
    .B2(\notblock$6645[0] ),
    .X(\sel_0$6647 ));
 sky130_fd_sc_hd__xor2_2 \U$$4389  (.A(net1814),
    .B(net1256),
    .X(\sel_1$6648 ));
 sky130_fd_sc_hd__a22o_1 \U$$439  (.A1(net1221),
    .A2(net427),
    .B1(net1211),
    .B2(net709),
    .X(\t$4630 ));
 sky130_fd_sc_hd__a22o_1 \U$$4390  (.A1(net1815),
    .A2(\sel_0$6647 ),
    .B1(net1233),
    .B2(net698),
    .X(\t$6649 ));
 sky130_fd_sc_hd__xor2_1 \U$$4391  (.A(\t$6649 ),
    .B(net1816),
    .X(booth_b64_m0));
 sky130_fd_sc_hd__a22o_1 \U$$4392  (.A1(net1234),
    .A2(\sel_0$6647 ),
    .B1(net1129),
    .B2(net698),
    .X(\t$6650 ));
 sky130_fd_sc_hd__xor2_1 \U$$4393  (.A(\t$6650 ),
    .B(net1817),
    .X(booth_b64_m1));
 sky130_fd_sc_hd__a22o_1 \U$$4394  (.A1(net76),
    .A2(\sel_0$6647 ),
    .B1(net1038),
    .B2(net698),
    .X(\t$6651 ));
 sky130_fd_sc_hd__xor2_1 \U$$4395  (.A(\t$6651 ),
    .B(net1818),
    .X(booth_b64_m2));
 sky130_fd_sc_hd__a22o_1 \U$$4396  (.A1(net1038),
    .A2(\sel_0$6647 ),
    .B1(net939),
    .B2(net698),
    .X(\t$6652 ));
 sky130_fd_sc_hd__xor2_1 \U$$4397  (.A(\t$6652 ),
    .B(net1819),
    .X(booth_b64_m3));
 sky130_fd_sc_hd__a22o_1 \U$$4398  (.A1(net939),
    .A2(\sel_0$6647 ),
    .B1(net1678),
    .B2(net698),
    .X(\t$6653 ));
 sky130_fd_sc_hd__xor2_1 \U$$4399  (.A(\t$6653 ),
    .B(net1820),
    .X(booth_b64_m4));
 sky130_fd_sc_hd__a22o_1 \U$$44  (.A1(net1143),
    .A2(net448),
    .B1(net1133),
    .B2(net690),
    .X(\t$4429 ));
 sky130_fd_sc_hd__xor2_1 \U$$440  (.A(\t$4630 ),
    .B(net1245),
    .X(booth_b6_m11));
 sky130_fd_sc_hd__a22o_1 \U$$4400  (.A1(net1677),
    .A2(\sel_0$6647 ),
    .B1(net1566),
    .B2(net696),
    .X(\t$6654 ));
 sky130_fd_sc_hd__xor2_1 \U$$4401  (.A(\t$6654 ),
    .B(net1821),
    .X(booth_b64_m5));
 sky130_fd_sc_hd__a22o_1 \U$$4402  (.A1(net1563),
    .A2(\sel_0$6647 ),
    .B1(net125),
    .B2(net695),
    .X(\t$6655 ));
 sky130_fd_sc_hd__xor2_1 \U$$4403  (.A(\t$6655 ),
    .B(net1822),
    .X(booth_b64_m6));
 sky130_fd_sc_hd__a22o_1 \U$$4404  (.A1(net125),
    .A2(\sel_0$6647 ),
    .B1(net1518),
    .B2(net696),
    .X(\t$6656 ));
 sky130_fd_sc_hd__xor2_1 \U$$4405  (.A(\t$6656 ),
    .B(net1823),
    .X(booth_b64_m7));
 sky130_fd_sc_hd__a22o_1 \U$$4406  (.A1(net1518),
    .A2(\sel_0$6647 ),
    .B1(net1507),
    .B2(net694),
    .X(\t$6657 ));
 sky130_fd_sc_hd__xor2_1 \U$$4407  (.A(\t$6657 ),
    .B(net1824),
    .X(booth_b64_m8));
 sky130_fd_sc_hd__a22o_1 \U$$4408  (.A1(net1507),
    .A2(\sel_0$6647 ),
    .B1(net1502),
    .B2(net694),
    .X(\t$6658 ));
 sky130_fd_sc_hd__xor2_1 \U$$4409  (.A(\t$6658 ),
    .B(net1825),
    .X(booth_b64_m9));
 sky130_fd_sc_hd__a22o_1 \U$$441  (.A1(net1211),
    .A2(net431),
    .B1(net1203),
    .B2(net713),
    .X(\t$4631 ));
 sky130_fd_sc_hd__a22o_1 \U$$4410  (.A1(net1502),
    .A2(\sel_0$6647 ),
    .B1(net1222),
    .B2(net694),
    .X(\t$6659 ));
 sky130_fd_sc_hd__xor2_1 \U$$4411  (.A(\t$6659 ),
    .B(net1826),
    .X(booth_b64_m10));
 sky130_fd_sc_hd__a22o_1 \U$$4412  (.A1(net1222),
    .A2(\sel_0$6647 ),
    .B1(net1214),
    .B2(net694),
    .X(\t$6660 ));
 sky130_fd_sc_hd__xor2_1 \U$$4413  (.A(\t$6660 ),
    .B(net1827),
    .X(booth_b64_m11));
 sky130_fd_sc_hd__a22o_1 \U$$4414  (.A1(net1214),
    .A2(\sel_0$6647 ),
    .B1(net1205),
    .B2(net694),
    .X(\t$6661 ));
 sky130_fd_sc_hd__xor2_1 \U$$4415  (.A(\t$6661 ),
    .B(net1828),
    .X(booth_b64_m12));
 sky130_fd_sc_hd__a22o_1 \U$$4416  (.A1(net1209),
    .A2(\sel_0$6647 ),
    .B1(net1197),
    .B2(net695),
    .X(\t$6662 ));
 sky130_fd_sc_hd__xor2_1 \U$$4417  (.A(\t$6662 ),
    .B(net1829),
    .X(booth_b64_m13));
 sky130_fd_sc_hd__a22o_1 \U$$4418  (.A1(net1196),
    .A2(\sel_0$6647 ),
    .B1(net1177),
    .B2(net694),
    .X(\t$6663 ));
 sky130_fd_sc_hd__xor2_1 \U$$4419  (.A(\t$6663 ),
    .B(net1830),
    .X(booth_b64_m14));
 sky130_fd_sc_hd__xor2_1 \U$$442  (.A(\t$4631 ),
    .B(net1250),
    .X(booth_b6_m12));
 sky130_fd_sc_hd__a22o_1 \U$$4420  (.A1(net1177),
    .A2(\sel_0$6647 ),
    .B1(net1168),
    .B2(net694),
    .X(\t$6664 ));
 sky130_fd_sc_hd__xor2_1 \U$$4421  (.A(\t$6664 ),
    .B(net1831),
    .X(booth_b64_m15));
 sky130_fd_sc_hd__a22o_1 \U$$4422  (.A1(net1169),
    .A2(\sel_0$6647 ),
    .B1(net1160),
    .B2(net695),
    .X(\t$6665 ));
 sky130_fd_sc_hd__xor2_1 \U$$4423  (.A(\t$6665 ),
    .B(net1832),
    .X(booth_b64_m16));
 sky130_fd_sc_hd__a22o_1 \U$$4424  (.A1(net1159),
    .A2(\sel_0$6647 ),
    .B1(net1152),
    .B2(net693),
    .X(\t$6666 ));
 sky130_fd_sc_hd__xor2_1 \U$$4425  (.A(\t$6666 ),
    .B(net1833),
    .X(booth_b64_m17));
 sky130_fd_sc_hd__a22o_1 \U$$4426  (.A1(net1152),
    .A2(\sel_0$6647 ),
    .B1(net1141),
    .B2(net693),
    .X(\t$6667 ));
 sky130_fd_sc_hd__xor2_1 \U$$4427  (.A(\t$6667 ),
    .B(net1834),
    .X(booth_b64_m18));
 sky130_fd_sc_hd__a22o_1 \U$$4428  (.A1(net1141),
    .A2(\sel_0$6647 ),
    .B1(net1135),
    .B2(net694),
    .X(\t$6668 ));
 sky130_fd_sc_hd__xor2_1 \U$$4429  (.A(\t$6668 ),
    .B(net1835),
    .X(booth_b64_m19));
 sky130_fd_sc_hd__a22o_1 \U$$443  (.A1(net1206),
    .A2(net431),
    .B1(net1198),
    .B2(net713),
    .X(\t$4632 ));
 sky130_fd_sc_hd__a22o_1 \U$$4430  (.A1(net1135),
    .A2(\sel_0$6647 ),
    .B1(net1119),
    .B2(net694),
    .X(\t$6669 ));
 sky130_fd_sc_hd__xor2_1 \U$$4431  (.A(\t$6669 ),
    .B(net1836),
    .X(booth_b64_m20));
 sky130_fd_sc_hd__a22o_1 \U$$4432  (.A1(net1119),
    .A2(\sel_0$6647 ),
    .B1(net1112),
    .B2(net693),
    .X(\t$6670 ));
 sky130_fd_sc_hd__xor2_1 \U$$4433  (.A(\t$6670 ),
    .B(net1837),
    .X(booth_b64_m21));
 sky130_fd_sc_hd__a22o_1 \U$$4434  (.A1(net1112),
    .A2(\sel_0$6647 ),
    .B1(net1103),
    .B2(net695),
    .X(\t$6671 ));
 sky130_fd_sc_hd__xor2_1 \U$$4435  (.A(\t$6671 ),
    .B(net1838),
    .X(booth_b64_m22));
 sky130_fd_sc_hd__a22o_1 \U$$4436  (.A1(net1103),
    .A2(\sel_0$6647 ),
    .B1(net1095),
    .B2(net693),
    .X(\t$6672 ));
 sky130_fd_sc_hd__xor2_1 \U$$4437  (.A(\t$6672 ),
    .B(net1839),
    .X(booth_b64_m23));
 sky130_fd_sc_hd__a22o_1 \U$$4438  (.A1(net1095),
    .A2(\sel_0$6647 ),
    .B1(net1086),
    .B2(net695),
    .X(\t$6673 ));
 sky130_fd_sc_hd__xor2_1 \U$$4439  (.A(\t$6673 ),
    .B(net1840),
    .X(booth_b64_m24));
 sky130_fd_sc_hd__xor2_1 \U$$444  (.A(\t$4632 ),
    .B(net1250),
    .X(booth_b6_m13));
 sky130_fd_sc_hd__a22o_1 \U$$4440  (.A1(net1086),
    .A2(\sel_0$6647 ),
    .B1(net1076),
    .B2(net695),
    .X(\t$6674 ));
 sky130_fd_sc_hd__xor2_1 \U$$4441  (.A(\t$6674 ),
    .B(net1841),
    .X(booth_b64_m25));
 sky130_fd_sc_hd__a22o_1 \U$$4442  (.A1(net1078),
    .A2(\sel_0$6647 ),
    .B1(net1070),
    .B2(net698),
    .X(\t$6675 ));
 sky130_fd_sc_hd__xor2_1 \U$$4443  (.A(\t$6675 ),
    .B(net1842),
    .X(booth_b64_m26));
 sky130_fd_sc_hd__a22o_1 \U$$4444  (.A1(net1070),
    .A2(\sel_0$6647 ),
    .B1(net1062),
    .B2(net698),
    .X(\t$6676 ));
 sky130_fd_sc_hd__xor2_1 \U$$4445  (.A(\t$6676 ),
    .B(net1843),
    .X(booth_b64_m27));
 sky130_fd_sc_hd__a22o_1 \U$$4446  (.A1(net84),
    .A2(\sel_0$6647 ),
    .B1(net1054),
    .B2(net698),
    .X(\t$6677 ));
 sky130_fd_sc_hd__xor2_1 \U$$4447  (.A(\t$6677 ),
    .B(net1844),
    .X(booth_b64_m28));
 sky130_fd_sc_hd__a22o_1 \U$$4448  (.A1(net1054),
    .A2(\sel_0$6647 ),
    .B1(net1046),
    .B2(net696),
    .X(\t$6678 ));
 sky130_fd_sc_hd__xor2_1 \U$$4449  (.A(\t$6678 ),
    .B(net1845),
    .X(booth_b64_m29));
 sky130_fd_sc_hd__a22o_1 \U$$445  (.A1(net1198),
    .A2(net429),
    .B1(net1179),
    .B2(net711),
    .X(\t$4633 ));
 sky130_fd_sc_hd__a22o_1 \U$$4450  (.A1(net1046),
    .A2(\sel_0$6647 ),
    .B1(net1029),
    .B2(net698),
    .X(\t$6679 ));
 sky130_fd_sc_hd__xor2_1 \U$$4451  (.A(\t$6679 ),
    .B(net1846),
    .X(booth_b64_m30));
 sky130_fd_sc_hd__a22o_1 \U$$4452  (.A1(net1030),
    .A2(\sel_0$6647 ),
    .B1(net1022),
    .B2(net698),
    .X(\t$6680 ));
 sky130_fd_sc_hd__xor2_1 \U$$4453  (.A(\t$6680 ),
    .B(net1847),
    .X(booth_b64_m31));
 sky130_fd_sc_hd__a22o_1 \U$$4454  (.A1(net1022),
    .A2(\sel_0$6647 ),
    .B1(net1005),
    .B2(net699),
    .X(\t$6681 ));
 sky130_fd_sc_hd__xor2_1 \U$$4455  (.A(\t$6681 ),
    .B(net1848),
    .X(booth_b64_m32));
 sky130_fd_sc_hd__a22o_1 \U$$4456  (.A1(net1005),
    .A2(\sel_0$6647 ),
    .B1(net997),
    .B2(net697),
    .X(\t$6682 ));
 sky130_fd_sc_hd__xor2_1 \U$$4457  (.A(\t$6682 ),
    .B(net1849),
    .X(booth_b64_m33));
 sky130_fd_sc_hd__a22o_1 \U$$4458  (.A1(net997),
    .A2(\sel_0$6647 ),
    .B1(net989),
    .B2(net697),
    .X(\t$6683 ));
 sky130_fd_sc_hd__xor2_1 \U$$4459  (.A(\t$6683 ),
    .B(net1850),
    .X(booth_b64_m34));
 sky130_fd_sc_hd__xor2_1 \U$$446  (.A(\t$4633 ),
    .B(net1249),
    .X(booth_b6_m14));
 sky130_fd_sc_hd__a22o_1 \U$$4460  (.A1(net989),
    .A2(\sel_0$6647 ),
    .B1(net980),
    .B2(net697),
    .X(\t$6684 ));
 sky130_fd_sc_hd__xor2_1 \U$$4461  (.A(\t$6684 ),
    .B(net1851),
    .X(booth_b64_m35));
 sky130_fd_sc_hd__a22o_1 \U$$4462  (.A1(net980),
    .A2(\sel_0$6647 ),
    .B1(net971),
    .B2(net697),
    .X(\t$6685 ));
 sky130_fd_sc_hd__xor2_1 \U$$4463  (.A(\t$6685 ),
    .B(net1852),
    .X(booth_b64_m36));
 sky130_fd_sc_hd__a22o_1 \U$$4464  (.A1(net971),
    .A2(\sel_0$6647 ),
    .B1(net963),
    .B2(net699),
    .X(\t$6686 ));
 sky130_fd_sc_hd__xor2_1 \U$$4465  (.A(\t$6686 ),
    .B(net1853),
    .X(booth_b64_m37));
 sky130_fd_sc_hd__a22o_1 \U$$4466  (.A1(net963),
    .A2(\sel_0$6647 ),
    .B1(net953),
    .B2(net697),
    .X(\t$6687 ));
 sky130_fd_sc_hd__xor2_1 \U$$4467  (.A(\t$6687 ),
    .B(net1854),
    .X(booth_b64_m38));
 sky130_fd_sc_hd__a22o_1 \U$$4468  (.A1(net954),
    .A2(\sel_0$6647 ),
    .B1(net945),
    .B2(net699),
    .X(\t$6688 ));
 sky130_fd_sc_hd__xor2_1 \U$$4469  (.A(\t$6688 ),
    .B(net1855),
    .X(booth_b64_m39));
 sky130_fd_sc_hd__a22o_1 \U$$447  (.A1(net1180),
    .A2(net429),
    .B1(net1171),
    .B2(net711),
    .X(\t$4634 ));
 sky130_fd_sc_hd__a22o_1 \U$$4470  (.A1(net946),
    .A2(\sel_0$6647 ),
    .B1(net930),
    .B2(net697),
    .X(\t$6689 ));
 sky130_fd_sc_hd__xor2_1 \U$$4471  (.A(\t$6689 ),
    .B(net1856),
    .X(booth_b64_m40));
 sky130_fd_sc_hd__a22o_1 \U$$4472  (.A1(net930),
    .A2(\sel_0$6647 ),
    .B1(net1751),
    .B2(net697),
    .X(\t$6690 ));
 sky130_fd_sc_hd__xor2_1 \U$$4473  (.A(\t$6690 ),
    .B(net1857),
    .X(booth_b64_m41));
 sky130_fd_sc_hd__a22o_1 \U$$4474  (.A1(net1747),
    .A2(\sel_0$6647 ),
    .B1(net1739),
    .B2(net693),
    .X(\t$6691 ));
 sky130_fd_sc_hd__xor2_1 \U$$4475  (.A(\t$6691 ),
    .B(net1858),
    .X(booth_b64_m42));
 sky130_fd_sc_hd__a22o_1 \U$$4476  (.A1(net1743),
    .A2(\sel_0$6647 ),
    .B1(net1735),
    .B2(net696),
    .X(\t$6692 ));
 sky130_fd_sc_hd__xor2_1 \U$$4477  (.A(\t$6692 ),
    .B(net1859),
    .X(booth_b64_m43));
 sky130_fd_sc_hd__a22o_1 \U$$4478  (.A1(net1735),
    .A2(\sel_0$6647 ),
    .B1(net1727),
    .B2(net696),
    .X(\t$6693 ));
 sky130_fd_sc_hd__xor2_1 \U$$4479  (.A(\t$6693 ),
    .B(net1860),
    .X(booth_b64_m44));
 sky130_fd_sc_hd__xor2_1 \U$$448  (.A(\t$4634 ),
    .B(net1248),
    .X(booth_b6_m15));
 sky130_fd_sc_hd__a22o_1 \U$$4480  (.A1(net1727),
    .A2(\sel_0$6647 ),
    .B1(net1719),
    .B2(net696),
    .X(\t$6694 ));
 sky130_fd_sc_hd__xor2_1 \U$$4481  (.A(\t$6694 ),
    .B(net1861),
    .X(booth_b64_m45));
 sky130_fd_sc_hd__a22o_1 \U$$4482  (.A1(net1719),
    .A2(\sel_0$6647 ),
    .B1(net1710),
    .B2(net699),
    .X(\t$6695 ));
 sky130_fd_sc_hd__xor2_1 \U$$4483  (.A(\t$6695 ),
    .B(net1862),
    .X(booth_b64_m46));
 sky130_fd_sc_hd__a22o_1 \U$$4484  (.A1(net1710),
    .A2(\sel_0$6647 ),
    .B1(net1702),
    .B2(net696),
    .X(\t$6696 ));
 sky130_fd_sc_hd__xor2_1 \U$$4485  (.A(\t$6696 ),
    .B(net1863),
    .X(booth_b64_m47));
 sky130_fd_sc_hd__a22o_1 \U$$4486  (.A1(net1696),
    .A2(\sel_0$6647 ),
    .B1(net1688),
    .B2(net693),
    .X(\t$6697 ));
 sky130_fd_sc_hd__xor2_1 \U$$4487  (.A(\t$6697 ),
    .B(net1864),
    .X(booth_b64_m48));
 sky130_fd_sc_hd__a22o_1 \U$$4488  (.A1(net1694),
    .A2(\sel_0$6647 ),
    .B1(net1685),
    .B2(net696),
    .X(\t$6698 ));
 sky130_fd_sc_hd__xor2_1 \U$$4489  (.A(\t$6698 ),
    .B(net1865),
    .X(booth_b64_m49));
 sky130_fd_sc_hd__a22o_1 \U$$449  (.A1(net1170),
    .A2(net429),
    .B1(net1161),
    .B2(net711),
    .X(\t$4635 ));
 sky130_fd_sc_hd__a22o_1 \U$$4490  (.A1(net1685),
    .A2(\sel_0$6647 ),
    .B1(net1659),
    .B2(net697),
    .X(\t$6699 ));
 sky130_fd_sc_hd__xor2_1 \U$$4491  (.A(\t$6699 ),
    .B(net1866),
    .X(booth_b64_m50));
 sky130_fd_sc_hd__a22o_1 \U$$4492  (.A1(net1661),
    .A2(\sel_0$6647 ),
    .B1(net1653),
    .B2(net697),
    .X(\t$6700 ));
 sky130_fd_sc_hd__xor2_1 \U$$4493  (.A(\t$6700 ),
    .B(net1867),
    .X(booth_b64_m51));
 sky130_fd_sc_hd__a22o_1 \U$$4494  (.A1(net1653),
    .A2(\sel_0$6647 ),
    .B1(net1645),
    .B2(net697),
    .X(\t$6701 ));
 sky130_fd_sc_hd__xor2_1 \U$$4495  (.A(\t$6701 ),
    .B(net1868),
    .X(booth_b64_m52));
 sky130_fd_sc_hd__a22o_1 \U$$4496  (.A1(net1640),
    .A2(\sel_0$6647 ),
    .B1(net1632),
    .B2(net695),
    .X(\t$6702 ));
 sky130_fd_sc_hd__xor2_1 \U$$4497  (.A(\t$6702 ),
    .B(net1869),
    .X(booth_b64_m53));
 sky130_fd_sc_hd__a22o_1 \U$$4498  (.A1(net1636),
    .A2(\sel_0$6647 ),
    .B1(net1625),
    .B2(net696),
    .X(\t$6703 ));
 sky130_fd_sc_hd__xor2_1 \U$$4499  (.A(\t$6703 ),
    .B(net1870),
    .X(booth_b64_m54));
 sky130_fd_sc_hd__xor2_1 \U$$45  (.A(\t$4429 ),
    .B(net1575),
    .X(booth_b0_m19));
 sky130_fd_sc_hd__xor2_1 \U$$450  (.A(\t$4635 ),
    .B(net1249),
    .X(booth_b6_m16));
 sky130_fd_sc_hd__a22o_1 \U$$4500  (.A1(net1625),
    .A2(\sel_0$6647 ),
    .B1(net1617),
    .B2(net699),
    .X(\t$6704 ));
 sky130_fd_sc_hd__xor2_1 \U$$4501  (.A(\t$6704 ),
    .B(net1871),
    .X(booth_b64_m55));
 sky130_fd_sc_hd__a22o_1 \U$$4502  (.A1(net1614),
    .A2(\sel_0$6647 ),
    .B1(net1606),
    .B2(net699),
    .X(\t$6705 ));
 sky130_fd_sc_hd__xor2_1 \U$$4503  (.A(\t$6705 ),
    .B(net1872),
    .X(booth_b64_m56));
 sky130_fd_sc_hd__a22o_1 \U$$4504  (.A1(net1605),
    .A2(\sel_0$6647 ),
    .B1(net1597),
    .B2(net693),
    .X(\t$6706 ));
 sky130_fd_sc_hd__xor2_1 \U$$4505  (.A(\t$6706 ),
    .B(net1873),
    .X(booth_b64_m57));
 sky130_fd_sc_hd__a22o_1 \U$$4506  (.A1(net1601),
    .A2(\sel_0$6647 ),
    .B1(net1592),
    .B2(net696),
    .X(\t$6707 ));
 sky130_fd_sc_hd__xor2_1 \U$$4507  (.A(\t$6707 ),
    .B(net1874),
    .X(booth_b64_m58));
 sky130_fd_sc_hd__a22o_1 \U$$4508  (.A1(net1589),
    .A2(\sel_0$6647 ),
    .B1(net1580),
    .B2(net695),
    .X(\t$6708 ));
 sky130_fd_sc_hd__xor2_1 \U$$4509  (.A(\t$6708 ),
    .B(net1875),
    .X(booth_b64_m59));
 sky130_fd_sc_hd__a22o_1 \U$$451  (.A1(net1161),
    .A2(net431),
    .B1(net1149),
    .B2(net713),
    .X(\t$4636 ));
 sky130_fd_sc_hd__a22o_1 \U$$4510  (.A1(net1580),
    .A2(\sel_0$6647 ),
    .B1(net1554),
    .B2(net695),
    .X(\t$6709 ));
 sky130_fd_sc_hd__xor2_1 \U$$4511  (.A(\t$6709 ),
    .B(net1876),
    .X(booth_b64_m60));
 sky130_fd_sc_hd__a22o_1 \U$$4512  (.A1(net1553),
    .A2(\sel_0$6647 ),
    .B1(net1544),
    .B2(net693),
    .X(\t$6710 ));
 sky130_fd_sc_hd__xor2_1 \U$$4513  (.A(\t$6710 ),
    .B(net1877),
    .X(booth_b64_m61));
 sky130_fd_sc_hd__a22o_1 \U$$4514  (.A1(net1544),
    .A2(\sel_0$6647 ),
    .B1(net1536),
    .B2(net693),
    .X(\t$6711 ));
 sky130_fd_sc_hd__xor2_1 \U$$4515  (.A(\t$6711 ),
    .B(net1878),
    .X(booth_b64_m62));
 sky130_fd_sc_hd__a22o_1 \U$$4516  (.A1(net1536),
    .A2(\sel_0$6647 ),
    .B1(net1528),
    .B2(net693),
    .X(\t$6712 ));
 sky130_fd_sc_hd__xor2_1 \U$$4517  (.A(\t$6712 ),
    .B(net1879),
    .X(booth_b64_m63));
 sky130_fd_sc_hd__xor2_1 \U$$452  (.A(\t$4636 ),
    .B(net1250),
    .X(booth_b6_m17));
 sky130_fd_sc_hd__a22o_1 \U$$453  (.A1(net1147),
    .A2(net427),
    .B1(net1139),
    .B2(net709),
    .X(\t$4637 ));
 sky130_fd_sc_hd__xor2_1 \U$$454  (.A(\t$4637 ),
    .B(net1245),
    .X(booth_b6_m18));
 sky130_fd_sc_hd__a22o_1 \U$$455  (.A1(net1139),
    .A2(net427),
    .B1(net1131),
    .B2(net709),
    .X(\t$4638 ));
 sky130_fd_sc_hd__xor2_1 \U$$456  (.A(\t$4638 ),
    .B(net1245),
    .X(booth_b6_m19));
 sky130_fd_sc_hd__a22o_1 \U$$457  (.A1(net1130),
    .A2(net426),
    .B1(net1114),
    .B2(net708),
    .X(\t$4639 ));
 sky130_fd_sc_hd__xor2_1 \U$$458  (.A(\t$4639 ),
    .B(net1244),
    .X(booth_b6_m20));
 sky130_fd_sc_hd__a22o_1 \U$$459  (.A1(net1114),
    .A2(net426),
    .B1(net1105),
    .B2(net708),
    .X(\t$4640 ));
 sky130_fd_sc_hd__a22o_1 \U$$46  (.A1(net1133),
    .A2(net448),
    .B1(net1117),
    .B2(net690),
    .X(\t$4430 ));
 sky130_fd_sc_hd__xor2_1 \U$$460  (.A(\t$4640 ),
    .B(net1244),
    .X(booth_b6_m21));
 sky130_fd_sc_hd__a22o_1 \U$$461  (.A1(net1105),
    .A2(net426),
    .B1(net1097),
    .B2(net708),
    .X(\t$4641 ));
 sky130_fd_sc_hd__xor2_1 \U$$462  (.A(\t$4641 ),
    .B(net1244),
    .X(booth_b6_m22));
 sky130_fd_sc_hd__a22o_1 \U$$463  (.A1(net1097),
    .A2(net426),
    .B1(net1088),
    .B2(net708),
    .X(\t$4642 ));
 sky130_fd_sc_hd__xor2_1 \U$$464  (.A(\t$4642 ),
    .B(net1244),
    .X(booth_b6_m23));
 sky130_fd_sc_hd__a22o_1 \U$$465  (.A1(net1088),
    .A2(net426),
    .B1(net1080),
    .B2(net708),
    .X(\t$4643 ));
 sky130_fd_sc_hd__xor2_1 \U$$466  (.A(\t$4643 ),
    .B(net1244),
    .X(booth_b6_m24));
 sky130_fd_sc_hd__a22o_1 \U$$467  (.A1(net1080),
    .A2(net428),
    .B1(net1071),
    .B2(net710),
    .X(\t$4644 ));
 sky130_fd_sc_hd__xor2_1 \U$$468  (.A(\t$4644 ),
    .B(net1245),
    .X(booth_b6_m25));
 sky130_fd_sc_hd__a22o_1 \U$$469  (.A1(net1072),
    .A2(net427),
    .B1(net1064),
    .B2(net709),
    .X(\t$4645 ));
 sky130_fd_sc_hd__xor2_1 \U$$47  (.A(\t$4430 ),
    .B(net1575),
    .X(booth_b0_m20));
 sky130_fd_sc_hd__xor2_1 \U$$470  (.A(\t$4645 ),
    .B(net1245),
    .X(booth_b6_m26));
 sky130_fd_sc_hd__a22o_1 \U$$471  (.A1(net1066),
    .A2(net429),
    .B1(net1057),
    .B2(net711),
    .X(\t$4646 ));
 sky130_fd_sc_hd__xor2_1 \U$$472  (.A(\t$4646 ),
    .B(net1249),
    .X(booth_b6_m27));
 sky130_fd_sc_hd__a22o_1 \U$$473  (.A1(net1058),
    .A2(net429),
    .B1(net1050),
    .B2(net711),
    .X(\t$4647 ));
 sky130_fd_sc_hd__xor2_1 \U$$474  (.A(\t$4647 ),
    .B(net1248),
    .X(booth_b6_m28));
 sky130_fd_sc_hd__a22o_1 \U$$475  (.A1(net1050),
    .A2(net429),
    .B1(net1042),
    .B2(net711),
    .X(\t$4648 ));
 sky130_fd_sc_hd__xor2_1 \U$$476  (.A(\t$4648 ),
    .B(net1249),
    .X(booth_b6_m29));
 sky130_fd_sc_hd__a22o_1 \U$$477  (.A1(net1041),
    .A2(net431),
    .B1(net1025),
    .B2(net713),
    .X(\t$4649 ));
 sky130_fd_sc_hd__xor2_1 \U$$478  (.A(\t$4649 ),
    .B(net1250),
    .X(booth_b6_m30));
 sky130_fd_sc_hd__a22o_1 \U$$479  (.A1(net1025),
    .A2(net431),
    .B1(net1017),
    .B2(net713),
    .X(\t$4650 ));
 sky130_fd_sc_hd__a22o_1 \U$$48  (.A1(net1117),
    .A2(net448),
    .B1(net1108),
    .B2(net690),
    .X(\t$4431 ));
 sky130_fd_sc_hd__xor2_1 \U$$480  (.A(\t$4650 ),
    .B(net1250),
    .X(booth_b6_m31));
 sky130_fd_sc_hd__a22o_1 \U$$481  (.A1(net1016),
    .A2(net427),
    .B1(net998),
    .B2(net709),
    .X(\t$4651 ));
 sky130_fd_sc_hd__xor2_1 \U$$482  (.A(\t$4651 ),
    .B(net1245),
    .X(booth_b6_m32));
 sky130_fd_sc_hd__a22o_1 \U$$483  (.A1(net1000),
    .A2(net431),
    .B1(net992),
    .B2(net713),
    .X(\t$4652 ));
 sky130_fd_sc_hd__xor2_1 \U$$484  (.A(\t$4652 ),
    .B(net1250),
    .X(booth_b6_m33));
 sky130_fd_sc_hd__a22o_1 \U$$485  (.A1(net990),
    .A2(net428),
    .B1(net986),
    .B2(net710),
    .X(\t$4653 ));
 sky130_fd_sc_hd__xor2_1 \U$$486  (.A(\t$4653 ),
    .B(net1245),
    .X(booth_b6_m34));
 sky130_fd_sc_hd__a22o_1 \U$$487  (.A1(net982),
    .A2(net426),
    .B1(net973),
    .B2(net708),
    .X(\t$4654 ));
 sky130_fd_sc_hd__xor2_1 \U$$488  (.A(\t$4654 ),
    .B(net1244),
    .X(booth_b6_m35));
 sky130_fd_sc_hd__a22o_1 \U$$489  (.A1(net973),
    .A2(net426),
    .B1(net964),
    .B2(net708),
    .X(\t$4655 ));
 sky130_fd_sc_hd__xor2_1 \U$$49  (.A(\t$4431 ),
    .B(net1575),
    .X(booth_b0_m21));
 sky130_fd_sc_hd__xor2_1 \U$$490  (.A(\t$4655 ),
    .B(net1244),
    .X(booth_b6_m36));
 sky130_fd_sc_hd__a22o_1 \U$$491  (.A1(net964),
    .A2(net426),
    .B1(net956),
    .B2(net708),
    .X(\t$4656 ));
 sky130_fd_sc_hd__xor2_1 \U$$492  (.A(\t$4656 ),
    .B(net1244),
    .X(booth_b6_m37));
 sky130_fd_sc_hd__a22o_1 \U$$493  (.A1(net956),
    .A2(net427),
    .B1(net948),
    .B2(net709),
    .X(\t$4657 ));
 sky130_fd_sc_hd__xor2_1 \U$$494  (.A(\t$4657 ),
    .B(net1253),
    .X(booth_b6_m38));
 sky130_fd_sc_hd__a22o_1 \U$$495  (.A1(net949),
    .A2(net427),
    .B1(net941),
    .B2(net709),
    .X(\t$4658 ));
 sky130_fd_sc_hd__xor2_1 \U$$496  (.A(\t$4658 ),
    .B(net1253),
    .X(booth_b6_m39));
 sky130_fd_sc_hd__a22o_1 \U$$497  (.A1(net940),
    .A2(net427),
    .B1(net924),
    .B2(net709),
    .X(\t$4659 ));
 sky130_fd_sc_hd__xor2_1 \U$$498  (.A(\t$4659 ),
    .B(net1244),
    .X(booth_b6_m40));
 sky130_fd_sc_hd__a22o_1 \U$$499  (.A1(net924),
    .A2(net426),
    .B1(net1745),
    .B2(net708),
    .X(\t$4660 ));
 sky130_fd_sc_hd__xor2_1 \U$$5  (.A(net1),
    .B(net1880),
    .X(sel_1));
 sky130_fd_sc_hd__a22o_1 \U$$50  (.A1(net1108),
    .A2(net448),
    .B1(net1100),
    .B2(net690),
    .X(\t$4432 ));
 sky130_fd_sc_hd__xor2_1 \U$$500  (.A(\t$4660 ),
    .B(net1244),
    .X(booth_b6_m41));
 sky130_fd_sc_hd__a22o_1 \U$$501  (.A1(net1745),
    .A2(net426),
    .B1(net1737),
    .B2(net708),
    .X(\t$4661 ));
 sky130_fd_sc_hd__xor2_1 \U$$502  (.A(\t$4661 ),
    .B(net1245),
    .X(booth_b6_m42));
 sky130_fd_sc_hd__a22o_1 \U$$503  (.A1(net1738),
    .A2(net428),
    .B1(net1730),
    .B2(net710),
    .X(\t$4662 ));
 sky130_fd_sc_hd__xor2_1 \U$$504  (.A(\t$4662 ),
    .B(net1247),
    .X(booth_b6_m43));
 sky130_fd_sc_hd__a22o_1 \U$$505  (.A1(net1729),
    .A2(net428),
    .B1(net1720),
    .B2(net710),
    .X(\t$4663 ));
 sky130_fd_sc_hd__xor2_1 \U$$506  (.A(\t$4663 ),
    .B(net1246),
    .X(booth_b6_m44));
 sky130_fd_sc_hd__a22o_1 \U$$507  (.A1(net1725),
    .A2(net432),
    .B1(net1716),
    .B2(net714),
    .X(\t$4664 ));
 sky130_fd_sc_hd__xor2_1 \U$$508  (.A(\t$4664 ),
    .B(net1251),
    .X(booth_b6_m45));
 sky130_fd_sc_hd__a22o_1 \U$$509  (.A1(net1716),
    .A2(net430),
    .B1(net1707),
    .B2(net712),
    .X(\t$4665 ));
 sky130_fd_sc_hd__xor2_1 \U$$51  (.A(\t$4432 ),
    .B(net1575),
    .X(booth_b0_m22));
 sky130_fd_sc_hd__xor2_1 \U$$510  (.A(\t$4665 ),
    .B(net1252),
    .X(booth_b6_m46));
 sky130_fd_sc_hd__a22o_1 \U$$511  (.A1(net1707),
    .A2(net430),
    .B1(net1699),
    .B2(net712),
    .X(\t$4666 ));
 sky130_fd_sc_hd__xor2_1 \U$$512  (.A(\t$4666 ),
    .B(net1250),
    .X(booth_b6_m47));
 sky130_fd_sc_hd__a22o_1 \U$$513  (.A1(net1699),
    .A2(net430),
    .B1(net1691),
    .B2(net712),
    .X(\t$4667 ));
 sky130_fd_sc_hd__xor2_1 \U$$514  (.A(\t$4667 ),
    .B(net1250),
    .X(booth_b6_m48));
 sky130_fd_sc_hd__a22o_1 \U$$515  (.A1(net1691),
    .A2(net432),
    .B1(net1683),
    .B2(net714),
    .X(\t$4668 ));
 sky130_fd_sc_hd__xor2_1 \U$$516  (.A(\t$4668 ),
    .B(net1251),
    .X(booth_b6_m49));
 sky130_fd_sc_hd__a22o_1 \U$$517  (.A1(net1682),
    .A2(net432),
    .B1(net1657),
    .B2(net714),
    .X(\t$4669 ));
 sky130_fd_sc_hd__xor2_1 \U$$518  (.A(\t$4669 ),
    .B(net1251),
    .X(booth_b6_m50));
 sky130_fd_sc_hd__a22o_1 \U$$519  (.A1(net1657),
    .A2(net433),
    .B1(net1649),
    .B2(net715),
    .X(\t$4670 ));
 sky130_fd_sc_hd__a22o_1 \U$$52  (.A1(net1100),
    .A2(net448),
    .B1(net1091),
    .B2(net690),
    .X(\t$4433 ));
 sky130_fd_sc_hd__xor2_1 \U$$520  (.A(\t$4670 ),
    .B(net1251),
    .X(booth_b6_m51));
 sky130_fd_sc_hd__a22o_1 \U$$521  (.A1(net1649),
    .A2(net432),
    .B1(net1641),
    .B2(net714),
    .X(\t$4671 ));
 sky130_fd_sc_hd__xor2_1 \U$$522  (.A(\t$4671 ),
    .B(net1251),
    .X(booth_b6_m52));
 sky130_fd_sc_hd__a22o_1 \U$$523  (.A1(net1638),
    .A2(net428),
    .B1(net1629),
    .B2(net710),
    .X(\t$4672 ));
 sky130_fd_sc_hd__xor2_1 \U$$524  (.A(\t$4672 ),
    .B(net1247),
    .X(booth_b6_m53));
 sky130_fd_sc_hd__a22o_1 \U$$525  (.A1(net1630),
    .A2(net428),
    .B1(net1621),
    .B2(net710),
    .X(\t$4673 ));
 sky130_fd_sc_hd__xor2_1 \U$$526  (.A(\t$4673 ),
    .B(net1247),
    .X(booth_b6_m54));
 sky130_fd_sc_hd__a22o_1 \U$$527  (.A1(net1620),
    .A2(net428),
    .B1(net1612),
    .B2(net710),
    .X(\t$4674 ));
 sky130_fd_sc_hd__xor2_1 \U$$528  (.A(\t$4674 ),
    .B(net1246),
    .X(booth_b6_m55));
 sky130_fd_sc_hd__a22o_1 \U$$529  (.A1(net1612),
    .A2(net428),
    .B1(net1604),
    .B2(net710),
    .X(\t$4675 ));
 sky130_fd_sc_hd__xor2_1 \U$$53  (.A(\t$4433 ),
    .B(net1575),
    .X(booth_b0_m23));
 sky130_fd_sc_hd__xor2_1 \U$$530  (.A(\t$4675 ),
    .B(net1246),
    .X(booth_b6_m56));
 sky130_fd_sc_hd__a22o_1 \U$$531  (.A1(net1604),
    .A2(net433),
    .B1(net1595),
    .B2(net715),
    .X(\t$4676 ));
 sky130_fd_sc_hd__xor2_1 \U$$532  (.A(\t$4676 ),
    .B(net1246),
    .X(booth_b6_m57));
 sky130_fd_sc_hd__a22o_1 \U$$533  (.A1(net1595),
    .A2(net428),
    .B1(net1586),
    .B2(net710),
    .X(\t$4677 ));
 sky130_fd_sc_hd__xor2_1 \U$$534  (.A(\t$4677 ),
    .B(net1246),
    .X(booth_b6_m58));
 sky130_fd_sc_hd__a22o_1 \U$$535  (.A1(net1590),
    .A2(net432),
    .B1(net1582),
    .B2(net714),
    .X(\t$4678 ));
 sky130_fd_sc_hd__xor2_1 \U$$536  (.A(\t$4678 ),
    .B(net1251),
    .X(booth_b6_m59));
 sky130_fd_sc_hd__a22o_1 \U$$537  (.A1(net1582),
    .A2(net432),
    .B1(net1555),
    .B2(net714),
    .X(\t$4679 ));
 sky130_fd_sc_hd__xor2_1 \U$$538  (.A(\t$4679 ),
    .B(net1251),
    .X(booth_b6_m60));
 sky130_fd_sc_hd__a22o_1 \U$$539  (.A1(net1559),
    .A2(net432),
    .B1(net122),
    .B2(net714),
    .X(\t$4680 ));
 sky130_fd_sc_hd__a22o_1 \U$$54  (.A1(net1089),
    .A2(net443),
    .B1(net1081),
    .B2(net685),
    .X(\t$4434 ));
 sky130_fd_sc_hd__xor2_1 \U$$540  (.A(\t$4680 ),
    .B(net1252),
    .X(booth_b6_m61));
 sky130_fd_sc_hd__a22o_1 \U$$541  (.A1(net1547),
    .A2(net432),
    .B1(net1539),
    .B2(net714),
    .X(\t$4681 ));
 sky130_fd_sc_hd__xor2_1 \U$$542  (.A(\t$4681 ),
    .B(net1251),
    .X(booth_b6_m62));
 sky130_fd_sc_hd__a22o_1 \U$$543  (.A1(net1539),
    .A2(net432),
    .B1(net1531),
    .B2(net714),
    .X(\t$4682 ));
 sky130_fd_sc_hd__xor2_1 \U$$544  (.A(\t$4682 ),
    .B(net1251),
    .X(booth_b6_m63));
 sky130_fd_sc_hd__a22o_1 \U$$545  (.A1(net1531),
    .A2(net432),
    .B1(net1881),
    .B2(net714),
    .X(\t$4683 ));
 sky130_fd_sc_hd__xor2_1 \U$$546  (.A(\t$4683 ),
    .B(net1251),
    .X(booth_b6_m64));
 sky130_fd_sc_hd__inv_1 \U$$547  (.A(net1246),
    .Y(\notsign$4684 ));
 sky130_fd_sc_hd__inv_1 \U$$548  (.A(net1246),
    .Y(\notblock$4685[0] ));
 sky130_fd_sc_hd__inv_1 \U$$549  (.A(net63),
    .Y(\notblock$4685[1] ));
 sky130_fd_sc_hd__xor2_1 \U$$55  (.A(\t$4434 ),
    .B(net1569),
    .X(booth_b0_m24));
 sky130_fd_sc_hd__inv_1 \U$$550  (.A(net1237),
    .Y(\notblock$4685[2] ));
 sky130_fd_sc_hd__and2_1 \U$$551  (.A(net1237),
    .B(\notblock$4685[1] ),
    .X(\t$4686 ));
 sky130_fd_sc_hd__a32o_1 \U$$552  (.A1(\notblock$4685[2] ),
    .A2(net63),
    .A3(net1246),
    .B1(\t$4686 ),
    .B2(\notblock$4685[0] ),
    .X(\sel_0$4687 ));
 sky130_fd_sc_hd__xor2_1 \U$$553  (.A(net63),
    .B(net1247),
    .X(\sel_1$4688 ));
 sky130_fd_sc_hd__a22o_1 \U$$554  (.A1(net1882),
    .A2(net413),
    .B1(net1231),
    .B2(net679),
    .X(\t$4689 ));
 sky130_fd_sc_hd__xor2_1 \U$$555  (.A(\t$4689 ),
    .B(net1239),
    .X(booth_b8_m0));
 sky130_fd_sc_hd__a22o_1 \U$$556  (.A1(net1231),
    .A2(net413),
    .B1(net1127),
    .B2(net679),
    .X(\t$4690 ));
 sky130_fd_sc_hd__xor2_1 \U$$557  (.A(\t$4690 ),
    .B(net1239),
    .X(booth_b8_m1));
 sky130_fd_sc_hd__a22o_1 \U$$558  (.A1(net1126),
    .A2(net414),
    .B1(net1036),
    .B2(net680),
    .X(\t$4691 ));
 sky130_fd_sc_hd__xor2_1 \U$$559  (.A(\t$4691 ),
    .B(net1239),
    .X(booth_b8_m2));
 sky130_fd_sc_hd__a22o_1 \U$$56  (.A1(net1080),
    .A2(net443),
    .B1(net1071),
    .B2(net685),
    .X(\t$4435 ));
 sky130_fd_sc_hd__a22o_1 \U$$560  (.A1(net1036),
    .A2(net414),
    .B1(net936),
    .B2(net680),
    .X(\t$4692 ));
 sky130_fd_sc_hd__xor2_1 \U$$561  (.A(\t$4692 ),
    .B(net1239),
    .X(booth_b8_m3));
 sky130_fd_sc_hd__a22o_1 \U$$562  (.A1(net937),
    .A2(net414),
    .B1(net1675),
    .B2(net680),
    .X(\t$4693 ));
 sky130_fd_sc_hd__xor2_1 \U$$563  (.A(\t$4693 ),
    .B(net1240),
    .X(booth_b8_m4));
 sky130_fd_sc_hd__a22o_1 \U$$564  (.A1(net1676),
    .A2(net414),
    .B1(net1564),
    .B2(net680),
    .X(\t$4694 ));
 sky130_fd_sc_hd__xor2_1 \U$$565  (.A(\t$4694 ),
    .B(net1240),
    .X(booth_b8_m5));
 sky130_fd_sc_hd__a22o_1 \U$$566  (.A1(net1561),
    .A2(net415),
    .B1(net1521),
    .B2(net681),
    .X(\t$4695 ));
 sky130_fd_sc_hd__xor2_1 \U$$567  (.A(\t$4695 ),
    .B(net1241),
    .X(booth_b8_m6));
 sky130_fd_sc_hd__a22o_1 \U$$568  (.A1(net1521),
    .A2(net415),
    .B1(net1513),
    .B2(net681),
    .X(\t$4696 ));
 sky130_fd_sc_hd__xor2_1 \U$$569  (.A(\t$4696 ),
    .B(net1241),
    .X(booth_b8_m7));
 sky130_fd_sc_hd__xor2_1 \U$$57  (.A(\t$4435 ),
    .B(net1569),
    .X(booth_b0_m25));
 sky130_fd_sc_hd__a22o_1 \U$$570  (.A1(net1513),
    .A2(net410),
    .B1(net1505),
    .B2(net676),
    .X(\t$4697 ));
 sky130_fd_sc_hd__xor2_1 \U$$571  (.A(\t$4697 ),
    .B(net1236),
    .X(booth_b8_m8));
 sky130_fd_sc_hd__a22o_1 \U$$572  (.A1(net1505),
    .A2(net410),
    .B1(net1496),
    .B2(net676),
    .X(\t$4698 ));
 sky130_fd_sc_hd__xor2_1 \U$$573  (.A(\t$4698 ),
    .B(net1236),
    .X(booth_b8_m9));
 sky130_fd_sc_hd__a22o_1 \U$$574  (.A1(net1496),
    .A2(net415),
    .B1(net1221),
    .B2(net681),
    .X(\t$4699 ));
 sky130_fd_sc_hd__xor2_1 \U$$575  (.A(\t$4699 ),
    .B(net1241),
    .X(booth_b8_m10));
 sky130_fd_sc_hd__a22o_1 \U$$576  (.A1(net1224),
    .A2(net413),
    .B1(net1216),
    .B2(net679),
    .X(\t$4700 ));
 sky130_fd_sc_hd__xor2_1 \U$$577  (.A(\t$4700 ),
    .B(net1239),
    .X(booth_b8_m11));
 sky130_fd_sc_hd__a22o_1 \U$$578  (.A1(net1216),
    .A2(net413),
    .B1(net1206),
    .B2(net679),
    .X(\t$4701 ));
 sky130_fd_sc_hd__xor2_1 \U$$579  (.A(\t$4701 ),
    .B(net1239),
    .X(booth_b8_m12));
 sky130_fd_sc_hd__a22o_1 \U$$58  (.A1(net1071),
    .A2(net442),
    .B1(net1063),
    .B2(net684),
    .X(\t$4436 ));
 sky130_fd_sc_hd__a22o_1 \U$$580  (.A1(net1207),
    .A2(net413),
    .B1(net1199),
    .B2(net679),
    .X(\t$4702 ));
 sky130_fd_sc_hd__xor2_1 \U$$581  (.A(\t$4702 ),
    .B(net1240),
    .X(booth_b8_m13));
 sky130_fd_sc_hd__a22o_1 \U$$582  (.A1(net1198),
    .A2(net413),
    .B1(net1179),
    .B2(net679),
    .X(\t$4703 ));
 sky130_fd_sc_hd__xor2_1 \U$$583  (.A(\t$4703 ),
    .B(net1239),
    .X(booth_b8_m14));
 sky130_fd_sc_hd__a22o_1 \U$$584  (.A1(net1179),
    .A2(net415),
    .B1(net1170),
    .B2(net681),
    .X(\t$4704 ));
 sky130_fd_sc_hd__xor2_1 \U$$585  (.A(\t$4704 ),
    .B(net1241),
    .X(booth_b8_m15));
 sky130_fd_sc_hd__a22o_1 \U$$586  (.A1(net1166),
    .A2(net409),
    .B1(net1157),
    .B2(net675),
    .X(\t$4705 ));
 sky130_fd_sc_hd__xor2_1 \U$$587  (.A(\t$4705 ),
    .B(net1241),
    .X(booth_b8_m16));
 sky130_fd_sc_hd__a22o_1 \U$$588  (.A1(net1155),
    .A2(net410),
    .B1(net1146),
    .B2(net676),
    .X(\t$4706 ));
 sky130_fd_sc_hd__xor2_1 \U$$589  (.A(\t$4706 ),
    .B(net1236),
    .X(booth_b8_m17));
 sky130_fd_sc_hd__xor2_1 \U$$59  (.A(\t$4436 ),
    .B(net1568),
    .X(booth_b0_m26));
 sky130_fd_sc_hd__a22o_1 \U$$590  (.A1(net1146),
    .A2(net409),
    .B1(net1138),
    .B2(net675),
    .X(\t$4707 ));
 sky130_fd_sc_hd__xor2_1 \U$$591  (.A(\t$4707 ),
    .B(net1235),
    .X(booth_b8_m18));
 sky130_fd_sc_hd__a22o_1 \U$$592  (.A1(net1138),
    .A2(net409),
    .B1(net1130),
    .B2(net675),
    .X(\t$4708 ));
 sky130_fd_sc_hd__xor2_1 \U$$593  (.A(\t$4708 ),
    .B(net1235),
    .X(booth_b8_m19));
 sky130_fd_sc_hd__a22o_1 \U$$594  (.A1(net1130),
    .A2(net409),
    .B1(net1114),
    .B2(net675),
    .X(\t$4709 ));
 sky130_fd_sc_hd__xor2_1 \U$$595  (.A(\t$4709 ),
    .B(net1235),
    .X(booth_b8_m20));
 sky130_fd_sc_hd__a22o_1 \U$$596  (.A1(net1114),
    .A2(net409),
    .B1(net1105),
    .B2(net675),
    .X(\t$4710 ));
 sky130_fd_sc_hd__xor2_1 \U$$597  (.A(\t$4710 ),
    .B(net1235),
    .X(booth_b8_m21));
 sky130_fd_sc_hd__a22o_1 \U$$598  (.A1(net1105),
    .A2(net409),
    .B1(net1097),
    .B2(net675),
    .X(\t$4711 ));
 sky130_fd_sc_hd__xor2_1 \U$$599  (.A(\t$4711 ),
    .B(net1235),
    .X(booth_b8_m22));
 sky130_fd_sc_hd__a22o_1 \U$$6  (.A1(net1883),
    .A2(net446),
    .B1(net1232),
    .B2(net688),
    .X(\t$4410 ));
 sky130_fd_sc_hd__a22o_1 \U$$60  (.A1(net1063),
    .A2(net442),
    .B1(net1055),
    .B2(net684),
    .X(\t$4437 ));
 sky130_fd_sc_hd__a22o_1 \U$$600  (.A1(net1097),
    .A2(net410),
    .B1(net1088),
    .B2(net676),
    .X(\t$4712 ));
 sky130_fd_sc_hd__xor2_1 \U$$601  (.A(\t$4712 ),
    .B(net1236),
    .X(booth_b8_m23));
 sky130_fd_sc_hd__a22o_1 \U$$602  (.A1(net1089),
    .A2(net410),
    .B1(net1081),
    .B2(net676),
    .X(\t$4713 ));
 sky130_fd_sc_hd__xor2_1 \U$$603  (.A(\t$4713 ),
    .B(net1236),
    .X(booth_b8_m24));
 sky130_fd_sc_hd__a22o_1 \U$$604  (.A1(net1083),
    .A2(net413),
    .B1(net1074),
    .B2(net679),
    .X(\t$4714 ));
 sky130_fd_sc_hd__xor2_1 \U$$605  (.A(\t$4714 ),
    .B(net1239),
    .X(booth_b8_m25));
 sky130_fd_sc_hd__a22o_1 \U$$606  (.A1(net1075),
    .A2(net413),
    .B1(net1067),
    .B2(net679),
    .X(\t$4715 ));
 sky130_fd_sc_hd__xor2_1 \U$$607  (.A(\t$4715 ),
    .B(net1240),
    .X(booth_b8_m26));
 sky130_fd_sc_hd__a22o_1 \U$$608  (.A1(net1066),
    .A2(net413),
    .B1(net1058),
    .B2(net679),
    .X(\t$4716 ));
 sky130_fd_sc_hd__xor2_1 \U$$609  (.A(\t$4716 ),
    .B(net1239),
    .X(booth_b8_m27));
 sky130_fd_sc_hd__xor2_1 \U$$61  (.A(\t$4437 ),
    .B(net1568),
    .X(booth_b0_m27));
 sky130_fd_sc_hd__a22o_1 \U$$610  (.A1(net1057),
    .A2(net413),
    .B1(net1049),
    .B2(net679),
    .X(\t$4717 ));
 sky130_fd_sc_hd__xor2_1 \U$$611  (.A(\t$4717 ),
    .B(net1239),
    .X(booth_b8_m28));
 sky130_fd_sc_hd__a22o_1 \U$$612  (.A1(net1049),
    .A2(net415),
    .B1(net1041),
    .B2(net681),
    .X(\t$4718 ));
 sky130_fd_sc_hd__xor2_1 \U$$613  (.A(\t$4718 ),
    .B(net1241),
    .X(booth_b8_m29));
 sky130_fd_sc_hd__a22o_1 \U$$614  (.A1(net1040),
    .A2(net410),
    .B1(net1024),
    .B2(net676),
    .X(\t$4719 ));
 sky130_fd_sc_hd__xor2_1 \U$$615  (.A(\t$4719 ),
    .B(net1236),
    .X(booth_b8_m30));
 sky130_fd_sc_hd__a22o_1 \U$$616  (.A1(net1025),
    .A2(net415),
    .B1(net1017),
    .B2(net681),
    .X(\t$4720 ));
 sky130_fd_sc_hd__xor2_1 \U$$617  (.A(\t$4720 ),
    .B(net1241),
    .X(booth_b8_m31));
 sky130_fd_sc_hd__a22o_1 \U$$618  (.A1(net1016),
    .A2(net410),
    .B1(net998),
    .B2(net676),
    .X(\t$4721 ));
 sky130_fd_sc_hd__xor2_1 \U$$619  (.A(\t$4721 ),
    .B(net1236),
    .X(booth_b8_m32));
 sky130_fd_sc_hd__a22o_1 \U$$62  (.A1(net1055),
    .A2(net442),
    .B1(net1047),
    .B2(net684),
    .X(\t$4438 ));
 sky130_fd_sc_hd__a22o_1 \U$$620  (.A1(net998),
    .A2(net409),
    .B1(net990),
    .B2(net675),
    .X(\t$4722 ));
 sky130_fd_sc_hd__xor2_1 \U$$621  (.A(\t$4722 ),
    .B(net1235),
    .X(booth_b8_m33));
 sky130_fd_sc_hd__a22o_1 \U$$622  (.A1(net990),
    .A2(net409),
    .B1(net982),
    .B2(net675),
    .X(\t$4723 ));
 sky130_fd_sc_hd__xor2_1 \U$$623  (.A(\t$4723 ),
    .B(net1235),
    .X(booth_b8_m34));
 sky130_fd_sc_hd__a22o_1 \U$$624  (.A1(net982),
    .A2(net409),
    .B1(net973),
    .B2(net675),
    .X(\t$4724 ));
 sky130_fd_sc_hd__xor2_1 \U$$625  (.A(\t$4724 ),
    .B(net1235),
    .X(booth_b8_m35));
 sky130_fd_sc_hd__a22o_1 \U$$626  (.A1(net973),
    .A2(net410),
    .B1(net964),
    .B2(net676),
    .X(\t$4725 ));
 sky130_fd_sc_hd__xor2_1 \U$$627  (.A(\t$4725 ),
    .B(net1236),
    .X(booth_b8_m36));
 sky130_fd_sc_hd__a22o_1 \U$$628  (.A1(net968),
    .A2(net415),
    .B1(net960),
    .B2(net681),
    .X(\t$4726 ));
 sky130_fd_sc_hd__xor2_1 \U$$629  (.A(\t$4726 ),
    .B(net1241),
    .X(booth_b8_m37));
 sky130_fd_sc_hd__xor2_1 \U$$63  (.A(\t$4438 ),
    .B(net1568),
    .X(booth_b0_m28));
 sky130_fd_sc_hd__a22o_1 \U$$630  (.A1(net956),
    .A2(net409),
    .B1(net948),
    .B2(net675),
    .X(\t$4727 ));
 sky130_fd_sc_hd__xor2_1 \U$$631  (.A(\t$4727 ),
    .B(net1235),
    .X(booth_b8_m38));
 sky130_fd_sc_hd__a22o_1 \U$$632  (.A1(net948),
    .A2(net411),
    .B1(net940),
    .B2(net677),
    .X(\t$4728 ));
 sky130_fd_sc_hd__xor2_1 \U$$633  (.A(\t$4728 ),
    .B(net1235),
    .X(booth_b8_m39));
 sky130_fd_sc_hd__a22o_1 \U$$634  (.A1(net940),
    .A2(net411),
    .B1(net924),
    .B2(net677),
    .X(\t$4729 ));
 sky130_fd_sc_hd__xor2_1 \U$$635  (.A(\t$4729 ),
    .B(net1237),
    .X(booth_b8_m40));
 sky130_fd_sc_hd__a22o_1 \U$$636  (.A1(net925),
    .A2(net412),
    .B1(net1746),
    .B2(net678),
    .X(\t$4730 ));
 sky130_fd_sc_hd__xor2_1 \U$$637  (.A(\t$4730 ),
    .B(net1238),
    .X(booth_b8_m41));
 sky130_fd_sc_hd__a22o_1 \U$$638  (.A1(net1745),
    .A2(net411),
    .B1(net1737),
    .B2(net677),
    .X(\t$4731 ));
 sky130_fd_sc_hd__xor2_1 \U$$639  (.A(\t$4731 ),
    .B(net1237),
    .X(booth_b8_m42));
 sky130_fd_sc_hd__a22o_1 \U$$64  (.A1(net1047),
    .A2(net442),
    .B1(net1039),
    .B2(net684),
    .X(\t$4439 ));
 sky130_fd_sc_hd__a22o_1 \U$$640  (.A1(net1744),
    .A2(net416),
    .B1(net1736),
    .B2(net682),
    .X(\t$4732 ));
 sky130_fd_sc_hd__xor2_1 \U$$641  (.A(\t$4732 ),
    .B(net1242),
    .X(booth_b8_m43));
 sky130_fd_sc_hd__a22o_1 \U$$642  (.A1(net1736),
    .A2(net414),
    .B1(net1725),
    .B2(net680),
    .X(\t$4733 ));
 sky130_fd_sc_hd__xor2_1 \U$$643  (.A(\t$4733 ),
    .B(net1241),
    .X(booth_b8_m44));
 sky130_fd_sc_hd__a22o_1 \U$$644  (.A1(net1725),
    .A2(net417),
    .B1(net1716),
    .B2(net683),
    .X(\t$4734 ));
 sky130_fd_sc_hd__xor2_1 \U$$645  (.A(\t$4734 ),
    .B(net1242),
    .X(booth_b8_m45));
 sky130_fd_sc_hd__a22o_1 \U$$646  (.A1(net1716),
    .A2(net414),
    .B1(net1707),
    .B2(net680),
    .X(\t$4735 ));
 sky130_fd_sc_hd__xor2_1 \U$$647  (.A(\t$4735 ),
    .B(net1241),
    .X(booth_b8_m46));
 sky130_fd_sc_hd__a22o_1 \U$$648  (.A1(net1707),
    .A2(net416),
    .B1(net1699),
    .B2(net682),
    .X(\t$4736 ));
 sky130_fd_sc_hd__xor2_1 \U$$649  (.A(\t$4736 ),
    .B(net1242),
    .X(booth_b8_m47));
 sky130_fd_sc_hd__xor2_1 \U$$65  (.A(\t$4439 ),
    .B(net1568),
    .X(booth_b0_m29));
 sky130_fd_sc_hd__a22o_1 \U$$650  (.A1(net1698),
    .A2(net416),
    .B1(net1690),
    .B2(net682),
    .X(\t$4737 ));
 sky130_fd_sc_hd__xor2_1 \U$$651  (.A(\t$4737 ),
    .B(net1242),
    .X(booth_b8_m48));
 sky130_fd_sc_hd__a22o_1 \U$$652  (.A1(net1690),
    .A2(net416),
    .B1(net1682),
    .B2(net682),
    .X(\t$4738 ));
 sky130_fd_sc_hd__xor2_1 \U$$653  (.A(\t$4738 ),
    .B(net1242),
    .X(booth_b8_m49));
 sky130_fd_sc_hd__a22o_1 \U$$654  (.A1(net1682),
    .A2(net416),
    .B1(net1657),
    .B2(net682),
    .X(\t$4739 ));
 sky130_fd_sc_hd__xor2_1 \U$$655  (.A(\t$4739 ),
    .B(net1242),
    .X(booth_b8_m50));
 sky130_fd_sc_hd__a22o_1 \U$$656  (.A1(net1654),
    .A2(net411),
    .B1(net1646),
    .B2(net677),
    .X(\t$4740 ));
 sky130_fd_sc_hd__xor2_1 \U$$657  (.A(\t$4740 ),
    .B(net1238),
    .X(booth_b8_m51));
 sky130_fd_sc_hd__a22o_1 \U$$658  (.A1(net1648),
    .A2(net411),
    .B1(net1640),
    .B2(net677),
    .X(\t$4741 ));
 sky130_fd_sc_hd__xor2_1 \U$$659  (.A(\t$4741 ),
    .B(net1238),
    .X(booth_b8_m52));
 sky130_fd_sc_hd__a22o_1 \U$$66  (.A1(net1039),
    .A2(net442),
    .B1(net1023),
    .B2(net684),
    .X(\t$4440 ));
 sky130_fd_sc_hd__a22o_1 \U$$660  (.A1(net1638),
    .A2(net411),
    .B1(net1629),
    .B2(net677),
    .X(\t$4742 ));
 sky130_fd_sc_hd__xor2_1 \U$$661  (.A(\t$4742 ),
    .B(net1237),
    .X(booth_b8_m53));
 sky130_fd_sc_hd__a22o_1 \U$$662  (.A1(net1629),
    .A2(net411),
    .B1(net1620),
    .B2(net677),
    .X(\t$4743 ));
 sky130_fd_sc_hd__xor2_1 \U$$663  (.A(\t$4743 ),
    .B(net1237),
    .X(booth_b8_m54));
 sky130_fd_sc_hd__a22o_1 \U$$664  (.A1(net1620),
    .A2(net411),
    .B1(net1612),
    .B2(net677),
    .X(\t$4744 ));
 sky130_fd_sc_hd__xor2_1 \U$$665  (.A(\t$4744 ),
    .B(net1237),
    .X(booth_b8_m55));
 sky130_fd_sc_hd__a22o_1 \U$$666  (.A1(net1612),
    .A2(net411),
    .B1(net1604),
    .B2(net677),
    .X(\t$4745 ));
 sky130_fd_sc_hd__xor2_1 \U$$667  (.A(\t$4745 ),
    .B(net1237),
    .X(booth_b8_m56));
 sky130_fd_sc_hd__a22o_1 \U$$668  (.A1(net1607),
    .A2(net417),
    .B1(net1599),
    .B2(net683),
    .X(\t$4746 ));
 sky130_fd_sc_hd__xor2_1 \U$$669  (.A(\t$4746 ),
    .B(net1242),
    .X(booth_b8_m57));
 sky130_fd_sc_hd__xor2_1 \U$$67  (.A(\t$4440 ),
    .B(net1568),
    .X(booth_b0_m30));
 sky130_fd_sc_hd__a22o_1 \U$$670  (.A1(net1599),
    .A2(net416),
    .B1(net1590),
    .B2(net682),
    .X(\t$4747 ));
 sky130_fd_sc_hd__xor2_1 \U$$671  (.A(\t$4747 ),
    .B(net1242),
    .X(booth_b8_m58));
 sky130_fd_sc_hd__a22o_1 \U$$672  (.A1(net1590),
    .A2(net416),
    .B1(net1582),
    .B2(net682),
    .X(\t$4748 ));
 sky130_fd_sc_hd__xor2_1 \U$$673  (.A(\t$4748 ),
    .B(net1243),
    .X(booth_b8_m59));
 sky130_fd_sc_hd__a22o_1 \U$$674  (.A1(net1582),
    .A2(net416),
    .B1(net1555),
    .B2(net682),
    .X(\t$4749 ));
 sky130_fd_sc_hd__xor2_1 \U$$675  (.A(\t$4749 ),
    .B(net1243),
    .X(booth_b8_m60));
 sky130_fd_sc_hd__a22o_1 \U$$676  (.A1(net1555),
    .A2(net416),
    .B1(net1547),
    .B2(net682),
    .X(\t$4750 ));
 sky130_fd_sc_hd__xor2_1 \U$$677  (.A(\t$4750 ),
    .B(net1242),
    .X(booth_b8_m61));
 sky130_fd_sc_hd__a22o_1 \U$$678  (.A1(net1547),
    .A2(net416),
    .B1(net1539),
    .B2(net682),
    .X(\t$4751 ));
 sky130_fd_sc_hd__xor2_1 \U$$679  (.A(\t$4751 ),
    .B(net1242),
    .X(booth_b8_m62));
 sky130_fd_sc_hd__a22o_1 \U$$68  (.A1(net1023),
    .A2(net442),
    .B1(net1015),
    .B2(net684),
    .X(\t$4441 ));
 sky130_fd_sc_hd__a22o_1 \U$$680  (.A1(net1535),
    .A2(net411),
    .B1(net1527),
    .B2(net677),
    .X(\t$4752 ));
 sky130_fd_sc_hd__xor2_1 \U$$681  (.A(\t$4752 ),
    .B(net1237),
    .X(booth_b8_m63));
 sky130_fd_sc_hd__a22o_1 \U$$682  (.A1(net1527),
    .A2(net412),
    .B1(net1884),
    .B2(net678),
    .X(\t$4753 ));
 sky130_fd_sc_hd__xor2_1 \U$$683  (.A(\t$4753 ),
    .B(net1238),
    .X(booth_b8_m64));
 sky130_fd_sc_hd__inv_1 \U$$684  (.A(net1237),
    .Y(\notsign$4754 ));
 sky130_fd_sc_hd__inv_1 \U$$685  (.A(net1238),
    .Y(\notblock$4755[0] ));
 sky130_fd_sc_hd__inv_1 \U$$686  (.A(net2),
    .Y(\notblock$4755[1] ));
 sky130_fd_sc_hd__inv_1 \U$$687  (.A(net1417),
    .Y(\notblock$4755[2] ));
 sky130_fd_sc_hd__and2_1 \U$$688  (.A(net1417),
    .B(\notblock$4755[1] ),
    .X(\t$4756 ));
 sky130_fd_sc_hd__a32o_1 \U$$689  (.A1(\notblock$4755[2] ),
    .A2(net2),
    .A3(net1238),
    .B1(\t$4756 ),
    .B2(\notblock$4755[0] ),
    .X(\sel_0$4757 ));
 sky130_fd_sc_hd__xor2_1 \U$$69  (.A(\t$4441 ),
    .B(net1568),
    .X(booth_b0_m31));
 sky130_fd_sc_hd__xor2_1 \U$$690  (.A(net2),
    .B(net1238),
    .X(\sel_1$4758 ));
 sky130_fd_sc_hd__a22o_1 \U$$691  (.A1(net1885),
    .A2(net404),
    .B1(net1231),
    .B2(net670),
    .X(\t$4759 ));
 sky130_fd_sc_hd__xor2_1 \U$$692  (.A(\t$4759 ),
    .B(net1414),
    .X(booth_b10_m0));
 sky130_fd_sc_hd__a22o_1 \U$$693  (.A1(net1230),
    .A2(net404),
    .B1(net1126),
    .B2(net670),
    .X(\t$4760 ));
 sky130_fd_sc_hd__xor2_1 \U$$694  (.A(\t$4760 ),
    .B(net1414),
    .X(booth_b10_m1));
 sky130_fd_sc_hd__a22o_1 \U$$695  (.A1(net1127),
    .A2(net404),
    .B1(net1035),
    .B2(net670),
    .X(\t$4761 ));
 sky130_fd_sc_hd__xor2_1 \U$$696  (.A(\t$4761 ),
    .B(net1414),
    .X(booth_b10_m2));
 sky130_fd_sc_hd__a22o_1 \U$$697  (.A1(net1036),
    .A2(net404),
    .B1(net936),
    .B2(net670),
    .X(\t$4762 ));
 sky130_fd_sc_hd__xor2_1 \U$$698  (.A(\t$4762 ),
    .B(net1414),
    .X(booth_b10_m3));
 sky130_fd_sc_hd__a22o_1 \U$$699  (.A1(net933),
    .A2(net406),
    .B1(net1672),
    .B2(net672),
    .X(\t$4763 ));
 sky130_fd_sc_hd__xor2_1 \U$$7  (.A(\t$4410 ),
    .B(net1574),
    .X(booth_b0_m0));
 sky130_fd_sc_hd__a22o_1 \U$$70  (.A1(net1016),
    .A2(net442),
    .B1(net999),
    .B2(net684),
    .X(\t$4442 ));
 sky130_fd_sc_hd__xor2_1 \U$$700  (.A(\t$4763 ),
    .B(net1415),
    .X(booth_b10_m4));
 sky130_fd_sc_hd__a22o_1 \U$$701  (.A1(net1672),
    .A2(net406),
    .B1(net1561),
    .B2(net672),
    .X(\t$4764 ));
 sky130_fd_sc_hd__xor2_1 \U$$702  (.A(\t$4764 ),
    .B(net1415),
    .X(booth_b10_m5));
 sky130_fd_sc_hd__a22o_1 \U$$703  (.A1(net1561),
    .A2(net402),
    .B1(net1522),
    .B2(net668),
    .X(\t$4765 ));
 sky130_fd_sc_hd__xor2_1 \U$$704  (.A(\t$4765 ),
    .B(net1412),
    .X(booth_b10_m6));
 sky130_fd_sc_hd__a22o_1 \U$$705  (.A1(net1519),
    .A2(net402),
    .B1(net1513),
    .B2(net668),
    .X(\t$4766 ));
 sky130_fd_sc_hd__xor2_1 \U$$706  (.A(\t$4766 ),
    .B(net1412),
    .X(booth_b10_m7));
 sky130_fd_sc_hd__a22o_1 \U$$707  (.A1(net1513),
    .A2(net406),
    .B1(net1505),
    .B2(net672),
    .X(\t$4767 ));
 sky130_fd_sc_hd__xor2_1 \U$$708  (.A(\t$4767 ),
    .B(net1415),
    .X(booth_b10_m8));
 sky130_fd_sc_hd__a22o_1 \U$$709  (.A1(net1508),
    .A2(net404),
    .B1(net1499),
    .B2(net670),
    .X(\t$4768 ));
 sky130_fd_sc_hd__xor2_1 \U$$71  (.A(\t$4442 ),
    .B(net1569),
    .X(booth_b0_m32));
 sky130_fd_sc_hd__xor2_1 \U$$710  (.A(\t$4768 ),
    .B(net1414),
    .X(booth_b10_m9));
 sky130_fd_sc_hd__a22o_1 \U$$711  (.A1(net1499),
    .A2(net404),
    .B1(net1224),
    .B2(net670),
    .X(\t$4769 ));
 sky130_fd_sc_hd__xor2_1 \U$$712  (.A(\t$4769 ),
    .B(net1414),
    .X(booth_b10_m10));
 sky130_fd_sc_hd__a22o_1 \U$$713  (.A1(net1224),
    .A2(net404),
    .B1(net1216),
    .B2(net670),
    .X(\t$4770 ));
 sky130_fd_sc_hd__xor2_1 \U$$714  (.A(\t$4770 ),
    .B(net1414),
    .X(booth_b10_m11));
 sky130_fd_sc_hd__a22o_1 \U$$715  (.A1(net1211),
    .A2(net406),
    .B1(net1204),
    .B2(net672),
    .X(\t$4771 ));
 sky130_fd_sc_hd__xor2_1 \U$$716  (.A(\t$4771 ),
    .B(net1415),
    .X(booth_b10_m12));
 sky130_fd_sc_hd__a22o_1 \U$$717  (.A1(net1204),
    .A2(net406),
    .B1(net1194),
    .B2(net672),
    .X(\t$4772 ));
 sky130_fd_sc_hd__xor2_1 \U$$718  (.A(\t$4772 ),
    .B(net1415),
    .X(booth_b10_m13));
 sky130_fd_sc_hd__a22o_1 \U$$719  (.A1(net1194),
    .A2(net402),
    .B1(net1175),
    .B2(net668),
    .X(\t$4773 ));
 sky130_fd_sc_hd__a22o_1 \U$$72  (.A1(net1000),
    .A2(net447),
    .B1(net992),
    .B2(net689),
    .X(\t$4443 ));
 sky130_fd_sc_hd__xor2_1 \U$$720  (.A(\t$4773 ),
    .B(net1415),
    .X(booth_b10_m14));
 sky130_fd_sc_hd__a22o_1 \U$$721  (.A1(net1174),
    .A2(net402),
    .B1(net1164),
    .B2(net668),
    .X(\t$4774 ));
 sky130_fd_sc_hd__xor2_1 \U$$722  (.A(\t$4774 ),
    .B(net1412),
    .X(booth_b10_m15));
 sky130_fd_sc_hd__a22o_1 \U$$723  (.A1(net1164),
    .A2(net401),
    .B1(net1155),
    .B2(net667),
    .X(\t$4775 ));
 sky130_fd_sc_hd__xor2_1 \U$$724  (.A(\t$4775 ),
    .B(net1412),
    .X(booth_b10_m16));
 sky130_fd_sc_hd__a22o_1 \U$$725  (.A1(net1155),
    .A2(net401),
    .B1(net1146),
    .B2(net667),
    .X(\t$4776 ));
 sky130_fd_sc_hd__xor2_1 \U$$726  (.A(\t$4776 ),
    .B(net1412),
    .X(booth_b10_m17));
 sky130_fd_sc_hd__a22o_1 \U$$727  (.A1(net1146),
    .A2(net401),
    .B1(net1138),
    .B2(net667),
    .X(\t$4777 ));
 sky130_fd_sc_hd__xor2_1 \U$$728  (.A(\t$4777 ),
    .B(net1412),
    .X(booth_b10_m18));
 sky130_fd_sc_hd__a22o_1 \U$$729  (.A1(net1138),
    .A2(net401),
    .B1(net1130),
    .B2(net667),
    .X(\t$4778 ));
 sky130_fd_sc_hd__xor2_1 \U$$73  (.A(\t$4443 ),
    .B(net1574),
    .X(booth_b0_m33));
 sky130_fd_sc_hd__xor2_1 \U$$730  (.A(\t$4778 ),
    .B(net1412),
    .X(booth_b10_m19));
 sky130_fd_sc_hd__a22o_1 \U$$731  (.A1(net1130),
    .A2(net401),
    .B1(net1114),
    .B2(net667),
    .X(\t$4779 ));
 sky130_fd_sc_hd__xor2_1 \U$$732  (.A(\t$4779 ),
    .B(net1412),
    .X(booth_b10_m20));
 sky130_fd_sc_hd__a22o_1 \U$$733  (.A1(net1114),
    .A2(net402),
    .B1(net1105),
    .B2(net668),
    .X(\t$4780 ));
 sky130_fd_sc_hd__xor2_1 \U$$734  (.A(\t$4780 ),
    .B(net1412),
    .X(booth_b10_m21));
 sky130_fd_sc_hd__a22o_1 \U$$735  (.A1(net1106),
    .A2(net402),
    .B1(net1099),
    .B2(net668),
    .X(\t$4781 ));
 sky130_fd_sc_hd__xor2_1 \U$$736  (.A(\t$4781 ),
    .B(net1413),
    .X(booth_b10_m22));
 sky130_fd_sc_hd__a22o_1 \U$$737  (.A1(net1100),
    .A2(net404),
    .B1(net1091),
    .B2(net670),
    .X(\t$4782 ));
 sky130_fd_sc_hd__xor2_1 \U$$738  (.A(\t$4782 ),
    .B(net1414),
    .X(booth_b10_m23));
 sky130_fd_sc_hd__a22o_1 \U$$739  (.A1(net1091),
    .A2(net405),
    .B1(net1083),
    .B2(net671),
    .X(\t$4783 ));
 sky130_fd_sc_hd__a22o_1 \U$$74  (.A1(net992),
    .A2(net448),
    .B1(net987),
    .B2(net690),
    .X(\t$4444 ));
 sky130_fd_sc_hd__xor2_1 \U$$740  (.A(\t$4783 ),
    .B(net1414),
    .X(booth_b10_m24));
 sky130_fd_sc_hd__a22o_1 \U$$741  (.A1(net1084),
    .A2(net404),
    .B1(net1075),
    .B2(net670),
    .X(\t$4784 ));
 sky130_fd_sc_hd__xor2_1 \U$$742  (.A(\t$4784 ),
    .B(net1414),
    .X(booth_b10_m25));
 sky130_fd_sc_hd__a22o_1 \U$$743  (.A1(net1074),
    .A2(net405),
    .B1(net1066),
    .B2(net671),
    .X(\t$4785 ));
 sky130_fd_sc_hd__xor2_1 \U$$744  (.A(\t$4785 ),
    .B(net1416),
    .X(booth_b10_m26));
 sky130_fd_sc_hd__a22o_1 \U$$745  (.A1(net1066),
    .A2(net406),
    .B1(net1057),
    .B2(net672),
    .X(\t$4786 ));
 sky130_fd_sc_hd__xor2_1 \U$$746  (.A(\t$4786 ),
    .B(net1416),
    .X(booth_b10_m27));
 sky130_fd_sc_hd__a22o_1 \U$$747  (.A1(net1056),
    .A2(net406),
    .B1(net1048),
    .B2(net672),
    .X(\t$4787 ));
 sky130_fd_sc_hd__xor2_1 \U$$748  (.A(\t$4787 ),
    .B(net1415),
    .X(booth_b10_m28));
 sky130_fd_sc_hd__a22o_1 \U$$749  (.A1(net1049),
    .A2(net406),
    .B1(net1041),
    .B2(net672),
    .X(\t$4788 ));
 sky130_fd_sc_hd__xor2_1 \U$$75  (.A(\t$4444 ),
    .B(net1574),
    .X(booth_b0_m34));
 sky130_fd_sc_hd__xor2_1 \U$$750  (.A(\t$4788 ),
    .B(net1415),
    .X(booth_b10_m29));
 sky130_fd_sc_hd__a22o_1 \U$$751  (.A1(net1040),
    .A2(net402),
    .B1(net1024),
    .B2(net668),
    .X(\t$4789 ));
 sky130_fd_sc_hd__xor2_1 \U$$752  (.A(\t$4789 ),
    .B(net1412),
    .X(booth_b10_m30));
 sky130_fd_sc_hd__a22o_1 \U$$753  (.A1(net1023),
    .A2(net401),
    .B1(net1015),
    .B2(net667),
    .X(\t$4790 ));
 sky130_fd_sc_hd__xor2_1 \U$$754  (.A(\t$4790 ),
    .B(net1413),
    .X(booth_b10_m31));
 sky130_fd_sc_hd__a22o_1 \U$$755  (.A1(net1015),
    .A2(net401),
    .B1(net998),
    .B2(net667),
    .X(\t$4791 ));
 sky130_fd_sc_hd__xor2_1 \U$$756  (.A(\t$4791 ),
    .B(net1413),
    .X(booth_b10_m32));
 sky130_fd_sc_hd__a22o_1 \U$$757  (.A1(net998),
    .A2(net402),
    .B1(net990),
    .B2(net668),
    .X(\t$4792 ));
 sky130_fd_sc_hd__xor2_1 \U$$758  (.A(\t$4792 ),
    .B(net1413),
    .X(booth_b10_m33));
 sky130_fd_sc_hd__a22o_1 \U$$759  (.A1(net990),
    .A2(net402),
    .B1(net982),
    .B2(net668),
    .X(\t$4793 ));
 sky130_fd_sc_hd__a22o_1 \U$$76  (.A1(net987),
    .A2(net448),
    .B1(net977),
    .B2(net690),
    .X(\t$4445 ));
 sky130_fd_sc_hd__xor2_1 \U$$760  (.A(\t$4793 ),
    .B(net1413),
    .X(booth_b10_m34));
 sky130_fd_sc_hd__a22o_1 \U$$761  (.A1(net986),
    .A2(net406),
    .B1(net981),
    .B2(net672),
    .X(\t$4794 ));
 sky130_fd_sc_hd__xor2_1 \U$$762  (.A(\t$4794 ),
    .B(net1416),
    .X(booth_b10_m35));
 sky130_fd_sc_hd__a22o_1 \U$$763  (.A1(net973),
    .A2(net401),
    .B1(net964),
    .B2(net667),
    .X(\t$4795 ));
 sky130_fd_sc_hd__xor2_1 \U$$764  (.A(\t$4795 ),
    .B(net1413),
    .X(booth_b10_m36));
 sky130_fd_sc_hd__a22o_1 \U$$765  (.A1(net964),
    .A2(net401),
    .B1(net956),
    .B2(net667),
    .X(\t$4796 ));
 sky130_fd_sc_hd__xor2_1 \U$$766  (.A(\t$4796 ),
    .B(net1413),
    .X(booth_b10_m37));
 sky130_fd_sc_hd__a22o_1 \U$$767  (.A1(net956),
    .A2(net401),
    .B1(net948),
    .B2(net667),
    .X(\t$4797 ));
 sky130_fd_sc_hd__xor2_1 \U$$768  (.A(\t$4797 ),
    .B(net1413),
    .X(booth_b10_m38));
 sky130_fd_sc_hd__a22o_1 \U$$769  (.A1(net949),
    .A2(net403),
    .B1(net941),
    .B2(net669),
    .X(\t$4798 ));
 sky130_fd_sc_hd__xor2_1 \U$$77  (.A(\t$4445 ),
    .B(net1575),
    .X(booth_b0_m35));
 sky130_fd_sc_hd__xor2_1 \U$$770  (.A(\t$4798 ),
    .B(net1418),
    .X(booth_b10_m39));
 sky130_fd_sc_hd__a22o_1 \U$$771  (.A1(net940),
    .A2(net403),
    .B1(net924),
    .B2(net669),
    .X(\t$4799 ));
 sky130_fd_sc_hd__xor2_1 \U$$772  (.A(\t$4799 ),
    .B(net1418),
    .X(booth_b10_m40));
 sky130_fd_sc_hd__a22o_1 \U$$773  (.A1(net931),
    .A2(net407),
    .B1(net1749),
    .B2(net673),
    .X(\t$4800 ));
 sky130_fd_sc_hd__xor2_1 \U$$774  (.A(\t$4800 ),
    .B(net1416),
    .X(booth_b10_m41));
 sky130_fd_sc_hd__a22o_1 \U$$775  (.A1(net1749),
    .A2(net405),
    .B1(net1741),
    .B2(net671),
    .X(\t$4801 ));
 sky130_fd_sc_hd__xor2_1 \U$$776  (.A(\t$4801 ),
    .B(net1416),
    .X(booth_b10_m42));
 sky130_fd_sc_hd__a22o_1 \U$$777  (.A1(net1744),
    .A2(net405),
    .B1(net1736),
    .B2(net671),
    .X(\t$4802 ));
 sky130_fd_sc_hd__xor2_1 \U$$778  (.A(\t$4802 ),
    .B(net1416),
    .X(booth_b10_m43));
 sky130_fd_sc_hd__a22o_1 \U$$779  (.A1(net1736),
    .A2(net405),
    .B1(net1725),
    .B2(net671),
    .X(\t$4803 ));
 sky130_fd_sc_hd__a22o_1 \U$$78  (.A1(net977),
    .A2(net448),
    .B1(net969),
    .B2(net690),
    .X(\t$4446 ));
 sky130_fd_sc_hd__xor2_1 \U$$780  (.A(\t$4803 ),
    .B(net1416),
    .X(booth_b10_m44));
 sky130_fd_sc_hd__a22o_1 \U$$781  (.A1(net1724),
    .A2(net404),
    .B1(net1715),
    .B2(net670),
    .X(\t$4804 ));
 sky130_fd_sc_hd__xor2_1 \U$$782  (.A(\t$4804 ),
    .B(net1416),
    .X(booth_b10_m45));
 sky130_fd_sc_hd__a22o_1 \U$$783  (.A1(net1716),
    .A2(net407),
    .B1(net1707),
    .B2(net673),
    .X(\t$4805 ));
 sky130_fd_sc_hd__xor2_1 \U$$784  (.A(\t$4805 ),
    .B(net1419),
    .X(booth_b10_m46));
 sky130_fd_sc_hd__a22o_1 \U$$785  (.A1(net1706),
    .A2(net405),
    .B1(net1698),
    .B2(net671),
    .X(\t$4806 ));
 sky130_fd_sc_hd__xor2_1 \U$$786  (.A(\t$4806 ),
    .B(net1416),
    .X(booth_b10_m47));
 sky130_fd_sc_hd__a22o_1 \U$$787  (.A1(net1698),
    .A2(net407),
    .B1(net1690),
    .B2(net673),
    .X(\t$4807 ));
 sky130_fd_sc_hd__xor2_1 \U$$788  (.A(\t$4807 ),
    .B(net1419),
    .X(booth_b10_m48));
 sky130_fd_sc_hd__a22o_1 \U$$789  (.A1(net1689),
    .A2(net408),
    .B1(net1679),
    .B2(net674),
    .X(\t$4808 ));
 sky130_fd_sc_hd__xor2_1 \U$$79  (.A(\t$4446 ),
    .B(net1575),
    .X(booth_b0_m36));
 sky130_fd_sc_hd__xor2_1 \U$$790  (.A(\t$4808 ),
    .B(net1418),
    .X(booth_b10_m49));
 sky130_fd_sc_hd__a22o_1 \U$$791  (.A1(net1681),
    .A2(net408),
    .B1(net1656),
    .B2(net674),
    .X(\t$4809 ));
 sky130_fd_sc_hd__xor2_1 \U$$792  (.A(\t$4809 ),
    .B(net1419),
    .X(booth_b10_m50));
 sky130_fd_sc_hd__a22o_1 \U$$793  (.A1(net1654),
    .A2(net403),
    .B1(net1646),
    .B2(net669),
    .X(\t$4810 ));
 sky130_fd_sc_hd__xor2_1 \U$$794  (.A(\t$4810 ),
    .B(net1418),
    .X(booth_b10_m51));
 sky130_fd_sc_hd__a22o_1 \U$$795  (.A1(net1646),
    .A2(net403),
    .B1(net1638),
    .B2(net669),
    .X(\t$4811 ));
 sky130_fd_sc_hd__xor2_1 \U$$796  (.A(\t$4811 ),
    .B(net1418),
    .X(booth_b10_m52));
 sky130_fd_sc_hd__a22o_1 \U$$797  (.A1(net1638),
    .A2(net403),
    .B1(net1629),
    .B2(net669),
    .X(\t$4812 ));
 sky130_fd_sc_hd__xor2_1 \U$$798  (.A(\t$4812 ),
    .B(net1418),
    .X(booth_b10_m53));
 sky130_fd_sc_hd__a22o_1 \U$$799  (.A1(net1630),
    .A2(net403),
    .B1(net1620),
    .B2(net669),
    .X(\t$4813 ));
 sky130_fd_sc_hd__a22o_1 \U$$8  (.A1(net1232),
    .A2(net446),
    .B1(net1127),
    .B2(net688),
    .X(\t$4411 ));
 sky130_fd_sc_hd__a22o_1 \U$$80  (.A1(net964),
    .A2(net442),
    .B1(net956),
    .B2(net684),
    .X(\t$4447 ));
 sky130_fd_sc_hd__xor2_1 \U$$800  (.A(\t$4813 ),
    .B(net1417),
    .X(booth_b10_m54));
 sky130_fd_sc_hd__a22o_1 \U$$801  (.A1(net1623),
    .A2(net407),
    .B1(net1615),
    .B2(net673),
    .X(\t$4814 ));
 sky130_fd_sc_hd__xor2_1 \U$$802  (.A(\t$4814 ),
    .B(net1419),
    .X(booth_b10_m55));
 sky130_fd_sc_hd__a22o_1 \U$$803  (.A1(net1615),
    .A2(net407),
    .B1(net1607),
    .B2(net673),
    .X(\t$4815 ));
 sky130_fd_sc_hd__xor2_1 \U$$804  (.A(\t$4815 ),
    .B(net1419),
    .X(booth_b10_m56));
 sky130_fd_sc_hd__a22o_1 \U$$805  (.A1(net1607),
    .A2(net407),
    .B1(net1599),
    .B2(net673),
    .X(\t$4816 ));
 sky130_fd_sc_hd__xor2_1 \U$$806  (.A(\t$4816 ),
    .B(net1419),
    .X(booth_b10_m57));
 sky130_fd_sc_hd__a22o_1 \U$$807  (.A1(net1599),
    .A2(net407),
    .B1(net1590),
    .B2(net673),
    .X(\t$4817 ));
 sky130_fd_sc_hd__xor2_1 \U$$808  (.A(\t$4817 ),
    .B(net1419),
    .X(booth_b10_m58));
 sky130_fd_sc_hd__a22o_1 \U$$809  (.A1(net1590),
    .A2(net407),
    .B1(net1582),
    .B2(net673),
    .X(\t$4818 ));
 sky130_fd_sc_hd__xor2_1 \U$$81  (.A(\t$4447 ),
    .B(net1568),
    .X(booth_b0_m37));
 sky130_fd_sc_hd__xor2_1 \U$$810  (.A(\t$4818 ),
    .B(net1419),
    .X(booth_b10_m59));
 sky130_fd_sc_hd__a22o_1 \U$$811  (.A1(net1582),
    .A2(net408),
    .B1(net1555),
    .B2(net674),
    .X(\t$4819 ));
 sky130_fd_sc_hd__xor2_1 \U$$812  (.A(\t$4819 ),
    .B(net1419),
    .X(booth_b10_m60));
 sky130_fd_sc_hd__a22o_1 \U$$813  (.A1(net1551),
    .A2(net403),
    .B1(net1543),
    .B2(net669),
    .X(\t$4820 ));
 sky130_fd_sc_hd__xor2_1 \U$$814  (.A(\t$4820 ),
    .B(net1417),
    .X(booth_b10_m61));
 sky130_fd_sc_hd__a22o_1 \U$$815  (.A1(net1543),
    .A2(net403),
    .B1(net1535),
    .B2(net669),
    .X(\t$4821 ));
 sky130_fd_sc_hd__xor2_1 \U$$816  (.A(\t$4821 ),
    .B(net1418),
    .X(booth_b10_m62));
 sky130_fd_sc_hd__a22o_1 \U$$817  (.A1(net1535),
    .A2(net403),
    .B1(net1527),
    .B2(net669),
    .X(\t$4822 ));
 sky130_fd_sc_hd__xor2_1 \U$$818  (.A(\t$4822 ),
    .B(net1417),
    .X(booth_b10_m63));
 sky130_fd_sc_hd__a22o_1 \U$$819  (.A1(net1527),
    .A2(net403),
    .B1(net1886),
    .B2(net669),
    .X(\t$4823 ));
 sky130_fd_sc_hd__a22o_1 \U$$82  (.A1(net960),
    .A2(net443),
    .B1(net952),
    .B2(net685),
    .X(\t$4448 ));
 sky130_fd_sc_hd__xor2_1 \U$$820  (.A(\t$4823 ),
    .B(net1417),
    .X(booth_b10_m64));
 sky130_fd_sc_hd__inv_1 \U$$821  (.A(net1417),
    .Y(\notsign$4824 ));
 sky130_fd_sc_hd__inv_1 \U$$822  (.A(net1417),
    .Y(\notblock$4825[0] ));
 sky130_fd_sc_hd__inv_1 \U$$823  (.A(net4),
    .Y(\notblock$4825[1] ));
 sky130_fd_sc_hd__inv_1 \U$$824  (.A(net1316),
    .Y(\notblock$4825[2] ));
 sky130_fd_sc_hd__and2_1 \U$$825  (.A(net1316),
    .B(\notblock$4825[1] ),
    .X(\t$4826 ));
 sky130_fd_sc_hd__a32o_1 \U$$826  (.A1(\notblock$4825[2] ),
    .A2(net4),
    .A3(net1417),
    .B1(\t$4826 ),
    .B2(\notblock$4825[0] ),
    .X(\sel_0$4827 ));
 sky130_fd_sc_hd__xor2_1 \U$$827  (.A(net4),
    .B(net1417),
    .X(\sel_1$4828 ));
 sky130_fd_sc_hd__a22o_1 \U$$828  (.A1(net1887),
    .A2(net397),
    .B1(net1231),
    .B2(net663),
    .X(\t$4829 ));
 sky130_fd_sc_hd__xor2_1 \U$$829  (.A(\t$4829 ),
    .B(net1312),
    .X(booth_b12_m0));
 sky130_fd_sc_hd__xor2_1 \U$$83  (.A(\t$4448 ),
    .B(net1569),
    .X(booth_b0_m38));
 sky130_fd_sc_hd__a22o_1 \U$$830  (.A1(net1231),
    .A2(net397),
    .B1(net1127),
    .B2(net663),
    .X(\t$4830 ));
 sky130_fd_sc_hd__xor2_1 \U$$831  (.A(\t$4830 ),
    .B(net1312),
    .X(booth_b12_m1));
 sky130_fd_sc_hd__a22o_1 \U$$832  (.A1(net1123),
    .A2(net396),
    .B1(net1032),
    .B2(net662),
    .X(\t$4831 ));
 sky130_fd_sc_hd__xor2_1 \U$$833  (.A(\t$4831 ),
    .B(net1312),
    .X(booth_b12_m2));
 sky130_fd_sc_hd__a22o_1 \U$$834  (.A1(net1032),
    .A2(net396),
    .B1(net933),
    .B2(net662),
    .X(\t$4832 ));
 sky130_fd_sc_hd__xor2_1 \U$$835  (.A(\t$4832 ),
    .B(net1312),
    .X(booth_b12_m3));
 sky130_fd_sc_hd__a22o_1 \U$$836  (.A1(net933),
    .A2(net394),
    .B1(net1672),
    .B2(net660),
    .X(\t$4833 ));
 sky130_fd_sc_hd__xor2_1 \U$$837  (.A(\t$4833 ),
    .B(net1310),
    .X(booth_b12_m4));
 sky130_fd_sc_hd__a22o_1 \U$$838  (.A1(net1672),
    .A2(net394),
    .B1(net1561),
    .B2(net660),
    .X(\t$4834 ));
 sky130_fd_sc_hd__xor2_1 \U$$839  (.A(\t$4834 ),
    .B(net1310),
    .X(booth_b12_m5));
 sky130_fd_sc_hd__a22o_1 \U$$84  (.A1(net952),
    .A2(net448),
    .B1(net947),
    .B2(net690),
    .X(\t$4449 ));
 sky130_fd_sc_hd__a22o_1 \U$$840  (.A1(net1561),
    .A2(net396),
    .B1(net1522),
    .B2(net662),
    .X(\t$4835 ));
 sky130_fd_sc_hd__xor2_1 \U$$841  (.A(\t$4835 ),
    .B(net1312),
    .X(booth_b12_m6));
 sky130_fd_sc_hd__a22o_1 \U$$842  (.A1(net1523),
    .A2(net396),
    .B1(net1515),
    .B2(net662),
    .X(\t$4836 ));
 sky130_fd_sc_hd__xor2_1 \U$$843  (.A(\t$4836 ),
    .B(net1312),
    .X(booth_b12_m7));
 sky130_fd_sc_hd__a22o_1 \U$$844  (.A1(net1515),
    .A2(net396),
    .B1(net1508),
    .B2(net662),
    .X(\t$4837 ));
 sky130_fd_sc_hd__xor2_1 \U$$845  (.A(\t$4837 ),
    .B(net1312),
    .X(booth_b12_m8));
 sky130_fd_sc_hd__a22o_1 \U$$846  (.A1(net1508),
    .A2(net397),
    .B1(net1499),
    .B2(net663),
    .X(\t$4838 ));
 sky130_fd_sc_hd__xor2_1 \U$$847  (.A(\t$4838 ),
    .B(net1313),
    .X(booth_b12_m9));
 sky130_fd_sc_hd__a22o_1 \U$$848  (.A1(net1496),
    .A2(net396),
    .B1(net1221),
    .B2(net662),
    .X(\t$4839 ));
 sky130_fd_sc_hd__xor2_1 \U$$849  (.A(\t$4839 ),
    .B(net1312),
    .X(booth_b12_m10));
 sky130_fd_sc_hd__xor2_1 \U$$85  (.A(\t$4449 ),
    .B(net1575),
    .X(booth_b0_m39));
 sky130_fd_sc_hd__a22o_1 \U$$850  (.A1(net1221),
    .A2(net396),
    .B1(net1212),
    .B2(net662),
    .X(\t$4840 ));
 sky130_fd_sc_hd__xor2_1 \U$$851  (.A(\t$4840 ),
    .B(net1312),
    .X(booth_b12_m11));
 sky130_fd_sc_hd__a22o_1 \U$$852  (.A1(net1211),
    .A2(net394),
    .B1(net1203),
    .B2(net660),
    .X(\t$4841 ));
 sky130_fd_sc_hd__xor2_1 \U$$853  (.A(\t$4841 ),
    .B(net1310),
    .X(booth_b12_m12));
 sky130_fd_sc_hd__a22o_1 \U$$854  (.A1(net1202),
    .A2(net394),
    .B1(net1193),
    .B2(net660),
    .X(\t$4842 ));
 sky130_fd_sc_hd__xor2_1 \U$$855  (.A(\t$4842 ),
    .B(net1310),
    .X(booth_b12_m13));
 sky130_fd_sc_hd__a22o_1 \U$$856  (.A1(net1192),
    .A2(net393),
    .B1(net1173),
    .B2(net659),
    .X(\t$4843 ));
 sky130_fd_sc_hd__xor2_1 \U$$857  (.A(\t$4843 ),
    .B(net1310),
    .X(booth_b12_m14));
 sky130_fd_sc_hd__a22o_1 \U$$858  (.A1(net1173),
    .A2(net393),
    .B1(net1164),
    .B2(net659),
    .X(\t$4844 ));
 sky130_fd_sc_hd__xor2_1 \U$$859  (.A(\t$4844 ),
    .B(net1310),
    .X(booth_b12_m15));
 sky130_fd_sc_hd__a22o_1 \U$$86  (.A1(net940),
    .A2(net442),
    .B1(net924),
    .B2(net684),
    .X(\t$4450 ));
 sky130_fd_sc_hd__a22o_1 \U$$860  (.A1(net1164),
    .A2(net393),
    .B1(net1155),
    .B2(net659),
    .X(\t$4845 ));
 sky130_fd_sc_hd__xor2_1 \U$$861  (.A(\t$4845 ),
    .B(net1310),
    .X(booth_b12_m16));
 sky130_fd_sc_hd__a22o_1 \U$$862  (.A1(net1155),
    .A2(net393),
    .B1(net1146),
    .B2(net659),
    .X(\t$4846 ));
 sky130_fd_sc_hd__xor2_1 \U$$863  (.A(\t$4846 ),
    .B(net1310),
    .X(booth_b12_m17));
 sky130_fd_sc_hd__a22o_1 \U$$864  (.A1(net1146),
    .A2(net393),
    .B1(net1138),
    .B2(net659),
    .X(\t$4847 ));
 sky130_fd_sc_hd__xor2_1 \U$$865  (.A(\t$4847 ),
    .B(net1310),
    .X(booth_b12_m18));
 sky130_fd_sc_hd__a22o_1 \U$$866  (.A1(net1138),
    .A2(net393),
    .B1(net1130),
    .B2(net659),
    .X(\t$4848 ));
 sky130_fd_sc_hd__xor2_1 \U$$867  (.A(\t$4848 ),
    .B(net1310),
    .X(booth_b12_m19));
 sky130_fd_sc_hd__a22o_1 \U$$868  (.A1(net1134),
    .A2(net396),
    .B1(net1118),
    .B2(net662),
    .X(\t$4849 ));
 sky130_fd_sc_hd__xor2_1 \U$$869  (.A(\t$4849 ),
    .B(net1314),
    .X(booth_b12_m20));
 sky130_fd_sc_hd__xor2_1 \U$$87  (.A(\t$4450 ),
    .B(net1568),
    .X(booth_b0_m40));
 sky130_fd_sc_hd__a22o_1 \U$$870  (.A1(net1117),
    .A2(net397),
    .B1(net1108),
    .B2(net663),
    .X(\t$4850 ));
 sky130_fd_sc_hd__xor2_1 \U$$871  (.A(\t$4850 ),
    .B(net1313),
    .X(booth_b12_m21));
 sky130_fd_sc_hd__a22o_1 \U$$872  (.A1(net1108),
    .A2(net397),
    .B1(net1100),
    .B2(net663),
    .X(\t$4851 ));
 sky130_fd_sc_hd__xor2_1 \U$$873  (.A(\t$4851 ),
    .B(net1313),
    .X(booth_b12_m22));
 sky130_fd_sc_hd__a22o_1 \U$$874  (.A1(net1101),
    .A2(net397),
    .B1(net1092),
    .B2(net663),
    .X(\t$4852 ));
 sky130_fd_sc_hd__xor2_1 \U$$875  (.A(\t$4852 ),
    .B(net1313),
    .X(booth_b12_m23));
 sky130_fd_sc_hd__a22o_1 \U$$876  (.A1(net1091),
    .A2(net397),
    .B1(net1083),
    .B2(net663),
    .X(\t$4853 ));
 sky130_fd_sc_hd__xor2_1 \U$$877  (.A(\t$4853 ),
    .B(net1314),
    .X(booth_b12_m24));
 sky130_fd_sc_hd__a22o_1 \U$$878  (.A1(net1083),
    .A2(net398),
    .B1(net1074),
    .B2(net664),
    .X(\t$4854 ));
 sky130_fd_sc_hd__xor2_1 \U$$879  (.A(\t$4854 ),
    .B(net1314),
    .X(booth_b12_m25));
 sky130_fd_sc_hd__a22o_1 \U$$88  (.A1(net924),
    .A2(net444),
    .B1(net1745),
    .B2(net686),
    .X(\t$4451 ));
 sky130_fd_sc_hd__a22o_1 \U$$880  (.A1(net1074),
    .A2(net396),
    .B1(net1066),
    .B2(net662),
    .X(\t$4855 ));
 sky130_fd_sc_hd__xor2_1 \U$$881  (.A(\t$4855 ),
    .B(net1312),
    .X(booth_b12_m26));
 sky130_fd_sc_hd__a22o_1 \U$$882  (.A1(net1064),
    .A2(net394),
    .B1(net1056),
    .B2(net660),
    .X(\t$4856 ));
 sky130_fd_sc_hd__xor2_1 \U$$883  (.A(\t$4856 ),
    .B(net1311),
    .X(booth_b12_m27));
 sky130_fd_sc_hd__a22o_1 \U$$884  (.A1(net1055),
    .A2(net394),
    .B1(net1047),
    .B2(net660),
    .X(\t$4857 ));
 sky130_fd_sc_hd__xor2_1 \U$$885  (.A(\t$4857 ),
    .B(net1311),
    .X(booth_b12_m28));
 sky130_fd_sc_hd__a22o_1 \U$$886  (.A1(net1047),
    .A2(net394),
    .B1(net1039),
    .B2(net660),
    .X(\t$4858 ));
 sky130_fd_sc_hd__xor2_1 \U$$887  (.A(\t$4858 ),
    .B(net1311),
    .X(booth_b12_m29));
 sky130_fd_sc_hd__a22o_1 \U$$888  (.A1(net1039),
    .A2(net393),
    .B1(net1023),
    .B2(net659),
    .X(\t$4859 ));
 sky130_fd_sc_hd__xor2_1 \U$$889  (.A(\t$4859 ),
    .B(net1311),
    .X(booth_b12_m30));
 sky130_fd_sc_hd__xor2_1 \U$$89  (.A(\t$4451 ),
    .B(net1570),
    .X(booth_b0_m41));
 sky130_fd_sc_hd__a22o_1 \U$$890  (.A1(net1023),
    .A2(net393),
    .B1(net1015),
    .B2(net659),
    .X(\t$4860 ));
 sky130_fd_sc_hd__xor2_1 \U$$891  (.A(\t$4860 ),
    .B(net1311),
    .X(booth_b12_m31));
 sky130_fd_sc_hd__a22o_1 \U$$892  (.A1(net1016),
    .A2(net394),
    .B1(net999),
    .B2(net660),
    .X(\t$4861 ));
 sky130_fd_sc_hd__xor2_1 \U$$893  (.A(\t$4861 ),
    .B(net1311),
    .X(booth_b12_m32));
 sky130_fd_sc_hd__a22o_1 \U$$894  (.A1(net999),
    .A2(net396),
    .B1(net991),
    .B2(net662),
    .X(\t$4862 ));
 sky130_fd_sc_hd__xor2_1 \U$$895  (.A(\t$4862 ),
    .B(net1314),
    .X(booth_b12_m33));
 sky130_fd_sc_hd__a22o_1 \U$$896  (.A1(net990),
    .A2(net393),
    .B1(net982),
    .B2(net659),
    .X(\t$4863 ));
 sky130_fd_sc_hd__xor2_1 \U$$897  (.A(\t$4863 ),
    .B(net1311),
    .X(booth_b12_m34));
 sky130_fd_sc_hd__a22o_1 \U$$898  (.A1(net982),
    .A2(net393),
    .B1(net973),
    .B2(net659),
    .X(\t$4864 ));
 sky130_fd_sc_hd__xor2_1 \U$$899  (.A(\t$4864 ),
    .B(net1311),
    .X(booth_b12_m35));
 sky130_fd_sc_hd__xor2_1 \U$$9  (.A(\t$4411 ),
    .B(net1574),
    .X(booth_b0_m1));
 sky130_fd_sc_hd__a22o_1 \U$$90  (.A1(net1745),
    .A2(net444),
    .B1(net1737),
    .B2(net686),
    .X(\t$4452 ));
 sky130_fd_sc_hd__a22o_1 \U$$900  (.A1(net973),
    .A2(net394),
    .B1(net964),
    .B2(net660),
    .X(\t$4865 ));
 sky130_fd_sc_hd__xor2_1 \U$$901  (.A(\t$4865 ),
    .B(net1311),
    .X(booth_b12_m36));
 sky130_fd_sc_hd__a22o_1 \U$$902  (.A1(net964),
    .A2(net395),
    .B1(net956),
    .B2(net661),
    .X(\t$4866 ));
 sky130_fd_sc_hd__xor2_1 \U$$903  (.A(\t$4866 ),
    .B(net1317),
    .X(booth_b12_m37));
 sky130_fd_sc_hd__a22o_1 \U$$904  (.A1(net960),
    .A2(net398),
    .B1(net952),
    .B2(net664),
    .X(\t$4867 ));
 sky130_fd_sc_hd__xor2_1 \U$$905  (.A(\t$4867 ),
    .B(net1314),
    .X(booth_b12_m38));
 sky130_fd_sc_hd__a22o_1 \U$$906  (.A1(net955),
    .A2(net397),
    .B1(net947),
    .B2(net663),
    .X(\t$4868 ));
 sky130_fd_sc_hd__xor2_1 \U$$907  (.A(\t$4868 ),
    .B(net1314),
    .X(booth_b12_m39));
 sky130_fd_sc_hd__a22o_1 \U$$908  (.A1(net944),
    .A2(net397),
    .B1(net928),
    .B2(net663),
    .X(\t$4869 ));
 sky130_fd_sc_hd__xor2_1 \U$$909  (.A(\t$4869 ),
    .B(net1314),
    .X(booth_b12_m40));
 sky130_fd_sc_hd__xor2_1 \U$$91  (.A(\t$4452 ),
    .B(net1570),
    .X(booth_b0_m42));
 sky130_fd_sc_hd__a22o_1 \U$$910  (.A1(net931),
    .A2(net397),
    .B1(net1752),
    .B2(net663),
    .X(\t$4870 ));
 sky130_fd_sc_hd__xor2_1 \U$$911  (.A(\t$4870 ),
    .B(net1314),
    .X(booth_b12_m41));
 sky130_fd_sc_hd__a22o_1 \U$$912  (.A1(net1752),
    .A2(net398),
    .B1(net1744),
    .B2(net664),
    .X(\t$4871 ));
 sky130_fd_sc_hd__xor2_1 \U$$913  (.A(\t$4871 ),
    .B(net1314),
    .X(booth_b12_m42));
 sky130_fd_sc_hd__a22o_1 \U$$914  (.A1(net1741),
    .A2(net398),
    .B1(net1733),
    .B2(net664),
    .X(\t$4872 ));
 sky130_fd_sc_hd__xor2_1 \U$$915  (.A(\t$4872 ),
    .B(net1315),
    .X(booth_b12_m43));
 sky130_fd_sc_hd__a22o_1 \U$$916  (.A1(net1733),
    .A2(net399),
    .B1(net1724),
    .B2(net665),
    .X(\t$4873 ));
 sky130_fd_sc_hd__xor2_1 \U$$917  (.A(\t$4873 ),
    .B(net1318),
    .X(booth_b12_m44));
 sky130_fd_sc_hd__a22o_1 \U$$918  (.A1(net1724),
    .A2(net398),
    .B1(net1715),
    .B2(net664),
    .X(\t$4874 ));
 sky130_fd_sc_hd__xor2_1 \U$$919  (.A(\t$4874 ),
    .B(net1315),
    .X(booth_b12_m45));
 sky130_fd_sc_hd__a22o_1 \U$$92  (.A1(net1737),
    .A2(net444),
    .B1(net1729),
    .B2(net686),
    .X(\t$4453 ));
 sky130_fd_sc_hd__a22o_1 \U$$920  (.A1(net1715),
    .A2(net399),
    .B1(net1706),
    .B2(net665),
    .X(\t$4875 ));
 sky130_fd_sc_hd__xor2_1 \U$$921  (.A(\t$4875 ),
    .B(net1314),
    .X(booth_b12_m46));
 sky130_fd_sc_hd__a22o_1 \U$$922  (.A1(net1705),
    .A2(net395),
    .B1(net1697),
    .B2(net661),
    .X(\t$4876 ));
 sky130_fd_sc_hd__xor2_1 \U$$923  (.A(\t$4876 ),
    .B(net1317),
    .X(booth_b12_m47));
 sky130_fd_sc_hd__a22o_1 \U$$924  (.A1(net1697),
    .A2(net400),
    .B1(net1689),
    .B2(net666),
    .X(\t$4877 ));
 sky130_fd_sc_hd__xor2_1 \U$$925  (.A(\t$4877 ),
    .B(net1317),
    .X(booth_b12_m48));
 sky130_fd_sc_hd__a22o_1 \U$$926  (.A1(net1687),
    .A2(net395),
    .B1(net1679),
    .B2(net661),
    .X(\t$4878 ));
 sky130_fd_sc_hd__xor2_1 \U$$927  (.A(\t$4878 ),
    .B(net1317),
    .X(booth_b12_m49));
 sky130_fd_sc_hd__a22o_1 \U$$928  (.A1(net1679),
    .A2(net395),
    .B1(net1654),
    .B2(net661),
    .X(\t$4879 ));
 sky130_fd_sc_hd__xor2_1 \U$$929  (.A(\t$4879 ),
    .B(net1317),
    .X(booth_b12_m50));
 sky130_fd_sc_hd__xor2_1 \U$$93  (.A(\t$4453 ),
    .B(net1570),
    .X(booth_b0_m43));
 sky130_fd_sc_hd__a22o_1 \U$$930  (.A1(net1656),
    .A2(net400),
    .B1(net1648),
    .B2(net666),
    .X(\t$4880 ));
 sky130_fd_sc_hd__xor2_1 \U$$931  (.A(\t$4880 ),
    .B(net1317),
    .X(booth_b12_m51));
 sky130_fd_sc_hd__a22o_1 \U$$932  (.A1(net1649),
    .A2(net399),
    .B1(net1641),
    .B2(net665),
    .X(\t$4881 ));
 sky130_fd_sc_hd__xor2_1 \U$$933  (.A(\t$4881 ),
    .B(net1318),
    .X(booth_b12_m52));
 sky130_fd_sc_hd__a22o_1 \U$$934  (.A1(net1641),
    .A2(net399),
    .B1(net1633),
    .B2(net665),
    .X(\t$4882 ));
 sky130_fd_sc_hd__xor2_1 \U$$935  (.A(\t$4882 ),
    .B(net1318),
    .X(booth_b12_m53));
 sky130_fd_sc_hd__a22o_1 \U$$936  (.A1(net1633),
    .A2(net399),
    .B1(net1623),
    .B2(net665),
    .X(\t$4883 ));
 sky130_fd_sc_hd__xor2_1 \U$$937  (.A(\t$4883 ),
    .B(net1318),
    .X(booth_b12_m54));
 sky130_fd_sc_hd__a22o_1 \U$$938  (.A1(net1623),
    .A2(net399),
    .B1(net1615),
    .B2(net665),
    .X(\t$4884 ));
 sky130_fd_sc_hd__xor2_1 \U$$939  (.A(\t$4884 ),
    .B(net1318),
    .X(booth_b12_m55));
 sky130_fd_sc_hd__a22o_1 \U$$94  (.A1(net1729),
    .A2(net445),
    .B1(net1720),
    .B2(net687),
    .X(\t$4454 ));
 sky130_fd_sc_hd__a22o_1 \U$$940  (.A1(net1615),
    .A2(net399),
    .B1(net1607),
    .B2(net665),
    .X(\t$4885 ));
 sky130_fd_sc_hd__xor2_1 \U$$941  (.A(\t$4885 ),
    .B(net1318),
    .X(booth_b12_m56));
 sky130_fd_sc_hd__a22o_1 \U$$942  (.A1(net1607),
    .A2(net399),
    .B1(net1599),
    .B2(net665),
    .X(\t$4886 ));
 sky130_fd_sc_hd__xor2_1 \U$$943  (.A(\t$4886 ),
    .B(net1318),
    .X(booth_b12_m57));
 sky130_fd_sc_hd__a22o_1 \U$$944  (.A1(net1599),
    .A2(net399),
    .B1(net1590),
    .B2(net665),
    .X(\t$4887 ));
 sky130_fd_sc_hd__xor2_1 \U$$945  (.A(\t$4887 ),
    .B(net1318),
    .X(booth_b12_m58));
 sky130_fd_sc_hd__a22o_1 \U$$946  (.A1(net1586),
    .A2(net395),
    .B1(net1578),
    .B2(net661),
    .X(\t$4888 ));
 sky130_fd_sc_hd__xor2_1 \U$$947  (.A(\t$4888 ),
    .B(net1316),
    .X(booth_b12_m59));
 sky130_fd_sc_hd__a22o_1 \U$$948  (.A1(net1581),
    .A2(net395),
    .B1(net1552),
    .B2(net661),
    .X(\t$4889 ));
 sky130_fd_sc_hd__xor2_1 \U$$949  (.A(\t$4889 ),
    .B(net1317),
    .X(booth_b12_m60));
 sky130_fd_sc_hd__xor2_1 \U$$95  (.A(\t$4454 ),
    .B(net1572),
    .X(booth_b0_m44));
 sky130_fd_sc_hd__a22o_1 \U$$950  (.A1(net1551),
    .A2(net395),
    .B1(net1543),
    .B2(net661),
    .X(\t$4890 ));
 sky130_fd_sc_hd__xor2_1 \U$$951  (.A(\t$4890 ),
    .B(net1316),
    .X(booth_b12_m61));
 sky130_fd_sc_hd__a22o_1 \U$$952  (.A1(net1546),
    .A2(net395),
    .B1(net1538),
    .B2(net661),
    .X(\t$4891 ));
 sky130_fd_sc_hd__xor2_1 \U$$953  (.A(\t$4891 ),
    .B(net1316),
    .X(booth_b12_m62));
 sky130_fd_sc_hd__a22o_1 \U$$954  (.A1(net1535),
    .A2(net395),
    .B1(net1527),
    .B2(net661),
    .X(\t$4892 ));
 sky130_fd_sc_hd__xor2_1 \U$$955  (.A(\t$4892 ),
    .B(net1316),
    .X(booth_b12_m63));
 sky130_fd_sc_hd__a22o_1 \U$$956  (.A1(net1530),
    .A2(net395),
    .B1(net1888),
    .B2(net661),
    .X(\t$4893 ));
 sky130_fd_sc_hd__xor2_1 \U$$957  (.A(\t$4893 ),
    .B(net1316),
    .X(booth_b12_m64));
 sky130_fd_sc_hd__inv_1 \U$$958  (.A(net1316),
    .Y(\notsign$4894 ));
 sky130_fd_sc_hd__inv_1 \U$$959  (.A(net1316),
    .Y(\notblock$4895[0] ));
 sky130_fd_sc_hd__a22o_1 \U$$96  (.A1(net1721),
    .A2(net445),
    .B1(net1712),
    .B2(net687),
    .X(\t$4455 ));
 sky130_fd_sc_hd__inv_1 \U$$960  (.A(net6),
    .Y(\notblock$4895[1] ));
 sky130_fd_sc_hd__inv_1 \U$$961  (.A(net1189),
    .Y(\notblock$4895[2] ));
 sky130_fd_sc_hd__and2_1 \U$$962  (.A(net1189),
    .B(\notblock$4895[1] ),
    .X(\t$4896 ));
 sky130_fd_sc_hd__a32o_1 \U$$963  (.A1(\notblock$4895[2] ),
    .A2(net6),
    .A3(net1316),
    .B1(\t$4896 ),
    .B2(\notblock$4895[0] ),
    .X(\sel_0$4897 ));
 sky130_fd_sc_hd__xor2_1 \U$$964  (.A(net6),
    .B(net1317),
    .X(\sel_1$4898 ));
 sky130_fd_sc_hd__a22o_1 \U$$965  (.A1(net1889),
    .A2(net387),
    .B1(net1228),
    .B2(net653),
    .X(\t$4899 ));
 sky130_fd_sc_hd__xor2_1 \U$$966  (.A(\t$4899 ),
    .B(net1185),
    .X(booth_b14_m0));
 sky130_fd_sc_hd__a22o_1 \U$$967  (.A1(net1230),
    .A2(net387),
    .B1(net1123),
    .B2(net653),
    .X(\t$4900 ));
 sky130_fd_sc_hd__xor2_1 \U$$968  (.A(\t$4900 ),
    .B(net1185),
    .X(booth_b14_m1));
 sky130_fd_sc_hd__a22o_1 \U$$969  (.A1(net1123),
    .A2(net385),
    .B1(net1032),
    .B2(net651),
    .X(\t$4901 ));
 sky130_fd_sc_hd__xor2_1 \U$$97  (.A(\t$4455 ),
    .B(net1572),
    .X(booth_b0_m45));
 sky130_fd_sc_hd__xor2_1 \U$$970  (.A(\t$4901 ),
    .B(net1183),
    .X(booth_b14_m2));
 sky130_fd_sc_hd__a22o_1 \U$$971  (.A1(net1032),
    .A2(net385),
    .B1(net933),
    .B2(net651),
    .X(\t$4902 ));
 sky130_fd_sc_hd__xor2_1 \U$$972  (.A(\t$4902 ),
    .B(net1183),
    .X(booth_b14_m3));
 sky130_fd_sc_hd__a22o_1 \U$$973  (.A1(net933),
    .A2(net387),
    .B1(net1672),
    .B2(net653),
    .X(\t$4903 ));
 sky130_fd_sc_hd__xor2_1 \U$$974  (.A(\t$4903 ),
    .B(net1185),
    .X(booth_b14_m4));
 sky130_fd_sc_hd__a22o_1 \U$$975  (.A1(net1676),
    .A2(net389),
    .B1(net1564),
    .B2(net655),
    .X(\t$4904 ));
 sky130_fd_sc_hd__xor2_1 \U$$976  (.A(\t$4904 ),
    .B(net1187),
    .X(booth_b14_m5));
 sky130_fd_sc_hd__a22o_1 \U$$977  (.A1(net1564),
    .A2(net389),
    .B1(net1523),
    .B2(net655),
    .X(\t$4905 ));
 sky130_fd_sc_hd__xor2_1 \U$$978  (.A(\t$4905 ),
    .B(net1187),
    .X(booth_b14_m6));
 sky130_fd_sc_hd__a22o_1 \U$$979  (.A1(net1523),
    .A2(net387),
    .B1(net1515),
    .B2(net653),
    .X(\t$4906 ));
 sky130_fd_sc_hd__a22o_1 \U$$98  (.A1(net1711),
    .A2(net444),
    .B1(net1703),
    .B2(net686),
    .X(\t$4456 ));
 sky130_fd_sc_hd__xor2_1 \U$$980  (.A(\t$4906 ),
    .B(net1187),
    .X(booth_b14_m7));
 sky130_fd_sc_hd__a22o_1 \U$$981  (.A1(net1513),
    .A2(net387),
    .B1(net1505),
    .B2(net653),
    .X(\t$4907 ));
 sky130_fd_sc_hd__xor2_1 \U$$982  (.A(\t$4907 ),
    .B(net1185),
    .X(booth_b14_m8));
 sky130_fd_sc_hd__a22o_1 \U$$983  (.A1(net1505),
    .A2(net387),
    .B1(net1496),
    .B2(net653),
    .X(\t$4908 ));
 sky130_fd_sc_hd__xor2_1 \U$$984  (.A(\t$4908 ),
    .B(net1185),
    .X(booth_b14_m9));
 sky130_fd_sc_hd__a22o_1 \U$$985  (.A1(net1496),
    .A2(net385),
    .B1(net1221),
    .B2(net651),
    .X(\t$4909 ));
 sky130_fd_sc_hd__xor2_1 \U$$986  (.A(\t$4909 ),
    .B(net1183),
    .X(booth_b14_m10));
 sky130_fd_sc_hd__a22o_1 \U$$987  (.A1(net1220),
    .A2(net385),
    .B1(net1210),
    .B2(net651),
    .X(\t$4910 ));
 sky130_fd_sc_hd__xor2_1 \U$$988  (.A(\t$4910 ),
    .B(net1184),
    .X(booth_b14_m11));
 sky130_fd_sc_hd__a22o_1 \U$$989  (.A1(net1210),
    .A2(net385),
    .B1(net1201),
    .B2(net651),
    .X(\t$4911 ));
 sky130_fd_sc_hd__xor2_1 \U$$99  (.A(\t$4456 ),
    .B(net1570),
    .X(booth_b0_m46));
 sky130_fd_sc_hd__xor2_1 \U$$990  (.A(\t$4911 ),
    .B(net1183),
    .X(booth_b14_m12));
 sky130_fd_sc_hd__a22o_1 \U$$991  (.A1(net1201),
    .A2(net385),
    .B1(net1192),
    .B2(net651),
    .X(\t$4912 ));
 sky130_fd_sc_hd__xor2_1 \U$$992  (.A(\t$4912 ),
    .B(net1183),
    .X(booth_b14_m13));
 sky130_fd_sc_hd__a22o_1 \U$$993  (.A1(net1192),
    .A2(net385),
    .B1(net1173),
    .B2(net651),
    .X(\t$4913 ));
 sky130_fd_sc_hd__xor2_1 \U$$994  (.A(\t$4913 ),
    .B(net1183),
    .X(booth_b14_m14));
 sky130_fd_sc_hd__a22o_1 \U$$995  (.A1(net1173),
    .A2(net385),
    .B1(net1164),
    .B2(net651),
    .X(\t$4914 ));
 sky130_fd_sc_hd__xor2_1 \U$$996  (.A(\t$4914 ),
    .B(net1183),
    .X(booth_b14_m15));
 sky130_fd_sc_hd__a22o_1 \U$$997  (.A1(net1164),
    .A2(net385),
    .B1(net1155),
    .B2(net651),
    .X(\t$4915 ));
 sky130_fd_sc_hd__xor2_1 \U$$998  (.A(\t$4915 ),
    .B(net1183),
    .X(booth_b14_m16));
 sky130_fd_sc_hd__a22o_1 \U$$999  (.A1(net1155),
    .A2(net385),
    .B1(net1146),
    .B2(net651),
    .X(\t$4916 ));
 sky130_fd_sc_hd__dfxtp_1 _0168_ (.CLK(clknet_leaf_147_clk),
    .D(booth_b44_m25),
    .Q(pp_row69_20));
 sky130_fd_sc_hd__dfxtp_1 _0169_ (.CLK(clknet_leaf_97_clk),
    .D(booth_b46_m23),
    .Q(pp_row69_21));
 sky130_fd_sc_hd__dfxtp_1 _0170_ (.CLK(clknet_leaf_97_clk),
    .D(booth_b48_m21),
    .Q(pp_row69_22));
 sky130_fd_sc_hd__dfxtp_1 _0171_ (.CLK(clknet_leaf_97_clk),
    .D(booth_b50_m19),
    .Q(pp_row69_23));
 sky130_fd_sc_hd__dfxtp_1 _0172_ (.CLK(clknet_leaf_101_clk),
    .D(booth_b52_m17),
    .Q(pp_row69_24));
 sky130_fd_sc_hd__dfxtp_1 _0173_ (.CLK(clknet_leaf_101_clk),
    .D(booth_b54_m15),
    .Q(pp_row69_25));
 sky130_fd_sc_hd__dfxtp_1 _0174_ (.CLK(clknet_leaf_101_clk),
    .D(booth_b56_m13),
    .Q(pp_row69_26));
 sky130_fd_sc_hd__dfxtp_1 _0175_ (.CLK(clknet_leaf_99_clk),
    .D(booth_b58_m11),
    .Q(pp_row69_27));
 sky130_fd_sc_hd__dfxtp_1 _0176_ (.CLK(clknet_leaf_99_clk),
    .D(booth_b60_m9),
    .Q(pp_row69_28));
 sky130_fd_sc_hd__dfxtp_1 _0177_ (.CLK(clknet_leaf_100_clk),
    .D(booth_b62_m7),
    .Q(pp_row69_29));
 sky130_fd_sc_hd__dfxtp_1 _0178_ (.CLK(clknet_leaf_125_clk),
    .D(booth_b60_m52),
    .Q(pp_row112_7));
 sky130_fd_sc_hd__dfxtp_1 _0179_ (.CLK(clknet_leaf_141_clk),
    .D(booth_b64_m5),
    .Q(pp_row69_30));
 sky130_fd_sc_hd__dfxtp_2 _0180_ (.CLK(clknet_leaf_197_clk),
    .D(net222),
    .Q(pp_row69_31));
 sky130_fd_sc_hd__dfxtp_1 _0181_ (.CLK(clknet_leaf_147_clk),
    .D(booth_b6_m64),
    .Q(pp_row70_1));
 sky130_fd_sc_hd__dfxtp_1 _0182_ (.CLK(clknet_leaf_147_clk),
    .D(booth_b8_m62),
    .Q(pp_row70_2));
 sky130_fd_sc_hd__dfxtp_1 _0183_ (.CLK(clknet_leaf_147_clk),
    .D(booth_b10_m60),
    .Q(pp_row70_3));
 sky130_fd_sc_hd__dfxtp_1 _0184_ (.CLK(clknet_leaf_147_clk),
    .D(booth_b12_m58),
    .Q(pp_row70_4));
 sky130_fd_sc_hd__dfxtp_1 _0185_ (.CLK(clknet_leaf_90_clk),
    .D(booth_b14_m56),
    .Q(pp_row70_5));
 sky130_fd_sc_hd__dfxtp_1 _0186_ (.CLK(clknet_leaf_148_clk),
    .D(booth_b16_m54),
    .Q(pp_row70_6));
 sky130_fd_sc_hd__dfxtp_1 _0187_ (.CLK(clknet_leaf_148_clk),
    .D(booth_b18_m52),
    .Q(pp_row70_7));
 sky130_fd_sc_hd__dfxtp_1 _0188_ (.CLK(clknet_leaf_148_clk),
    .D(booth_b20_m50),
    .Q(pp_row70_8));
 sky130_fd_sc_hd__dfxtp_1 _0189_ (.CLK(clknet_leaf_180_clk),
    .D(booth_b62_m50),
    .Q(pp_row112_8));
 sky130_fd_sc_hd__dfxtp_1 _0190_ (.CLK(clknet_leaf_148_clk),
    .D(booth_b22_m48),
    .Q(pp_row70_9));
 sky130_fd_sc_hd__dfxtp_1 _0191_ (.CLK(clknet_leaf_148_clk),
    .D(booth_b24_m46),
    .Q(pp_row70_10));
 sky130_fd_sc_hd__dfxtp_1 _0192_ (.CLK(clknet_leaf_148_clk),
    .D(booth_b26_m44),
    .Q(pp_row70_11));
 sky130_fd_sc_hd__dfxtp_1 _0193_ (.CLK(clknet_leaf_146_clk),
    .D(booth_b28_m42),
    .Q(pp_row70_12));
 sky130_fd_sc_hd__dfxtp_1 _0194_ (.CLK(clknet_leaf_146_clk),
    .D(booth_b30_m40),
    .Q(pp_row70_13));
 sky130_fd_sc_hd__dfxtp_1 _0195_ (.CLK(clknet_leaf_155_clk),
    .D(booth_b32_m38),
    .Q(pp_row70_14));
 sky130_fd_sc_hd__dfxtp_1 _0196_ (.CLK(clknet_leaf_154_clk),
    .D(booth_b34_m36),
    .Q(pp_row70_15));
 sky130_fd_sc_hd__dfxtp_1 _0197_ (.CLK(clknet_leaf_155_clk),
    .D(booth_b36_m34),
    .Q(pp_row70_16));
 sky130_fd_sc_hd__dfxtp_1 _0198_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b38_m32),
    .Q(pp_row70_17));
 sky130_fd_sc_hd__dfxtp_1 _0199_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b40_m30),
    .Q(pp_row70_18));
 sky130_fd_sc_hd__dfxtp_1 _0200_ (.CLK(clknet_leaf_180_clk),
    .D(booth_b64_m48),
    .Q(pp_row112_9));
 sky130_fd_sc_hd__dfxtp_1 _0201_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b42_m28),
    .Q(pp_row70_19));
 sky130_fd_sc_hd__dfxtp_1 _0202_ (.CLK(clknet_leaf_152_clk),
    .D(booth_b44_m26),
    .Q(pp_row70_20));
 sky130_fd_sc_hd__dfxtp_1 _0203_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b46_m24),
    .Q(pp_row70_21));
 sky130_fd_sc_hd__dfxtp_1 _0204_ (.CLK(clknet_leaf_152_clk),
    .D(booth_b48_m22),
    .Q(pp_row70_22));
 sky130_fd_sc_hd__dfxtp_1 _0205_ (.CLK(clknet_leaf_152_clk),
    .D(booth_b50_m20),
    .Q(pp_row70_23));
 sky130_fd_sc_hd__dfxtp_1 _0206_ (.CLK(clknet_leaf_152_clk),
    .D(booth_b52_m18),
    .Q(pp_row70_24));
 sky130_fd_sc_hd__dfxtp_1 _0207_ (.CLK(clknet_leaf_152_clk),
    .D(booth_b54_m16),
    .Q(pp_row70_25));
 sky130_fd_sc_hd__dfxtp_1 _0208_ (.CLK(clknet_leaf_151_clk),
    .D(booth_b56_m14),
    .Q(pp_row70_26));
 sky130_fd_sc_hd__dfxtp_1 _0209_ (.CLK(clknet_leaf_152_clk),
    .D(booth_b58_m12),
    .Q(pp_row70_27));
 sky130_fd_sc_hd__dfxtp_1 _0210_ (.CLK(clknet_leaf_154_clk),
    .D(booth_b60_m10),
    .Q(pp_row70_28));
 sky130_fd_sc_hd__dfxtp_1 _0211_ (.CLK(clknet_leaf_184_clk),
    .D(net143),
    .Q(pp_row112_10));
 sky130_fd_sc_hd__dfxtp_1 _0212_ (.CLK(clknet_leaf_145_clk),
    .D(booth_b62_m8),
    .Q(pp_row70_29));
 sky130_fd_sc_hd__dfxtp_1 _0213_ (.CLK(clknet_leaf_152_clk),
    .D(booth_b64_m6),
    .Q(pp_row70_30));
 sky130_fd_sc_hd__dfxtp_2 _0214_ (.CLK(clknet_leaf_198_clk),
    .D(net224),
    .Q(pp_row70_31));
 sky130_fd_sc_hd__dfxtp_1 _0215_ (.CLK(clknet_leaf_198_clk),
    .D(\notsign$4684 ),
    .Q(pp_row71_0));
 sky130_fd_sc_hd__dfxtp_1 _0216_ (.CLK(clknet_leaf_198_clk),
    .D(booth_b8_m63),
    .Q(pp_row71_1));
 sky130_fd_sc_hd__dfxtp_1 _0217_ (.CLK(clknet_leaf_198_clk),
    .D(booth_b10_m61),
    .Q(pp_row71_2));
 sky130_fd_sc_hd__dfxtp_1 _0218_ (.CLK(clknet_leaf_199_clk),
    .D(booth_b12_m59),
    .Q(pp_row71_3));
 sky130_fd_sc_hd__dfxtp_1 _0219_ (.CLK(clknet_leaf_200_clk),
    .D(booth_b14_m57),
    .Q(pp_row71_4));
 sky130_fd_sc_hd__dfxtp_1 _0220_ (.CLK(clknet_leaf_199_clk),
    .D(booth_b16_m55),
    .Q(pp_row71_5));
 sky130_fd_sc_hd__dfxtp_1 _0221_ (.CLK(clknet_leaf_200_clk),
    .D(booth_b18_m53),
    .Q(pp_row71_6));
 sky130_fd_sc_hd__dfxtp_1 _0222_ (.CLK(clknet_leaf_126_clk),
    .D(\notsign$6154 ),
    .Q(pp_row113_0));
 sky130_fd_sc_hd__dfxtp_1 _0223_ (.CLK(clknet_leaf_196_clk),
    .D(booth_b20_m51),
    .Q(pp_row71_7));
 sky130_fd_sc_hd__dfxtp_1 _0224_ (.CLK(clknet_leaf_196_clk),
    .D(booth_b22_m49),
    .Q(pp_row71_8));
 sky130_fd_sc_hd__dfxtp_1 _0225_ (.CLK(clknet_leaf_208_clk),
    .D(booth_b24_m47),
    .Q(pp_row71_9));
 sky130_fd_sc_hd__dfxtp_1 _0226_ (.CLK(clknet_leaf_208_clk),
    .D(booth_b26_m45),
    .Q(pp_row71_10));
 sky130_fd_sc_hd__dfxtp_1 _0227_ (.CLK(clknet_leaf_208_clk),
    .D(booth_b28_m43),
    .Q(pp_row71_11));
 sky130_fd_sc_hd__dfxtp_1 _0228_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b30_m41),
    .Q(pp_row71_12));
 sky130_fd_sc_hd__dfxtp_1 _0229_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b32_m39),
    .Q(pp_row71_13));
 sky130_fd_sc_hd__dfxtp_1 _0230_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b34_m37),
    .Q(pp_row71_14));
 sky130_fd_sc_hd__dfxtp_1 _0231_ (.CLK(clknet_leaf_151_clk),
    .D(booth_b36_m35),
    .Q(pp_row71_15));
 sky130_fd_sc_hd__dfxtp_1 _0232_ (.CLK(clknet_leaf_151_clk),
    .D(booth_b38_m33),
    .Q(pp_row71_16));
 sky130_fd_sc_hd__dfxtp_1 _0233_ (.CLK(clknet_leaf_125_clk),
    .D(booth_b50_m63),
    .Q(pp_row113_1));
 sky130_fd_sc_hd__dfxtp_1 _0234_ (.CLK(clknet_leaf_151_clk),
    .D(booth_b40_m31),
    .Q(pp_row71_17));
 sky130_fd_sc_hd__dfxtp_1 _0235_ (.CLK(clknet_leaf_151_clk),
    .D(booth_b42_m29),
    .Q(pp_row71_18));
 sky130_fd_sc_hd__dfxtp_1 _0236_ (.CLK(clknet_leaf_151_clk),
    .D(booth_b44_m27),
    .Q(pp_row71_19));
 sky130_fd_sc_hd__dfxtp_1 _0237_ (.CLK(clknet_leaf_211_clk),
    .D(booth_b46_m25),
    .Q(pp_row71_20));
 sky130_fd_sc_hd__dfxtp_1 _0238_ (.CLK(clknet_leaf_150_clk),
    .D(booth_b48_m23),
    .Q(pp_row71_21));
 sky130_fd_sc_hd__dfxtp_1 _0239_ (.CLK(clknet_leaf_150_clk),
    .D(booth_b50_m21),
    .Q(pp_row71_22));
 sky130_fd_sc_hd__dfxtp_1 _0240_ (.CLK(clknet_leaf_150_clk),
    .D(booth_b52_m19),
    .Q(pp_row71_23));
 sky130_fd_sc_hd__dfxtp_1 _0241_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b54_m17),
    .Q(pp_row71_24));
 sky130_fd_sc_hd__dfxtp_1 _0242_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b56_m15),
    .Q(pp_row71_25));
 sky130_fd_sc_hd__dfxtp_1 _0243_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b58_m13),
    .Q(pp_row71_26));
 sky130_fd_sc_hd__dfxtp_1 _0244_ (.CLK(clknet_leaf_126_clk),
    .D(booth_b52_m61),
    .Q(pp_row113_2));
 sky130_fd_sc_hd__dfxtp_1 _0245_ (.CLK(clknet_leaf_145_clk),
    .D(booth_b60_m11),
    .Q(pp_row71_27));
 sky130_fd_sc_hd__dfxtp_1 _0246_ (.CLK(clknet_leaf_145_clk),
    .D(booth_b62_m9),
    .Q(pp_row71_28));
 sky130_fd_sc_hd__dfxtp_1 _0247_ (.CLK(clknet_leaf_146_clk),
    .D(booth_b64_m7),
    .Q(pp_row71_29));
 sky130_fd_sc_hd__dfxtp_2 _0248_ (.CLK(clknet_leaf_197_clk),
    .D(net225),
    .Q(pp_row71_30));
 sky130_fd_sc_hd__dfxtp_1 _0249_ (.CLK(clknet_leaf_209_clk),
    .D(booth_b8_m64),
    .Q(pp_row72_1));
 sky130_fd_sc_hd__dfxtp_1 _0250_ (.CLK(clknet_leaf_209_clk),
    .D(booth_b10_m62),
    .Q(pp_row72_2));
 sky130_fd_sc_hd__dfxtp_1 _0251_ (.CLK(clknet_leaf_210_clk),
    .D(booth_b12_m60),
    .Q(pp_row72_3));
 sky130_fd_sc_hd__dfxtp_1 _0252_ (.CLK(clknet_leaf_209_clk),
    .D(booth_b14_m58),
    .Q(pp_row72_4));
 sky130_fd_sc_hd__dfxtp_1 _0253_ (.CLK(clknet_leaf_210_clk),
    .D(booth_b16_m56),
    .Q(pp_row72_5));
 sky130_fd_sc_hd__dfxtp_1 _0254_ (.CLK(clknet_leaf_209_clk),
    .D(booth_b18_m54),
    .Q(pp_row72_6));
 sky130_fd_sc_hd__dfxtp_1 _0255_ (.CLK(clknet_leaf_124_clk),
    .D(booth_b54_m59),
    .Q(pp_row113_3));
 sky130_fd_sc_hd__dfxtp_1 _0256_ (.CLK(clknet_leaf_209_clk),
    .D(booth_b20_m52),
    .Q(pp_row72_7));
 sky130_fd_sc_hd__dfxtp_1 _0257_ (.CLK(clknet_leaf_209_clk),
    .D(booth_b22_m50),
    .Q(pp_row72_8));
 sky130_fd_sc_hd__dfxtp_1 _0258_ (.CLK(clknet_leaf_211_clk),
    .D(booth_b24_m48),
    .Q(pp_row72_9));
 sky130_fd_sc_hd__dfxtp_1 _0259_ (.CLK(clknet_leaf_211_clk),
    .D(booth_b26_m46),
    .Q(pp_row72_10));
 sky130_fd_sc_hd__dfxtp_1 _0260_ (.CLK(clknet_leaf_210_clk),
    .D(booth_b28_m44),
    .Q(pp_row72_11));
 sky130_fd_sc_hd__dfxtp_1 _0261_ (.CLK(clknet_leaf_210_clk),
    .D(booth_b30_m42),
    .Q(pp_row72_12));
 sky130_fd_sc_hd__dfxtp_1 _0262_ (.CLK(clknet_leaf_210_clk),
    .D(booth_b32_m40),
    .Q(pp_row72_13));
 sky130_fd_sc_hd__dfxtp_1 _0263_ (.CLK(clknet_leaf_150_clk),
    .D(booth_b34_m38),
    .Q(pp_row72_14));
 sky130_fd_sc_hd__dfxtp_1 _0264_ (.CLK(clknet_leaf_150_clk),
    .D(booth_b36_m36),
    .Q(pp_row72_15));
 sky130_fd_sc_hd__dfxtp_1 _0265_ (.CLK(clknet_leaf_150_clk),
    .D(booth_b38_m34),
    .Q(pp_row72_16));
 sky130_fd_sc_hd__dfxtp_1 _0266_ (.CLK(clknet_leaf_124_clk),
    .D(booth_b56_m57),
    .Q(pp_row113_4));
 sky130_fd_sc_hd__dfxtp_1 _0267_ (.CLK(clknet_leaf_209_clk),
    .D(booth_b40_m32),
    .Q(pp_row72_17));
 sky130_fd_sc_hd__dfxtp_1 _0268_ (.CLK(clknet_leaf_209_clk),
    .D(booth_b42_m30),
    .Q(pp_row72_18));
 sky130_fd_sc_hd__dfxtp_1 _0269_ (.CLK(clknet_leaf_217_clk),
    .D(booth_b44_m28),
    .Q(pp_row72_19));
 sky130_fd_sc_hd__dfxtp_1 _0270_ (.CLK(clknet_leaf_217_clk),
    .D(booth_b46_m26),
    .Q(pp_row72_20));
 sky130_fd_sc_hd__dfxtp_1 _0271_ (.CLK(clknet_leaf_217_clk),
    .D(booth_b48_m24),
    .Q(pp_row72_21));
 sky130_fd_sc_hd__dfxtp_1 _0272_ (.CLK(clknet_leaf_217_clk),
    .D(booth_b50_m22),
    .Q(pp_row72_22));
 sky130_fd_sc_hd__dfxtp_1 _0273_ (.CLK(clknet_leaf_226_clk),
    .D(booth_b52_m20),
    .Q(pp_row72_23));
 sky130_fd_sc_hd__dfxtp_1 _0274_ (.CLK(clknet_leaf_217_clk),
    .D(booth_b54_m18),
    .Q(pp_row72_24));
 sky130_fd_sc_hd__dfxtp_1 _0275_ (.CLK(clknet_leaf_217_clk),
    .D(booth_b56_m16),
    .Q(pp_row72_25));
 sky130_fd_sc_hd__dfxtp_1 _0276_ (.CLK(clknet_leaf_202_clk),
    .D(booth_b58_m14),
    .Q(pp_row72_26));
 sky130_fd_sc_hd__dfxtp_1 _0277_ (.CLK(clknet_leaf_124_clk),
    .D(booth_b58_m55),
    .Q(pp_row113_5));
 sky130_fd_sc_hd__dfxtp_1 _0278_ (.CLK(clknet_leaf_179_clk),
    .D(booth_b64_m61),
    .Q(pp_row125_2));
 sky130_fd_sc_hd__dfxtp_1 _0279_ (.CLK(clknet_leaf_201_clk),
    .D(booth_b60_m12),
    .Q(pp_row72_27));
 sky130_fd_sc_hd__dfxtp_1 _0280_ (.CLK(clknet_leaf_201_clk),
    .D(booth_b62_m10),
    .Q(pp_row72_28));
 sky130_fd_sc_hd__dfxtp_1 _0281_ (.CLK(clknet_leaf_196_clk),
    .D(booth_b64_m8),
    .Q(pp_row72_29));
 sky130_fd_sc_hd__dfxtp_1 _0282_ (.CLK(clknet_leaf_198_clk),
    .D(net226),
    .Q(pp_row72_30));
 sky130_fd_sc_hd__dfxtp_1 _0283_ (.CLK(clknet_leaf_202_clk),
    .D(\notsign$4754 ),
    .Q(pp_row73_0));
 sky130_fd_sc_hd__dfxtp_1 _0284_ (.CLK(clknet_leaf_202_clk),
    .D(booth_b10_m63),
    .Q(pp_row73_1));
 sky130_fd_sc_hd__dfxtp_1 _0285_ (.CLK(clknet_leaf_202_clk),
    .D(booth_b12_m61),
    .Q(pp_row73_2));
 sky130_fd_sc_hd__dfxtp_1 _0286_ (.CLK(clknet_leaf_203_clk),
    .D(booth_b14_m59),
    .Q(pp_row73_3));
 sky130_fd_sc_hd__dfxtp_1 _0287_ (.CLK(clknet_leaf_202_clk),
    .D(booth_b16_m57),
    .Q(pp_row73_4));
 sky130_fd_sc_hd__dfxtp_1 _0288_ (.CLK(clknet_leaf_202_clk),
    .D(booth_b18_m55),
    .Q(pp_row73_5));
 sky130_fd_sc_hd__dfxtp_1 _0289_ (.CLK(clknet_leaf_128_clk),
    .D(booth_b60_m53),
    .Q(pp_row113_6));
 sky130_fd_sc_hd__dfxtp_1 _0290_ (.CLK(clknet_leaf_199_clk),
    .D(booth_b20_m53),
    .Q(pp_row73_6));
 sky130_fd_sc_hd__dfxtp_1 _0291_ (.CLK(clknet_leaf_199_clk),
    .D(booth_b22_m51),
    .Q(pp_row73_7));
 sky130_fd_sc_hd__dfxtp_1 _0292_ (.CLK(clknet_leaf_199_clk),
    .D(booth_b24_m49),
    .Q(pp_row73_8));
 sky130_fd_sc_hd__dfxtp_1 _0293_ (.CLK(clknet_leaf_199_clk),
    .D(booth_b26_m47),
    .Q(pp_row73_9));
 sky130_fd_sc_hd__dfxtp_1 _0294_ (.CLK(clknet_leaf_199_clk),
    .D(booth_b28_m45),
    .Q(pp_row73_10));
 sky130_fd_sc_hd__dfxtp_1 _0295_ (.CLK(clknet_leaf_199_clk),
    .D(booth_b30_m43),
    .Q(pp_row73_11));
 sky130_fd_sc_hd__dfxtp_1 _0296_ (.CLK(clknet_leaf_201_clk),
    .D(booth_b32_m41),
    .Q(pp_row73_12));
 sky130_fd_sc_hd__dfxtp_1 _0297_ (.CLK(clknet_leaf_201_clk),
    .D(booth_b34_m39),
    .Q(pp_row73_13));
 sky130_fd_sc_hd__dfxtp_1 _0298_ (.CLK(clknet_leaf_201_clk),
    .D(booth_b36_m37),
    .Q(pp_row73_14));
 sky130_fd_sc_hd__dfxtp_1 _0299_ (.CLK(clknet_leaf_226_clk),
    .D(booth_b38_m35),
    .Q(pp_row73_15));
 sky130_fd_sc_hd__dfxtp_1 _0300_ (.CLK(clknet_leaf_128_clk),
    .D(booth_b62_m51),
    .Q(pp_row113_7));
 sky130_fd_sc_hd__dfxtp_1 _0301_ (.CLK(clknet_leaf_227_clk),
    .D(booth_b40_m33),
    .Q(pp_row73_16));
 sky130_fd_sc_hd__dfxtp_1 _0302_ (.CLK(clknet_leaf_227_clk),
    .D(booth_b42_m31),
    .Q(pp_row73_17));
 sky130_fd_sc_hd__dfxtp_1 _0303_ (.CLK(clknet_leaf_227_clk),
    .D(booth_b44_m29),
    .Q(pp_row73_18));
 sky130_fd_sc_hd__dfxtp_1 _0304_ (.CLK(clknet_leaf_225_clk),
    .D(booth_b46_m27),
    .Q(pp_row73_19));
 sky130_fd_sc_hd__dfxtp_1 _0305_ (.CLK(clknet_leaf_225_clk),
    .D(booth_b48_m25),
    .Q(pp_row73_20));
 sky130_fd_sc_hd__dfxtp_1 _0306_ (.CLK(clknet_leaf_226_clk),
    .D(booth_b50_m23),
    .Q(pp_row73_21));
 sky130_fd_sc_hd__dfxtp_1 _0307_ (.CLK(clknet_leaf_226_clk),
    .D(booth_b52_m21),
    .Q(pp_row73_22));
 sky130_fd_sc_hd__dfxtp_1 _0308_ (.CLK(clknet_leaf_226_clk),
    .D(booth_b54_m19),
    .Q(pp_row73_23));
 sky130_fd_sc_hd__dfxtp_1 _0309_ (.CLK(clknet_leaf_209_clk),
    .D(booth_b56_m17),
    .Q(pp_row73_24));
 sky130_fd_sc_hd__dfxtp_1 _0310_ (.CLK(clknet_leaf_202_clk),
    .D(booth_b58_m15),
    .Q(pp_row73_25));
 sky130_fd_sc_hd__dfxtp_1 _0311_ (.CLK(clknet_leaf_128_clk),
    .D(booth_b64_m49),
    .Q(pp_row113_8));
 sky130_fd_sc_hd__dfxtp_1 _0312_ (.CLK(clknet_leaf_202_clk),
    .D(booth_b60_m13),
    .Q(pp_row73_26));
 sky130_fd_sc_hd__dfxtp_1 _0313_ (.CLK(clknet_leaf_201_clk),
    .D(booth_b62_m11),
    .Q(pp_row73_27));
 sky130_fd_sc_hd__dfxtp_1 _0314_ (.CLK(clknet_leaf_200_clk),
    .D(booth_b64_m9),
    .Q(pp_row73_28));
 sky130_fd_sc_hd__dfxtp_1 _0315_ (.CLK(clknet_leaf_197_clk),
    .D(net227),
    .Q(pp_row73_29));
 sky130_fd_sc_hd__dfxtp_1 _0316_ (.CLK(clknet_leaf_196_clk),
    .D(booth_b10_m64),
    .Q(pp_row74_1));
 sky130_fd_sc_hd__dfxtp_1 _0317_ (.CLK(clknet_leaf_196_clk),
    .D(booth_b12_m62),
    .Q(pp_row74_2));
 sky130_fd_sc_hd__dfxtp_1 _0318_ (.CLK(clknet_leaf_200_clk),
    .D(booth_b14_m60),
    .Q(pp_row74_3));
 sky130_fd_sc_hd__dfxtp_1 _0319_ (.CLK(clknet_leaf_200_clk),
    .D(booth_b16_m58),
    .Q(pp_row74_4));
 sky130_fd_sc_hd__dfxtp_1 _0320_ (.CLK(clknet_leaf_200_clk),
    .D(booth_b18_m56),
    .Q(pp_row74_5));
 sky130_fd_sc_hd__dfxtp_1 _0321_ (.CLK(clknet_leaf_200_clk),
    .D(booth_b20_m54),
    .Q(pp_row74_6));
 sky130_fd_sc_hd__dfxtp_2 _0322_ (.CLK(clknet_leaf_182_clk),
    .D(net144),
    .Q(pp_row113_9));
 sky130_fd_sc_hd__dfxtp_1 _0323_ (.CLK(clknet_leaf_201_clk),
    .D(booth_b22_m52),
    .Q(pp_row74_7));
 sky130_fd_sc_hd__dfxtp_1 _0324_ (.CLK(clknet_leaf_199_clk),
    .D(booth_b24_m50),
    .Q(pp_row74_8));
 sky130_fd_sc_hd__dfxtp_1 _0325_ (.CLK(clknet_leaf_199_clk),
    .D(booth_b26_m48),
    .Q(pp_row74_9));
 sky130_fd_sc_hd__dfxtp_1 _0326_ (.CLK(clknet_leaf_201_clk),
    .D(booth_b28_m46),
    .Q(pp_row74_10));
 sky130_fd_sc_hd__dfxtp_1 _0327_ (.CLK(clknet_leaf_227_clk),
    .D(booth_b30_m44),
    .Q(pp_row74_11));
 sky130_fd_sc_hd__dfxtp_1 _0328_ (.CLK(clknet_leaf_227_clk),
    .D(booth_b32_m42),
    .Q(pp_row74_12));
 sky130_fd_sc_hd__dfxtp_1 _0329_ (.CLK(clknet_leaf_201_clk),
    .D(booth_b34_m40),
    .Q(pp_row74_13));
 sky130_fd_sc_hd__dfxtp_1 _0330_ (.CLK(clknet_leaf_224_clk),
    .D(booth_b36_m38),
    .Q(pp_row74_14));
 sky130_fd_sc_hd__dfxtp_1 _0331_ (.CLK(clknet_leaf_224_clk),
    .D(booth_b38_m36),
    .Q(pp_row74_15));
 sky130_fd_sc_hd__dfxtp_1 _0332_ (.CLK(clknet_leaf_224_clk),
    .D(booth_b40_m34),
    .Q(pp_row74_16));
 sky130_fd_sc_hd__dfxtp_1 _0333_ (.CLK(clknet_leaf_128_clk),
    .D(booth_b50_m64),
    .Q(pp_row114_1));
 sky130_fd_sc_hd__dfxtp_1 _0334_ (.CLK(clknet_leaf_225_clk),
    .D(booth_b42_m32),
    .Q(pp_row74_17));
 sky130_fd_sc_hd__dfxtp_1 _0335_ (.CLK(clknet_leaf_225_clk),
    .D(booth_b44_m30),
    .Q(pp_row74_18));
 sky130_fd_sc_hd__dfxtp_1 _0336_ (.CLK(clknet_leaf_225_clk),
    .D(booth_b46_m28),
    .Q(pp_row74_19));
 sky130_fd_sc_hd__dfxtp_1 _0337_ (.CLK(clknet_leaf_226_clk),
    .D(booth_b48_m26),
    .Q(pp_row74_20));
 sky130_fd_sc_hd__dfxtp_1 _0338_ (.CLK(clknet_leaf_225_clk),
    .D(booth_b50_m24),
    .Q(pp_row74_21));
 sky130_fd_sc_hd__dfxtp_1 _0339_ (.CLK(clknet_leaf_226_clk),
    .D(booth_b52_m22),
    .Q(pp_row74_22));
 sky130_fd_sc_hd__dfxtp_1 _0340_ (.CLK(clknet_leaf_202_clk),
    .D(booth_b54_m20),
    .Q(pp_row74_23));
 sky130_fd_sc_hd__dfxtp_1 _0341_ (.CLK(clknet_leaf_202_clk),
    .D(booth_b56_m18),
    .Q(pp_row74_24));
 sky130_fd_sc_hd__dfxtp_1 _0342_ (.CLK(clknet_leaf_202_clk),
    .D(booth_b58_m16),
    .Q(pp_row74_25));
 sky130_fd_sc_hd__dfxtp_1 _0343_ (.CLK(clknet_leaf_203_clk),
    .D(booth_b60_m14),
    .Q(pp_row74_26));
 sky130_fd_sc_hd__dfxtp_1 _0344_ (.CLK(clknet_leaf_129_clk),
    .D(booth_b52_m62),
    .Q(pp_row114_2));
 sky130_fd_sc_hd__dfxtp_1 _0345_ (.CLK(clknet_leaf_203_clk),
    .D(booth_b62_m12),
    .Q(pp_row74_27));
 sky130_fd_sc_hd__dfxtp_1 _0346_ (.CLK(clknet_leaf_203_clk),
    .D(booth_b64_m10),
    .Q(pp_row74_28));
 sky130_fd_sc_hd__dfxtp_1 _0347_ (.CLK(clknet_leaf_197_clk),
    .D(net228),
    .Q(pp_row74_29));
 sky130_fd_sc_hd__dfxtp_1 _0348_ (.CLK(clknet_leaf_203_clk),
    .D(\notsign$4824 ),
    .Q(pp_row75_0));
 sky130_fd_sc_hd__dfxtp_1 _0349_ (.CLK(clknet_leaf_200_clk),
    .D(booth_b12_m63),
    .Q(pp_row75_1));
 sky130_fd_sc_hd__dfxtp_1 _0350_ (.CLK(clknet_leaf_200_clk),
    .D(booth_b14_m61),
    .Q(pp_row75_2));
 sky130_fd_sc_hd__dfxtp_1 _0351_ (.CLK(clknet_leaf_200_clk),
    .D(booth_b16_m59),
    .Q(pp_row75_3));
 sky130_fd_sc_hd__dfxtp_1 _0352_ (.CLK(clknet_leaf_200_clk),
    .D(booth_b18_m57),
    .Q(pp_row75_4));
 sky130_fd_sc_hd__dfxtp_1 _0353_ (.CLK(clknet_leaf_200_clk),
    .D(booth_b20_m55),
    .Q(pp_row75_5));
 sky130_fd_sc_hd__dfxtp_1 _0354_ (.CLK(clknet_leaf_196_clk),
    .D(booth_b22_m53),
    .Q(pp_row75_6));
 sky130_fd_sc_hd__dfxtp_1 _0355_ (.CLK(clknet_leaf_125_clk),
    .D(booth_b54_m60),
    .Q(pp_row114_3));
 sky130_fd_sc_hd__dfxtp_1 _0356_ (.CLK(clknet_leaf_196_clk),
    .D(booth_b24_m51),
    .Q(pp_row75_7));
 sky130_fd_sc_hd__dfxtp_1 _0357_ (.CLK(clknet_leaf_196_clk),
    .D(booth_b26_m49),
    .Q(pp_row75_8));
 sky130_fd_sc_hd__dfxtp_1 _0358_ (.CLK(clknet_leaf_192_clk),
    .D(booth_b28_m47),
    .Q(pp_row75_9));
 sky130_fd_sc_hd__dfxtp_1 _0359_ (.CLK(clknet_leaf_192_clk),
    .D(booth_b30_m45),
    .Q(pp_row75_10));
 sky130_fd_sc_hd__dfxtp_1 _0360_ (.CLK(clknet_leaf_192_clk),
    .D(booth_b32_m43),
    .Q(pp_row75_11));
 sky130_fd_sc_hd__dfxtp_1 _0361_ (.CLK(clknet_leaf_204_clk),
    .D(booth_b34_m41),
    .Q(pp_row75_12));
 sky130_fd_sc_hd__dfxtp_1 _0362_ (.CLK(clknet_leaf_192_clk),
    .D(booth_b36_m39),
    .Q(pp_row75_13));
 sky130_fd_sc_hd__dfxtp_1 _0363_ (.CLK(clknet_leaf_204_clk),
    .D(booth_b38_m37),
    .Q(pp_row75_14));
 sky130_fd_sc_hd__dfxtp_1 _0364_ (.CLK(clknet_leaf_204_clk),
    .D(booth_b40_m35),
    .Q(pp_row75_15));
 sky130_fd_sc_hd__dfxtp_1 _0365_ (.CLK(clknet_leaf_204_clk),
    .D(booth_b42_m33),
    .Q(pp_row75_16));
 sky130_fd_sc_hd__dfxtp_1 _0366_ (.CLK(clknet_leaf_125_clk),
    .D(booth_b56_m58),
    .Q(pp_row114_4));
 sky130_fd_sc_hd__dfxtp_1 _0367_ (.CLK(clknet_leaf_190_clk),
    .D(booth_b44_m31),
    .Q(pp_row75_17));
 sky130_fd_sc_hd__dfxtp_1 _0368_ (.CLK(clknet_leaf_205_clk),
    .D(booth_b46_m29),
    .Q(pp_row75_18));
 sky130_fd_sc_hd__dfxtp_1 _0369_ (.CLK(clknet_leaf_205_clk),
    .D(booth_b48_m27),
    .Q(pp_row75_19));
 sky130_fd_sc_hd__dfxtp_1 _0370_ (.CLK(clknet_leaf_205_clk),
    .D(booth_b50_m25),
    .Q(pp_row75_20));
 sky130_fd_sc_hd__dfxtp_1 _0371_ (.CLK(clknet_leaf_203_clk),
    .D(booth_b52_m23),
    .Q(pp_row75_21));
 sky130_fd_sc_hd__dfxtp_1 _0372_ (.CLK(clknet_leaf_203_clk),
    .D(booth_b54_m21),
    .Q(pp_row75_22));
 sky130_fd_sc_hd__dfxtp_1 _0373_ (.CLK(clknet_leaf_204_clk),
    .D(booth_b56_m19),
    .Q(pp_row75_23));
 sky130_fd_sc_hd__dfxtp_1 _0374_ (.CLK(clknet_leaf_204_clk),
    .D(booth_b58_m17),
    .Q(pp_row75_24));
 sky130_fd_sc_hd__dfxtp_1 _0375_ (.CLK(clknet_leaf_203_clk),
    .D(booth_b60_m15),
    .Q(pp_row75_25));
 sky130_fd_sc_hd__dfxtp_1 _0376_ (.CLK(clknet_leaf_203_clk),
    .D(booth_b62_m13),
    .Q(pp_row75_26));
 sky130_fd_sc_hd__dfxtp_1 _0377_ (.CLK(clknet_leaf_126_clk),
    .D(booth_b58_m56),
    .Q(pp_row114_5));
 sky130_fd_sc_hd__dfxtp_1 _0378_ (.CLK(clknet_leaf_200_clk),
    .D(booth_b64_m11),
    .Q(pp_row75_27));
 sky130_fd_sc_hd__dfxtp_1 _0379_ (.CLK(clknet_leaf_197_clk),
    .D(net229),
    .Q(pp_row75_28));
 sky130_fd_sc_hd__dfxtp_1 _0380_ (.CLK(clknet_leaf_204_clk),
    .D(booth_b12_m64),
    .Q(pp_row76_1));
 sky130_fd_sc_hd__dfxtp_1 _0381_ (.CLK(clknet_leaf_204_clk),
    .D(booth_b14_m62),
    .Q(pp_row76_2));
 sky130_fd_sc_hd__dfxtp_1 _0382_ (.CLK(clknet_leaf_204_clk),
    .D(booth_b16_m60),
    .Q(pp_row76_3));
 sky130_fd_sc_hd__dfxtp_1 _0383_ (.CLK(clknet_leaf_204_clk),
    .D(booth_b18_m58),
    .Q(pp_row76_4));
 sky130_fd_sc_hd__dfxtp_1 _0384_ (.CLK(clknet_leaf_193_clk),
    .D(booth_b20_m56),
    .Q(pp_row76_5));
 sky130_fd_sc_hd__dfxtp_1 _0385_ (.CLK(clknet_leaf_195_clk),
    .D(booth_b22_m54),
    .Q(pp_row76_6));
 sky130_fd_sc_hd__dfxtp_1 _0386_ (.CLK(clknet_leaf_195_clk),
    .D(booth_b24_m52),
    .Q(pp_row76_7));
 sky130_fd_sc_hd__dfxtp_1 _0387_ (.CLK(clknet_leaf_196_clk),
    .D(booth_b26_m50),
    .Q(pp_row76_8));
 sky130_fd_sc_hd__dfxtp_1 _0388_ (.CLK(clknet_leaf_127_clk),
    .D(booth_b60_m54),
    .Q(pp_row114_6));
 sky130_fd_sc_hd__dfxtp_2 _0389_ (.CLK(clknet_leaf_181_clk),
    .D(net157),
    .Q(pp_row125_3));
 sky130_fd_sc_hd__dfxtp_1 _0390_ (.CLK(clknet_leaf_196_clk),
    .D(booth_b28_m48),
    .Q(pp_row76_9));
 sky130_fd_sc_hd__dfxtp_1 _0391_ (.CLK(clknet_leaf_196_clk),
    .D(booth_b30_m46),
    .Q(pp_row76_10));
 sky130_fd_sc_hd__dfxtp_1 _0392_ (.CLK(clknet_leaf_191_clk),
    .D(booth_b32_m44),
    .Q(pp_row76_11));
 sky130_fd_sc_hd__dfxtp_1 _0393_ (.CLK(clknet_leaf_191_clk),
    .D(booth_b34_m42),
    .Q(pp_row76_12));
 sky130_fd_sc_hd__dfxtp_1 _0394_ (.CLK(clknet_leaf_191_clk),
    .D(booth_b36_m40),
    .Q(pp_row76_13));
 sky130_fd_sc_hd__dfxtp_1 _0395_ (.CLK(clknet_leaf_192_clk),
    .D(booth_b38_m38),
    .Q(pp_row76_14));
 sky130_fd_sc_hd__dfxtp_1 _0396_ (.CLK(clknet_leaf_191_clk),
    .D(booth_b40_m36),
    .Q(pp_row76_15));
 sky130_fd_sc_hd__dfxtp_1 _0397_ (.CLK(clknet_leaf_191_clk),
    .D(booth_b42_m34),
    .Q(pp_row76_16));
 sky130_fd_sc_hd__dfxtp_1 _0398_ (.CLK(clknet_leaf_190_clk),
    .D(booth_b44_m32),
    .Q(pp_row76_17));
 sky130_fd_sc_hd__dfxtp_1 _0399_ (.CLK(clknet_leaf_191_clk),
    .D(booth_b46_m30),
    .Q(pp_row76_18));
 sky130_fd_sc_hd__dfxtp_1 _0400_ (.CLK(clknet_leaf_127_clk),
    .D(booth_b62_m52),
    .Q(pp_row114_7));
 sky130_fd_sc_hd__dfxtp_1 _0401_ (.CLK(clknet_leaf_190_clk),
    .D(booth_b48_m28),
    .Q(pp_row76_19));
 sky130_fd_sc_hd__dfxtp_1 _0402_ (.CLK(clknet_leaf_208_clk),
    .D(booth_b50_m26),
    .Q(pp_row76_20));
 sky130_fd_sc_hd__dfxtp_1 _0403_ (.CLK(clknet_leaf_208_clk),
    .D(booth_b52_m24),
    .Q(pp_row76_21));
 sky130_fd_sc_hd__dfxtp_1 _0404_ (.CLK(clknet_leaf_208_clk),
    .D(booth_b54_m22),
    .Q(pp_row76_22));
 sky130_fd_sc_hd__dfxtp_1 _0405_ (.CLK(clknet_leaf_205_clk),
    .D(booth_b56_m20),
    .Q(pp_row76_23));
 sky130_fd_sc_hd__dfxtp_1 _0406_ (.CLK(clknet_leaf_206_clk),
    .D(booth_b58_m18),
    .Q(pp_row76_24));
 sky130_fd_sc_hd__dfxtp_1 _0407_ (.CLK(clknet_leaf_205_clk),
    .D(booth_b60_m16),
    .Q(pp_row76_25));
 sky130_fd_sc_hd__dfxtp_1 _0408_ (.CLK(clknet_leaf_206_clk),
    .D(booth_b62_m14),
    .Q(pp_row76_26));
 sky130_fd_sc_hd__dfxtp_1 _0409_ (.CLK(clknet_leaf_208_clk),
    .D(booth_b64_m12),
    .Q(pp_row76_27));
 sky130_fd_sc_hd__dfxtp_1 _0410_ (.CLK(clknet_leaf_197_clk),
    .D(net230),
    .Q(pp_row76_28));
 sky130_fd_sc_hd__dfxtp_1 _0411_ (.CLK(clknet_leaf_125_clk),
    .D(booth_b64_m50),
    .Q(pp_row114_8));
 sky130_fd_sc_hd__dfxtp_1 _0412_ (.CLK(clknet_leaf_192_clk),
    .D(\notsign$4894 ),
    .Q(pp_row77_0));
 sky130_fd_sc_hd__dfxtp_1 _0413_ (.CLK(clknet_leaf_192_clk),
    .D(booth_b14_m63),
    .Q(pp_row77_1));
 sky130_fd_sc_hd__dfxtp_1 _0414_ (.CLK(clknet_leaf_193_clk),
    .D(booth_b16_m61),
    .Q(pp_row77_2));
 sky130_fd_sc_hd__dfxtp_1 _0415_ (.CLK(clknet_leaf_155_clk),
    .D(booth_b18_m59),
    .Q(pp_row77_3));
 sky130_fd_sc_hd__dfxtp_1 _0416_ (.CLK(clknet_leaf_155_clk),
    .D(booth_b20_m57),
    .Q(pp_row77_4));
 sky130_fd_sc_hd__dfxtp_1 _0417_ (.CLK(clknet_leaf_155_clk),
    .D(booth_b22_m55),
    .Q(pp_row77_5));
 sky130_fd_sc_hd__dfxtp_1 _0418_ (.CLK(clknet_leaf_145_clk),
    .D(booth_b24_m53),
    .Q(pp_row77_6));
 sky130_fd_sc_hd__dfxtp_1 _0419_ (.CLK(clknet_leaf_145_clk),
    .D(booth_b26_m51),
    .Q(pp_row77_7));
 sky130_fd_sc_hd__dfxtp_1 _0420_ (.CLK(clknet_leaf_145_clk),
    .D(booth_b28_m49),
    .Q(pp_row77_8));
 sky130_fd_sc_hd__dfxtp_1 _0421_ (.CLK(clknet_leaf_207_clk),
    .D(booth_b30_m47),
    .Q(pp_row77_9));
 sky130_fd_sc_hd__dfxtp_2 _0422_ (.CLK(clknet_leaf_181_clk),
    .D(net145),
    .Q(pp_row114_9));
 sky130_fd_sc_hd__dfxtp_1 _0423_ (.CLK(clknet_leaf_207_clk),
    .D(booth_b32_m45),
    .Q(pp_row77_10));
 sky130_fd_sc_hd__dfxtp_1 _0424_ (.CLK(clknet_leaf_211_clk),
    .D(booth_b34_m43),
    .Q(pp_row77_11));
 sky130_fd_sc_hd__dfxtp_1 _0425_ (.CLK(clknet_leaf_207_clk),
    .D(booth_b36_m41),
    .Q(pp_row77_12));
 sky130_fd_sc_hd__dfxtp_1 _0426_ (.CLK(clknet_leaf_207_clk),
    .D(booth_b38_m39),
    .Q(pp_row77_13));
 sky130_fd_sc_hd__dfxtp_1 _0427_ (.CLK(clknet_leaf_207_clk),
    .D(booth_b40_m37),
    .Q(pp_row77_14));
 sky130_fd_sc_hd__dfxtp_1 _0428_ (.CLK(clknet_leaf_207_clk),
    .D(booth_b42_m35),
    .Q(pp_row77_15));
 sky130_fd_sc_hd__dfxtp_1 _0429_ (.CLK(clknet_leaf_207_clk),
    .D(booth_b44_m33),
    .Q(pp_row77_16));
 sky130_fd_sc_hd__dfxtp_1 _0430_ (.CLK(clknet_leaf_207_clk),
    .D(booth_b46_m31),
    .Q(pp_row77_17));
 sky130_fd_sc_hd__dfxtp_1 _0431_ (.CLK(clknet_leaf_154_clk),
    .D(booth_b48_m29),
    .Q(pp_row77_18));
 sky130_fd_sc_hd__dfxtp_1 _0432_ (.CLK(clknet_leaf_154_clk),
    .D(booth_b50_m27),
    .Q(pp_row77_19));
 sky130_fd_sc_hd__dfxtp_1 _0433_ (.CLK(clknet_leaf_131_clk),
    .D(\notsign$6224 ),
    .Q(pp_row115_0));
 sky130_fd_sc_hd__dfxtp_1 _0434_ (.CLK(clknet_leaf_154_clk),
    .D(booth_b52_m25),
    .Q(pp_row77_20));
 sky130_fd_sc_hd__dfxtp_1 _0435_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b54_m23),
    .Q(pp_row77_21));
 sky130_fd_sc_hd__dfxtp_1 _0436_ (.CLK(clknet_leaf_154_clk),
    .D(booth_b56_m21),
    .Q(pp_row77_22));
 sky130_fd_sc_hd__dfxtp_1 _0437_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b58_m19),
    .Q(pp_row77_23));
 sky130_fd_sc_hd__dfxtp_1 _0438_ (.CLK(clknet_leaf_160_clk),
    .D(booth_b60_m17),
    .Q(pp_row77_24));
 sky130_fd_sc_hd__dfxtp_1 _0439_ (.CLK(clknet_leaf_154_clk),
    .D(booth_b62_m15),
    .Q(pp_row77_25));
 sky130_fd_sc_hd__dfxtp_1 _0440_ (.CLK(clknet_leaf_161_clk),
    .D(booth_b64_m13),
    .Q(pp_row77_26));
 sky130_fd_sc_hd__dfxtp_1 _0441_ (.CLK(clknet_leaf_197_clk),
    .D(net231),
    .Q(pp_row77_27));
 sky130_fd_sc_hd__dfxtp_1 _0442_ (.CLK(clknet_leaf_151_clk),
    .D(booth_b14_m64),
    .Q(pp_row78_1));
 sky130_fd_sc_hd__dfxtp_1 _0443_ (.CLK(clknet_leaf_155_clk),
    .D(booth_b16_m62),
    .Q(pp_row78_2));
 sky130_fd_sc_hd__dfxtp_1 _0444_ (.CLK(clknet_leaf_131_clk),
    .D(booth_b52_m63),
    .Q(pp_row115_1));
 sky130_fd_sc_hd__dfxtp_1 _0445_ (.CLK(clknet_leaf_207_clk),
    .D(booth_b18_m60),
    .Q(pp_row78_3));
 sky130_fd_sc_hd__dfxtp_1 _0446_ (.CLK(clknet_leaf_207_clk),
    .D(booth_b20_m58),
    .Q(pp_row78_4));
 sky130_fd_sc_hd__dfxtp_1 _0447_ (.CLK(clknet_leaf_206_clk),
    .D(booth_b22_m56),
    .Q(pp_row78_5));
 sky130_fd_sc_hd__dfxtp_1 _0448_ (.CLK(clknet_leaf_206_clk),
    .D(booth_b24_m54),
    .Q(pp_row78_6));
 sky130_fd_sc_hd__dfxtp_1 _0449_ (.CLK(clknet_leaf_206_clk),
    .D(booth_b26_m52),
    .Q(pp_row78_7));
 sky130_fd_sc_hd__dfxtp_1 _0450_ (.CLK(clknet_leaf_158_clk),
    .D(booth_b28_m50),
    .Q(pp_row78_8));
 sky130_fd_sc_hd__dfxtp_1 _0451_ (.CLK(clknet_leaf_158_clk),
    .D(booth_b30_m48),
    .Q(pp_row78_9));
 sky130_fd_sc_hd__dfxtp_1 _0452_ (.CLK(clknet_leaf_158_clk),
    .D(booth_b32_m46),
    .Q(pp_row78_10));
 sky130_fd_sc_hd__dfxtp_1 _0453_ (.CLK(clknet_leaf_158_clk),
    .D(booth_b34_m44),
    .Q(pp_row78_11));
 sky130_fd_sc_hd__dfxtp_1 _0454_ (.CLK(clknet_leaf_158_clk),
    .D(booth_b36_m42),
    .Q(pp_row78_12));
 sky130_fd_sc_hd__dfxtp_1 _0455_ (.CLK(clknet_leaf_131_clk),
    .D(booth_b54_m61),
    .Q(pp_row115_2));
 sky130_fd_sc_hd__dfxtp_1 _0456_ (.CLK(clknet_leaf_158_clk),
    .D(booth_b38_m40),
    .Q(pp_row78_13));
 sky130_fd_sc_hd__dfxtp_1 _0457_ (.CLK(clknet_leaf_157_clk),
    .D(booth_b40_m38),
    .Q(pp_row78_14));
 sky130_fd_sc_hd__dfxtp_1 _0458_ (.CLK(clknet_leaf_157_clk),
    .D(booth_b42_m36),
    .Q(pp_row78_15));
 sky130_fd_sc_hd__dfxtp_1 _0459_ (.CLK(clknet_leaf_157_clk),
    .D(booth_b44_m34),
    .Q(pp_row78_16));
 sky130_fd_sc_hd__dfxtp_1 _0460_ (.CLK(clknet_leaf_157_clk),
    .D(booth_b46_m32),
    .Q(pp_row78_17));
 sky130_fd_sc_hd__dfxtp_1 _0461_ (.CLK(clknet_leaf_157_clk),
    .D(booth_b48_m30),
    .Q(pp_row78_18));
 sky130_fd_sc_hd__dfxtp_1 _0462_ (.CLK(clknet_leaf_157_clk),
    .D(booth_b50_m28),
    .Q(pp_row78_19));
 sky130_fd_sc_hd__dfxtp_1 _0463_ (.CLK(clknet_leaf_206_clk),
    .D(booth_b52_m26),
    .Q(pp_row78_20));
 sky130_fd_sc_hd__dfxtp_1 _0464_ (.CLK(clknet_leaf_206_clk),
    .D(booth_b54_m24),
    .Q(pp_row78_21));
 sky130_fd_sc_hd__dfxtp_1 _0465_ (.CLK(clknet_leaf_205_clk),
    .D(booth_b56_m22),
    .Q(pp_row78_22));
 sky130_fd_sc_hd__dfxtp_1 _0466_ (.CLK(clknet_leaf_130_clk),
    .D(booth_b56_m59),
    .Q(pp_row115_3));
 sky130_fd_sc_hd__dfxtp_1 _0467_ (.CLK(clknet_leaf_155_clk),
    .D(booth_b58_m20),
    .Q(pp_row78_23));
 sky130_fd_sc_hd__dfxtp_1 _0468_ (.CLK(clknet_leaf_155_clk),
    .D(booth_b60_m18),
    .Q(pp_row78_24));
 sky130_fd_sc_hd__dfxtp_1 _0469_ (.CLK(clknet_leaf_155_clk),
    .D(booth_b62_m16),
    .Q(pp_row78_25));
 sky130_fd_sc_hd__dfxtp_1 _0470_ (.CLK(clknet_leaf_192_clk),
    .D(booth_b64_m14),
    .Q(pp_row78_26));
 sky130_fd_sc_hd__dfxtp_1 _0471_ (.CLK(clknet_leaf_197_clk),
    .D(net232),
    .Q(pp_row78_27));
 sky130_fd_sc_hd__dfxtp_1 _0472_ (.CLK(clknet_leaf_193_clk),
    .D(\notsign$4964 ),
    .Q(pp_row79_0));
 sky130_fd_sc_hd__dfxtp_1 _0473_ (.CLK(clknet_leaf_193_clk),
    .D(booth_b16_m63),
    .Q(pp_row79_1));
 sky130_fd_sc_hd__dfxtp_1 _0474_ (.CLK(clknet_leaf_193_clk),
    .D(booth_b18_m61),
    .Q(pp_row79_2));
 sky130_fd_sc_hd__dfxtp_1 _0475_ (.CLK(clknet_leaf_186_clk),
    .D(booth_b20_m59),
    .Q(pp_row79_3));
 sky130_fd_sc_hd__dfxtp_1 _0476_ (.CLK(clknet_leaf_193_clk),
    .D(booth_b22_m57),
    .Q(pp_row79_4));
 sky130_fd_sc_hd__dfxtp_1 _0477_ (.CLK(clknet_leaf_129_clk),
    .D(booth_b58_m57),
    .Q(pp_row115_4));
 sky130_fd_sc_hd__dfxtp_1 _0478_ (.CLK(clknet_leaf_193_clk),
    .D(booth_b24_m55),
    .Q(pp_row79_5));
 sky130_fd_sc_hd__dfxtp_1 _0479_ (.CLK(clknet_leaf_205_clk),
    .D(booth_b26_m53),
    .Q(pp_row79_6));
 sky130_fd_sc_hd__dfxtp_1 _0480_ (.CLK(clknet_leaf_205_clk),
    .D(booth_b28_m51),
    .Q(pp_row79_7));
 sky130_fd_sc_hd__dfxtp_1 _0481_ (.CLK(clknet_leaf_205_clk),
    .D(booth_b30_m49),
    .Q(pp_row79_8));
 sky130_fd_sc_hd__dfxtp_1 _0482_ (.CLK(clknet_leaf_157_clk),
    .D(booth_b32_m47),
    .Q(pp_row79_9));
 sky130_fd_sc_hd__dfxtp_1 _0483_ (.CLK(clknet_leaf_156_clk),
    .D(booth_b34_m45),
    .Q(pp_row79_10));
 sky130_fd_sc_hd__dfxtp_1 _0484_ (.CLK(clknet_leaf_156_clk),
    .D(booth_b36_m43),
    .Q(pp_row79_11));
 sky130_fd_sc_hd__dfxtp_1 _0485_ (.CLK(clknet_leaf_205_clk),
    .D(booth_b38_m41),
    .Q(pp_row79_12));
 sky130_fd_sc_hd__dfxtp_1 _0486_ (.CLK(clknet_leaf_205_clk),
    .D(booth_b40_m39),
    .Q(pp_row79_13));
 sky130_fd_sc_hd__dfxtp_1 _0487_ (.CLK(clknet_leaf_205_clk),
    .D(booth_b42_m37),
    .Q(pp_row79_14));
 sky130_fd_sc_hd__dfxtp_1 _0488_ (.CLK(clknet_leaf_129_clk),
    .D(booth_b60_m55),
    .Q(pp_row115_5));
 sky130_fd_sc_hd__dfxtp_1 _0489_ (.CLK(clknet_leaf_159_clk),
    .D(booth_b44_m35),
    .Q(pp_row79_15));
 sky130_fd_sc_hd__dfxtp_1 _0490_ (.CLK(clknet_leaf_159_clk),
    .D(booth_b46_m33),
    .Q(pp_row79_16));
 sky130_fd_sc_hd__dfxtp_1 _0491_ (.CLK(clknet_leaf_159_clk),
    .D(booth_b48_m31),
    .Q(pp_row79_17));
 sky130_fd_sc_hd__dfxtp_1 _0492_ (.CLK(clknet_leaf_159_clk),
    .D(booth_b50_m29),
    .Q(pp_row79_18));
 sky130_fd_sc_hd__dfxtp_1 _0493_ (.CLK(clknet_leaf_161_clk),
    .D(booth_b52_m27),
    .Q(pp_row79_19));
 sky130_fd_sc_hd__dfxtp_1 _0494_ (.CLK(clknet_leaf_159_clk),
    .D(booth_b54_m25),
    .Q(pp_row79_20));
 sky130_fd_sc_hd__dfxtp_1 _0495_ (.CLK(clknet_leaf_158_clk),
    .D(booth_b56_m23),
    .Q(pp_row79_21));
 sky130_fd_sc_hd__dfxtp_1 _0496_ (.CLK(clknet_leaf_158_clk),
    .D(booth_b58_m21),
    .Q(pp_row79_22));
 sky130_fd_sc_hd__dfxtp_1 _0497_ (.CLK(clknet_leaf_158_clk),
    .D(booth_b60_m19),
    .Q(pp_row79_23));
 sky130_fd_sc_hd__dfxtp_1 _0498_ (.CLK(clknet_leaf_208_clk),
    .D(booth_b62_m17),
    .Q(pp_row79_24));
 sky130_fd_sc_hd__dfxtp_1 _0499_ (.CLK(clknet_leaf_126_clk),
    .D(booth_b62_m53),
    .Q(pp_row115_6));
 sky130_fd_sc_hd__dfxtp_1 _0500_ (.CLK(clknet_leaf_179_clk),
    .D(booth_b62_m64),
    .Q(pp_row126_1));
 sky130_fd_sc_hd__dfxtp_1 _0501_ (.CLK(clknet_leaf_208_clk),
    .D(booth_b64_m15),
    .Q(pp_row79_25));
 sky130_fd_sc_hd__dfxtp_1 _0502_ (.CLK(clknet_leaf_195_clk),
    .D(net233),
    .Q(pp_row79_26));
 sky130_fd_sc_hd__dfxtp_1 _0503_ (.CLK(clknet_leaf_206_clk),
    .D(booth_b16_m64),
    .Q(pp_row80_1));
 sky130_fd_sc_hd__dfxtp_1 _0504_ (.CLK(clknet_leaf_157_clk),
    .D(booth_b18_m62),
    .Q(pp_row80_2));
 sky130_fd_sc_hd__dfxtp_1 _0505_ (.CLK(clknet_leaf_172_clk),
    .D(booth_b20_m60),
    .Q(pp_row80_3));
 sky130_fd_sc_hd__dfxtp_1 _0506_ (.CLK(clknet_leaf_172_clk),
    .D(booth_b22_m58),
    .Q(pp_row80_4));
 sky130_fd_sc_hd__dfxtp_1 _0507_ (.CLK(clknet_leaf_172_clk),
    .D(booth_b24_m56),
    .Q(pp_row80_5));
 sky130_fd_sc_hd__dfxtp_1 _0508_ (.CLK(clknet_leaf_173_clk),
    .D(booth_b26_m54),
    .Q(pp_row80_6));
 sky130_fd_sc_hd__dfxtp_1 _0509_ (.CLK(clknet_leaf_173_clk),
    .D(booth_b28_m52),
    .Q(pp_row80_7));
 sky130_fd_sc_hd__dfxtp_1 _0510_ (.CLK(clknet_leaf_173_clk),
    .D(booth_b30_m50),
    .Q(pp_row80_8));
 sky130_fd_sc_hd__dfxtp_1 _0511_ (.CLK(clknet_leaf_126_clk),
    .D(booth_b64_m51),
    .Q(pp_row115_7));
 sky130_fd_sc_hd__dfxtp_1 _0512_ (.CLK(clknet_leaf_190_clk),
    .D(booth_b32_m48),
    .Q(pp_row80_9));
 sky130_fd_sc_hd__dfxtp_1 _0513_ (.CLK(clknet_leaf_191_clk),
    .D(booth_b34_m46),
    .Q(pp_row80_10));
 sky130_fd_sc_hd__dfxtp_1 _0514_ (.CLK(clknet_leaf_191_clk),
    .D(booth_b36_m44),
    .Q(pp_row80_11));
 sky130_fd_sc_hd__dfxtp_1 _0515_ (.CLK(clknet_leaf_156_clk),
    .D(booth_b38_m42),
    .Q(pp_row80_12));
 sky130_fd_sc_hd__dfxtp_1 _0516_ (.CLK(clknet_leaf_160_clk),
    .D(booth_b40_m40),
    .Q(pp_row80_13));
 sky130_fd_sc_hd__dfxtp_1 _0517_ (.CLK(clknet_leaf_155_clk),
    .D(booth_b42_m38),
    .Q(pp_row80_14));
 sky130_fd_sc_hd__dfxtp_1 _0518_ (.CLK(clknet_leaf_166_clk),
    .D(booth_b44_m36),
    .Q(pp_row80_15));
 sky130_fd_sc_hd__dfxtp_1 _0519_ (.CLK(clknet_leaf_166_clk),
    .D(booth_b46_m34),
    .Q(pp_row80_16));
 sky130_fd_sc_hd__dfxtp_1 _0520_ (.CLK(clknet_leaf_166_clk),
    .D(booth_b48_m32),
    .Q(pp_row80_17));
 sky130_fd_sc_hd__dfxtp_1 _0521_ (.CLK(clknet_leaf_159_clk),
    .D(booth_b50_m30),
    .Q(pp_row80_18));
 sky130_fd_sc_hd__dfxtp_2 _0522_ (.CLK(clknet_leaf_181_clk),
    .D(net146),
    .Q(pp_row115_8));
 sky130_fd_sc_hd__dfxtp_1 _0523_ (.CLK(clknet_leaf_163_clk),
    .D(booth_b52_m28),
    .Q(pp_row80_19));
 sky130_fd_sc_hd__dfxtp_1 _0524_ (.CLK(clknet_leaf_167_clk),
    .D(booth_b54_m26),
    .Q(pp_row80_20));
 sky130_fd_sc_hd__dfxtp_1 _0525_ (.CLK(clknet_leaf_162_clk),
    .D(booth_b56_m24),
    .Q(pp_row80_21));
 sky130_fd_sc_hd__dfxtp_1 _0526_ (.CLK(clknet_leaf_162_clk),
    .D(booth_b58_m22),
    .Q(pp_row80_22));
 sky130_fd_sc_hd__dfxtp_1 _0527_ (.CLK(clknet_leaf_162_clk),
    .D(booth_b60_m20),
    .Q(pp_row80_23));
 sky130_fd_sc_hd__dfxtp_1 _0528_ (.CLK(clknet_leaf_159_clk),
    .D(booth_b62_m18),
    .Q(pp_row80_24));
 sky130_fd_sc_hd__dfxtp_1 _0529_ (.CLK(clknet_leaf_159_clk),
    .D(booth_b64_m16),
    .Q(pp_row80_25));
 sky130_fd_sc_hd__dfxtp_1 _0530_ (.CLK(clknet_leaf_194_clk),
    .D(net235),
    .Q(pp_row80_26));
 sky130_fd_sc_hd__dfxtp_1 _0531_ (.CLK(clknet_leaf_162_clk),
    .D(\notsign$5034 ),
    .Q(pp_row81_0));
 sky130_fd_sc_hd__dfxtp_1 _0532_ (.CLK(clknet_leaf_159_clk),
    .D(booth_b18_m63),
    .Q(pp_row81_1));
 sky130_fd_sc_hd__dfxtp_1 _0533_ (.CLK(clknet_leaf_131_clk),
    .D(booth_b52_m64),
    .Q(pp_row116_1));
 sky130_fd_sc_hd__dfxtp_1 _0534_ (.CLK(clknet_leaf_159_clk),
    .D(booth_b20_m61),
    .Q(pp_row81_2));
 sky130_fd_sc_hd__dfxtp_1 _0535_ (.CLK(clknet_leaf_166_clk),
    .D(booth_b22_m59),
    .Q(pp_row81_3));
 sky130_fd_sc_hd__dfxtp_1 _0536_ (.CLK(clknet_leaf_163_clk),
    .D(booth_b24_m57),
    .Q(pp_row81_4));
 sky130_fd_sc_hd__dfxtp_1 _0537_ (.CLK(clknet_leaf_163_clk),
    .D(booth_b26_m55),
    .Q(pp_row81_5));
 sky130_fd_sc_hd__dfxtp_1 _0538_ (.CLK(clknet_leaf_166_clk),
    .D(booth_b28_m53),
    .Q(pp_row81_6));
 sky130_fd_sc_hd__dfxtp_1 _0539_ (.CLK(clknet_leaf_163_clk),
    .D(booth_b30_m51),
    .Q(pp_row81_7));
 sky130_fd_sc_hd__dfxtp_1 _0540_ (.CLK(clknet_leaf_165_clk),
    .D(booth_b32_m49),
    .Q(pp_row81_8));
 sky130_fd_sc_hd__dfxtp_1 _0541_ (.CLK(clknet_leaf_169_clk),
    .D(booth_b34_m47),
    .Q(pp_row81_9));
 sky130_fd_sc_hd__dfxtp_1 _0542_ (.CLK(clknet_leaf_170_clk),
    .D(booth_b36_m45),
    .Q(pp_row81_10));
 sky130_fd_sc_hd__dfxtp_1 _0543_ (.CLK(clknet_leaf_170_clk),
    .D(booth_b38_m43),
    .Q(pp_row81_11));
 sky130_fd_sc_hd__dfxtp_1 _0544_ (.CLK(clknet_leaf_126_clk),
    .D(booth_b54_m62),
    .Q(pp_row116_2));
 sky130_fd_sc_hd__dfxtp_1 _0545_ (.CLK(clknet_leaf_167_clk),
    .D(booth_b40_m41),
    .Q(pp_row81_12));
 sky130_fd_sc_hd__dfxtp_1 _0546_ (.CLK(clknet_leaf_171_clk),
    .D(booth_b42_m39),
    .Q(pp_row81_13));
 sky130_fd_sc_hd__dfxtp_1 _0547_ (.CLK(clknet_leaf_171_clk),
    .D(booth_b44_m37),
    .Q(pp_row81_14));
 sky130_fd_sc_hd__dfxtp_1 _0548_ (.CLK(clknet_leaf_171_clk),
    .D(booth_b46_m35),
    .Q(pp_row81_15));
 sky130_fd_sc_hd__dfxtp_1 _0549_ (.CLK(clknet_leaf_171_clk),
    .D(booth_b48_m33),
    .Q(pp_row81_16));
 sky130_fd_sc_hd__dfxtp_1 _0550_ (.CLK(clknet_leaf_172_clk),
    .D(booth_b50_m31),
    .Q(pp_row81_17));
 sky130_fd_sc_hd__dfxtp_1 _0551_ (.CLK(clknet_leaf_171_clk),
    .D(booth_b52_m29),
    .Q(pp_row81_18));
 sky130_fd_sc_hd__dfxtp_1 _0552_ (.CLK(clknet_leaf_171_clk),
    .D(booth_b54_m27),
    .Q(pp_row81_19));
 sky130_fd_sc_hd__dfxtp_1 _0553_ (.CLK(clknet_leaf_171_clk),
    .D(booth_b56_m25),
    .Q(pp_row81_20));
 sky130_fd_sc_hd__dfxtp_1 _0554_ (.CLK(clknet_leaf_189_clk),
    .D(booth_b58_m23),
    .Q(pp_row81_21));
 sky130_fd_sc_hd__dfxtp_1 _0555_ (.CLK(clknet_leaf_126_clk),
    .D(booth_b56_m60),
    .Q(pp_row116_3));
 sky130_fd_sc_hd__dfxtp_1 _0556_ (.CLK(clknet_leaf_189_clk),
    .D(booth_b60_m21),
    .Q(pp_row81_22));
 sky130_fd_sc_hd__dfxtp_1 _0557_ (.CLK(clknet_leaf_189_clk),
    .D(booth_b62_m19),
    .Q(pp_row81_23));
 sky130_fd_sc_hd__dfxtp_1 _0558_ (.CLK(clknet_leaf_157_clk),
    .D(booth_b64_m17),
    .Q(pp_row81_24));
 sky130_fd_sc_hd__dfxtp_2 _0559_ (.CLK(clknet_leaf_195_clk),
    .D(net236),
    .Q(pp_row81_25));
 sky130_fd_sc_hd__dfxtp_1 _0560_ (.CLK(clknet_leaf_186_clk),
    .D(booth_b18_m64),
    .Q(pp_row82_1));
 sky130_fd_sc_hd__dfxtp_1 _0561_ (.CLK(clknet_leaf_186_clk),
    .D(booth_b20_m62),
    .Q(pp_row82_2));
 sky130_fd_sc_hd__dfxtp_1 _0562_ (.CLK(clknet_leaf_186_clk),
    .D(booth_b22_m60),
    .Q(pp_row82_3));
 sky130_fd_sc_hd__dfxtp_1 _0563_ (.CLK(clknet_leaf_186_clk),
    .D(booth_b24_m58),
    .Q(pp_row82_4));
 sky130_fd_sc_hd__dfxtp_1 _0564_ (.CLK(clknet_leaf_186_clk),
    .D(booth_b26_m56),
    .Q(pp_row82_5));
 sky130_fd_sc_hd__dfxtp_1 _0565_ (.CLK(clknet_leaf_188_clk),
    .D(booth_b28_m54),
    .Q(pp_row82_6));
 sky130_fd_sc_hd__dfxtp_1 _0566_ (.CLK(clknet_leaf_126_clk),
    .D(booth_b58_m58),
    .Q(pp_row116_4));
 sky130_fd_sc_hd__dfxtp_1 _0567_ (.CLK(clknet_leaf_188_clk),
    .D(booth_b30_m52),
    .Q(pp_row82_7));
 sky130_fd_sc_hd__dfxtp_1 _0568_ (.CLK(clknet_leaf_188_clk),
    .D(booth_b32_m50),
    .Q(pp_row82_8));
 sky130_fd_sc_hd__dfxtp_1 _0569_ (.CLK(clknet_leaf_188_clk),
    .D(booth_b34_m48),
    .Q(pp_row82_9));
 sky130_fd_sc_hd__dfxtp_1 _0570_ (.CLK(clknet_leaf_188_clk),
    .D(booth_b36_m46),
    .Q(pp_row82_10));
 sky130_fd_sc_hd__dfxtp_1 _0571_ (.CLK(clknet_leaf_188_clk),
    .D(booth_b38_m44),
    .Q(pp_row82_11));
 sky130_fd_sc_hd__dfxtp_1 _0572_ (.CLK(clknet_leaf_189_clk),
    .D(booth_b40_m42),
    .Q(pp_row82_12));
 sky130_fd_sc_hd__dfxtp_1 _0573_ (.CLK(clknet_leaf_190_clk),
    .D(booth_b42_m40),
    .Q(pp_row82_13));
 sky130_fd_sc_hd__dfxtp_1 _0574_ (.CLK(clknet_leaf_190_clk),
    .D(booth_b44_m38),
    .Q(pp_row82_14));
 sky130_fd_sc_hd__dfxtp_1 _0575_ (.CLK(clknet_leaf_189_clk),
    .D(booth_b46_m36),
    .Q(pp_row82_15));
 sky130_fd_sc_hd__dfxtp_1 _0576_ (.CLK(clknet_leaf_189_clk),
    .D(booth_b48_m34),
    .Q(pp_row82_16));
 sky130_fd_sc_hd__dfxtp_1 _0577_ (.CLK(clknet_leaf_120_clk),
    .D(booth_b60_m56),
    .Q(pp_row116_5));
 sky130_fd_sc_hd__dfxtp_1 _0578_ (.CLK(clknet_leaf_189_clk),
    .D(booth_b50_m32),
    .Q(pp_row82_17));
 sky130_fd_sc_hd__dfxtp_1 _0579_ (.CLK(clknet_leaf_205_clk),
    .D(booth_b52_m30),
    .Q(pp_row82_18));
 sky130_fd_sc_hd__dfxtp_1 _0580_ (.CLK(clknet_leaf_189_clk),
    .D(booth_b54_m28),
    .Q(pp_row82_19));
 sky130_fd_sc_hd__dfxtp_1 _0581_ (.CLK(clknet_leaf_205_clk),
    .D(booth_b56_m26),
    .Q(pp_row82_20));
 sky130_fd_sc_hd__dfxtp_1 _0582_ (.CLK(clknet_leaf_173_clk),
    .D(booth_b58_m24),
    .Q(pp_row82_21));
 sky130_fd_sc_hd__dfxtp_1 _0583_ (.CLK(clknet_leaf_173_clk),
    .D(booth_b60_m22),
    .Q(pp_row82_22));
 sky130_fd_sc_hd__dfxtp_1 _0584_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b62_m20),
    .Q(pp_row82_23));
 sky130_fd_sc_hd__dfxtp_1 _0585_ (.CLK(clknet_leaf_188_clk),
    .D(booth_b64_m18),
    .Q(pp_row82_24));
 sky130_fd_sc_hd__dfxtp_1 _0586_ (.CLK(clknet_leaf_194_clk),
    .D(net237),
    .Q(pp_row82_25));
 sky130_fd_sc_hd__dfxtp_1 _0587_ (.CLK(clknet_leaf_186_clk),
    .D(\notsign$5104 ),
    .Q(pp_row83_0));
 sky130_fd_sc_hd__dfxtp_1 _0588_ (.CLK(clknet_leaf_120_clk),
    .D(booth_b62_m54),
    .Q(pp_row116_6));
 sky130_fd_sc_hd__dfxtp_1 _0589_ (.CLK(clknet_leaf_186_clk),
    .D(booth_b20_m63),
    .Q(pp_row83_1));
 sky130_fd_sc_hd__dfxtp_1 _0590_ (.CLK(clknet_leaf_186_clk),
    .D(booth_b22_m61),
    .Q(pp_row83_2));
 sky130_fd_sc_hd__dfxtp_1 _0591_ (.CLK(clknet_leaf_186_clk),
    .D(booth_b24_m59),
    .Q(pp_row83_3));
 sky130_fd_sc_hd__dfxtp_1 _0592_ (.CLK(clknet_leaf_186_clk),
    .D(booth_b26_m57),
    .Q(pp_row83_4));
 sky130_fd_sc_hd__dfxtp_1 _0593_ (.CLK(clknet_leaf_186_clk),
    .D(booth_b28_m55),
    .Q(pp_row83_5));
 sky130_fd_sc_hd__dfxtp_1 _0594_ (.CLK(clknet_leaf_193_clk),
    .D(booth_b30_m53),
    .Q(pp_row83_6));
 sky130_fd_sc_hd__dfxtp_1 _0595_ (.CLK(clknet_leaf_193_clk),
    .D(booth_b32_m51),
    .Q(pp_row83_7));
 sky130_fd_sc_hd__dfxtp_1 _0596_ (.CLK(clknet_leaf_193_clk),
    .D(booth_b34_m49),
    .Q(pp_row83_8));
 sky130_fd_sc_hd__dfxtp_1 _0597_ (.CLK(clknet_leaf_188_clk),
    .D(booth_b36_m47),
    .Q(pp_row83_9));
 sky130_fd_sc_hd__dfxtp_1 _0598_ (.CLK(clknet_leaf_188_clk),
    .D(booth_b38_m45),
    .Q(pp_row83_10));
 sky130_fd_sc_hd__dfxtp_1 _0599_ (.CLK(clknet_leaf_126_clk),
    .D(booth_b64_m52),
    .Q(pp_row116_7));
 sky130_fd_sc_hd__dfxtp_1 _0600_ (.CLK(clknet_leaf_188_clk),
    .D(booth_b40_m43),
    .Q(pp_row83_11));
 sky130_fd_sc_hd__dfxtp_1 _0601_ (.CLK(clknet_leaf_188_clk),
    .D(booth_b42_m41),
    .Q(pp_row83_12));
 sky130_fd_sc_hd__dfxtp_1 _0602_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b44_m39),
    .Q(pp_row83_13));
 sky130_fd_sc_hd__dfxtp_1 _0603_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b46_m37),
    .Q(pp_row83_14));
 sky130_fd_sc_hd__dfxtp_1 _0604_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b48_m35),
    .Q(pp_row83_15));
 sky130_fd_sc_hd__dfxtp_1 _0605_ (.CLK(clknet_leaf_188_clk),
    .D(booth_b50_m33),
    .Q(pp_row83_16));
 sky130_fd_sc_hd__dfxtp_1 _0606_ (.CLK(clknet_leaf_173_clk),
    .D(booth_b52_m31),
    .Q(pp_row83_17));
 sky130_fd_sc_hd__dfxtp_1 _0607_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b54_m29),
    .Q(pp_row83_18));
 sky130_fd_sc_hd__dfxtp_1 _0608_ (.CLK(clknet_leaf_172_clk),
    .D(booth_b56_m27),
    .Q(pp_row83_19));
 sky130_fd_sc_hd__dfxtp_1 _0609_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b58_m25),
    .Q(pp_row83_20));
 sky130_fd_sc_hd__dfxtp_2 _0610_ (.CLK(clknet_leaf_181_clk),
    .D(net147),
    .Q(pp_row116_8));
 sky130_fd_sc_hd__dfxtp_1 _0611_ (.CLK(clknet_leaf_179_clk),
    .D(booth_b64_m62),
    .Q(pp_row126_2));
 sky130_fd_sc_hd__dfxtp_1 _0612_ (.CLK(clknet_leaf_173_clk),
    .D(booth_b60_m23),
    .Q(pp_row83_21));
 sky130_fd_sc_hd__dfxtp_1 _0613_ (.CLK(clknet_leaf_173_clk),
    .D(booth_b62_m21),
    .Q(pp_row83_22));
 sky130_fd_sc_hd__dfxtp_1 _0614_ (.CLK(clknet_leaf_189_clk),
    .D(booth_b64_m19),
    .Q(pp_row83_23));
 sky130_fd_sc_hd__dfxtp_1 _0615_ (.CLK(clknet_leaf_195_clk),
    .D(net238),
    .Q(pp_row83_24));
 sky130_fd_sc_hd__dfxtp_1 _0616_ (.CLK(clknet_leaf_187_clk),
    .D(booth_b20_m64),
    .Q(pp_row84_1));
 sky130_fd_sc_hd__dfxtp_1 _0617_ (.CLK(clknet_leaf_187_clk),
    .D(booth_b22_m62),
    .Q(pp_row84_2));
 sky130_fd_sc_hd__dfxtp_1 _0618_ (.CLK(clknet_leaf_187_clk),
    .D(booth_b24_m60),
    .Q(pp_row84_3));
 sky130_fd_sc_hd__dfxtp_1 _0619_ (.CLK(clknet_leaf_187_clk),
    .D(booth_b26_m58),
    .Q(pp_row84_4));
 sky130_fd_sc_hd__dfxtp_1 _0620_ (.CLK(clknet_leaf_187_clk),
    .D(booth_b28_m56),
    .Q(pp_row84_5));
 sky130_fd_sc_hd__dfxtp_1 _0621_ (.CLK(clknet_leaf_187_clk),
    .D(booth_b30_m54),
    .Q(pp_row84_6));
 sky130_fd_sc_hd__dfxtp_1 _0622_ (.CLK(clknet_leaf_164_clk),
    .D(\notsign$6294 ),
    .Q(pp_row117_0));
 sky130_fd_sc_hd__dfxtp_1 _0623_ (.CLK(clknet_leaf_187_clk),
    .D(booth_b32_m52),
    .Q(pp_row84_7));
 sky130_fd_sc_hd__dfxtp_1 _0624_ (.CLK(clknet_leaf_187_clk),
    .D(booth_b34_m50),
    .Q(pp_row84_8));
 sky130_fd_sc_hd__dfxtp_1 _0625_ (.CLK(clknet_leaf_176_clk),
    .D(booth_b36_m48),
    .Q(pp_row84_9));
 sky130_fd_sc_hd__dfxtp_1 _0626_ (.CLK(clknet_leaf_176_clk),
    .D(booth_b38_m46),
    .Q(pp_row84_10));
 sky130_fd_sc_hd__dfxtp_1 _0627_ (.CLK(clknet_leaf_177_clk),
    .D(booth_b40_m44),
    .Q(pp_row84_11));
 sky130_fd_sc_hd__dfxtp_1 _0628_ (.CLK(clknet_leaf_179_clk),
    .D(booth_b42_m42),
    .Q(pp_row84_12));
 sky130_fd_sc_hd__dfxtp_1 _0629_ (.CLK(clknet_leaf_177_clk),
    .D(booth_b44_m40),
    .Q(pp_row84_13));
 sky130_fd_sc_hd__dfxtp_1 _0630_ (.CLK(clknet_leaf_178_clk),
    .D(booth_b46_m38),
    .Q(pp_row84_14));
 sky130_fd_sc_hd__dfxtp_1 _0631_ (.CLK(clknet_leaf_178_clk),
    .D(booth_b48_m36),
    .Q(pp_row84_15));
 sky130_fd_sc_hd__dfxtp_1 _0632_ (.CLK(clknet_leaf_178_clk),
    .D(booth_b50_m34),
    .Q(pp_row84_16));
 sky130_fd_sc_hd__dfxtp_1 _0633_ (.CLK(clknet_leaf_164_clk),
    .D(booth_b54_m63),
    .Q(pp_row117_1));
 sky130_fd_sc_hd__dfxtp_1 _0634_ (.CLK(clknet_leaf_178_clk),
    .D(booth_b52_m32),
    .Q(pp_row84_17));
 sky130_fd_sc_hd__dfxtp_1 _0635_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b54_m30),
    .Q(pp_row84_18));
 sky130_fd_sc_hd__dfxtp_1 _0636_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b56_m28),
    .Q(pp_row84_19));
 sky130_fd_sc_hd__dfxtp_1 _0637_ (.CLK(clknet_leaf_188_clk),
    .D(booth_b58_m26),
    .Q(pp_row84_20));
 sky130_fd_sc_hd__dfxtp_1 _0638_ (.CLK(clknet_leaf_188_clk),
    .D(booth_b60_m24),
    .Q(pp_row84_21));
 sky130_fd_sc_hd__dfxtp_1 _0639_ (.CLK(clknet_leaf_188_clk),
    .D(booth_b62_m22),
    .Q(pp_row84_22));
 sky130_fd_sc_hd__dfxtp_1 _0640_ (.CLK(clknet_leaf_186_clk),
    .D(booth_b64_m20),
    .Q(pp_row84_23));
 sky130_fd_sc_hd__dfxtp_1 _0641_ (.CLK(clknet_leaf_185_clk),
    .D(net239),
    .Q(pp_row84_24));
 sky130_fd_sc_hd__dfxtp_1 _0642_ (.CLK(clknet_leaf_183_clk),
    .D(\notsign$5174 ),
    .Q(pp_row85_0));
 sky130_fd_sc_hd__dfxtp_1 _0643_ (.CLK(clknet_leaf_180_clk),
    .D(booth_b22_m63),
    .Q(pp_row85_1));
 sky130_fd_sc_hd__dfxtp_1 _0644_ (.CLK(clknet_leaf_164_clk),
    .D(booth_b56_m61),
    .Q(pp_row117_2));
 sky130_fd_sc_hd__dfxtp_1 _0645_ (.CLK(clknet_leaf_183_clk),
    .D(booth_b24_m61),
    .Q(pp_row85_2));
 sky130_fd_sc_hd__dfxtp_1 _0646_ (.CLK(clknet_leaf_182_clk),
    .D(booth_b26_m59),
    .Q(pp_row85_3));
 sky130_fd_sc_hd__dfxtp_1 _0647_ (.CLK(clknet_leaf_183_clk),
    .D(booth_b28_m57),
    .Q(pp_row85_4));
 sky130_fd_sc_hd__dfxtp_1 _0648_ (.CLK(clknet_leaf_183_clk),
    .D(booth_b30_m55),
    .Q(pp_row85_5));
 sky130_fd_sc_hd__dfxtp_1 _0649_ (.CLK(clknet_leaf_165_clk),
    .D(booth_b32_m53),
    .Q(pp_row85_6));
 sky130_fd_sc_hd__dfxtp_1 _0650_ (.CLK(clknet_leaf_165_clk),
    .D(booth_b34_m51),
    .Q(pp_row85_7));
 sky130_fd_sc_hd__dfxtp_1 _0651_ (.CLK(clknet_leaf_168_clk),
    .D(booth_b36_m49),
    .Q(pp_row85_8));
 sky130_fd_sc_hd__dfxtp_1 _0652_ (.CLK(clknet_leaf_169_clk),
    .D(booth_b38_m47),
    .Q(pp_row85_9));
 sky130_fd_sc_hd__dfxtp_1 _0653_ (.CLK(clknet_leaf_169_clk),
    .D(booth_b40_m45),
    .Q(pp_row85_10));
 sky130_fd_sc_hd__dfxtp_1 _0654_ (.CLK(clknet_leaf_169_clk),
    .D(booth_b42_m43),
    .Q(pp_row85_11));
 sky130_fd_sc_hd__dfxtp_1 _0655_ (.CLK(clknet_leaf_131_clk),
    .D(booth_b58_m59),
    .Q(pp_row117_3));
 sky130_fd_sc_hd__dfxtp_1 _0656_ (.CLK(clknet_leaf_178_clk),
    .D(booth_b44_m41),
    .Q(pp_row85_12));
 sky130_fd_sc_hd__dfxtp_1 _0657_ (.CLK(clknet_leaf_178_clk),
    .D(booth_b46_m39),
    .Q(pp_row85_13));
 sky130_fd_sc_hd__dfxtp_1 _0658_ (.CLK(clknet_leaf_177_clk),
    .D(booth_b48_m37),
    .Q(pp_row85_14));
 sky130_fd_sc_hd__dfxtp_1 _0659_ (.CLK(clknet_leaf_175_clk),
    .D(booth_b50_m35),
    .Q(pp_row85_15));
 sky130_fd_sc_hd__dfxtp_1 _0660_ (.CLK(clknet_leaf_175_clk),
    .D(booth_b52_m33),
    .Q(pp_row85_16));
 sky130_fd_sc_hd__dfxtp_1 _0661_ (.CLK(clknet_leaf_176_clk),
    .D(booth_b54_m31),
    .Q(pp_row85_17));
 sky130_fd_sc_hd__dfxtp_1 _0662_ (.CLK(clknet_leaf_172_clk),
    .D(booth_b56_m29),
    .Q(pp_row85_18));
 sky130_fd_sc_hd__dfxtp_1 _0663_ (.CLK(clknet_leaf_172_clk),
    .D(booth_b58_m27),
    .Q(pp_row85_19));
 sky130_fd_sc_hd__dfxtp_1 _0664_ (.CLK(clknet_leaf_169_clk),
    .D(booth_b60_m25),
    .Q(pp_row85_20));
 sky130_fd_sc_hd__dfxtp_1 _0665_ (.CLK(clknet_leaf_187_clk),
    .D(booth_b62_m23),
    .Q(pp_row85_21));
 sky130_fd_sc_hd__dfxtp_1 _0666_ (.CLK(clknet_leaf_131_clk),
    .D(booth_b60_m57),
    .Q(pp_row117_4));
 sky130_fd_sc_hd__dfxtp_1 _0667_ (.CLK(clknet_leaf_187_clk),
    .D(booth_b64_m21),
    .Q(pp_row85_22));
 sky130_fd_sc_hd__dfxtp_1 _0668_ (.CLK(clknet_leaf_184_clk),
    .D(net240),
    .Q(pp_row85_23));
 sky130_fd_sc_hd__dfxtp_1 _0669_ (.CLK(clknet_leaf_180_clk),
    .D(booth_b22_m64),
    .Q(pp_row86_1));
 sky130_fd_sc_hd__dfxtp_1 _0670_ (.CLK(clknet_leaf_180_clk),
    .D(booth_b24_m62),
    .Q(pp_row86_2));
 sky130_fd_sc_hd__dfxtp_1 _0671_ (.CLK(clknet_leaf_175_clk),
    .D(booth_b26_m60),
    .Q(pp_row86_3));
 sky130_fd_sc_hd__dfxtp_1 _0672_ (.CLK(clknet_leaf_175_clk),
    .D(booth_b28_m58),
    .Q(pp_row86_4));
 sky130_fd_sc_hd__dfxtp_1 _0673_ (.CLK(clknet_leaf_175_clk),
    .D(booth_b30_m56),
    .Q(pp_row86_5));
 sky130_fd_sc_hd__dfxtp_1 _0674_ (.CLK(clknet_leaf_170_clk),
    .D(booth_b32_m54),
    .Q(pp_row86_6));
 sky130_fd_sc_hd__dfxtp_1 _0675_ (.CLK(clknet_leaf_170_clk),
    .D(booth_b34_m52),
    .Q(pp_row86_7));
 sky130_fd_sc_hd__dfxtp_1 _0676_ (.CLK(clknet_leaf_176_clk),
    .D(booth_b36_m50),
    .Q(pp_row86_8));
 sky130_fd_sc_hd__dfxtp_1 _0677_ (.CLK(clknet_leaf_131_clk),
    .D(booth_b62_m55),
    .Q(pp_row117_5));
 sky130_fd_sc_hd__dfxtp_1 _0678_ (.CLK(clknet_leaf_179_clk),
    .D(booth_b38_m48),
    .Q(pp_row86_9));
 sky130_fd_sc_hd__dfxtp_1 _0679_ (.CLK(clknet_leaf_179_clk),
    .D(booth_b40_m46),
    .Q(pp_row86_10));
 sky130_fd_sc_hd__dfxtp_1 _0680_ (.CLK(clknet_leaf_180_clk),
    .D(booth_b42_m44),
    .Q(pp_row86_11));
 sky130_fd_sc_hd__dfxtp_1 _0681_ (.CLK(clknet_leaf_169_clk),
    .D(booth_b44_m42),
    .Q(pp_row86_12));
 sky130_fd_sc_hd__dfxtp_1 _0682_ (.CLK(clknet_leaf_176_clk),
    .D(booth_b46_m40),
    .Q(pp_row86_13));
 sky130_fd_sc_hd__dfxtp_1 _0683_ (.CLK(clknet_leaf_176_clk),
    .D(booth_b48_m38),
    .Q(pp_row86_14));
 sky130_fd_sc_hd__dfxtp_1 _0684_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b50_m36),
    .Q(pp_row86_15));
 sky130_fd_sc_hd__dfxtp_1 _0685_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b52_m34),
    .Q(pp_row86_16));
 sky130_fd_sc_hd__dfxtp_1 _0686_ (.CLK(clknet_leaf_168_clk),
    .D(booth_b54_m32),
    .Q(pp_row86_17));
 sky130_fd_sc_hd__dfxtp_1 _0687_ (.CLK(clknet_leaf_168_clk),
    .D(booth_b56_m30),
    .Q(pp_row86_18));
 sky130_fd_sc_hd__dfxtp_1 _0688_ (.CLK(clknet_leaf_131_clk),
    .D(booth_b64_m53),
    .Q(pp_row117_6));
 sky130_fd_sc_hd__dfxtp_1 _0689_ (.CLK(clknet_leaf_168_clk),
    .D(booth_b58_m28),
    .Q(pp_row86_19));
 sky130_fd_sc_hd__dfxtp_1 _0690_ (.CLK(clknet_leaf_168_clk),
    .D(booth_b60_m26),
    .Q(pp_row86_20));
 sky130_fd_sc_hd__dfxtp_1 _0691_ (.CLK(clknet_leaf_168_clk),
    .D(booth_b62_m24),
    .Q(pp_row86_21));
 sky130_fd_sc_hd__dfxtp_1 _0692_ (.CLK(clknet_leaf_167_clk),
    .D(booth_b64_m22),
    .Q(pp_row86_22));
 sky130_fd_sc_hd__dfxtp_1 _0693_ (.CLK(clknet_leaf_184_clk),
    .D(net241),
    .Q(pp_row86_23));
 sky130_fd_sc_hd__dfxtp_1 _0694_ (.CLK(clknet_leaf_175_clk),
    .D(\notsign$5244 ),
    .Q(pp_row87_0));
 sky130_fd_sc_hd__dfxtp_1 _0695_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b24_m63),
    .Q(pp_row87_1));
 sky130_fd_sc_hd__dfxtp_1 _0696_ (.CLK(clknet_leaf_175_clk),
    .D(booth_b26_m61),
    .Q(pp_row87_2));
 sky130_fd_sc_hd__dfxtp_1 _0697_ (.CLK(clknet_leaf_187_clk),
    .D(booth_b28_m59),
    .Q(pp_row87_3));
 sky130_fd_sc_hd__dfxtp_1 _0698_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b30_m57),
    .Q(pp_row87_4));
 sky130_fd_sc_hd__dfxtp_2 _0699_ (.CLK(clknet_leaf_181_clk),
    .D(net148),
    .Q(pp_row117_7));
 sky130_fd_sc_hd__dfxtp_1 _0700_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b32_m55),
    .Q(pp_row87_5));
 sky130_fd_sc_hd__dfxtp_1 _0701_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b34_m53),
    .Q(pp_row87_6));
 sky130_fd_sc_hd__dfxtp_1 _0702_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b36_m51),
    .Q(pp_row87_7));
 sky130_fd_sc_hd__dfxtp_1 _0703_ (.CLK(clknet_leaf_174_clk),
    .D(booth_b38_m49),
    .Q(pp_row87_8));
 sky130_fd_sc_hd__dfxtp_1 _0704_ (.CLK(clknet_leaf_170_clk),
    .D(booth_b40_m47),
    .Q(pp_row87_9));
 sky130_fd_sc_hd__dfxtp_1 _0705_ (.CLK(clknet_leaf_172_clk),
    .D(booth_b42_m45),
    .Q(pp_row87_10));
 sky130_fd_sc_hd__dfxtp_1 _0706_ (.CLK(clknet_leaf_171_clk),
    .D(booth_b44_m43),
    .Q(pp_row87_11));
 sky130_fd_sc_hd__dfxtp_1 _0707_ (.CLK(clknet_leaf_167_clk),
    .D(booth_b46_m41),
    .Q(pp_row87_12));
 sky130_fd_sc_hd__dfxtp_1 _0708_ (.CLK(clknet_leaf_168_clk),
    .D(booth_b48_m39),
    .Q(pp_row87_13));
 sky130_fd_sc_hd__dfxtp_1 _0709_ (.CLK(clknet_leaf_168_clk),
    .D(booth_b50_m37),
    .Q(pp_row87_14));
 sky130_fd_sc_hd__dfxtp_1 _0710_ (.CLK(clknet_leaf_132_clk),
    .D(booth_b54_m64),
    .Q(pp_row118_1));
 sky130_fd_sc_hd__dfxtp_1 _0711_ (.CLK(clknet_leaf_165_clk),
    .D(booth_b52_m35),
    .Q(pp_row87_15));
 sky130_fd_sc_hd__dfxtp_1 _0712_ (.CLK(clknet_leaf_165_clk),
    .D(booth_b54_m33),
    .Q(pp_row87_16));
 sky130_fd_sc_hd__dfxtp_1 _0713_ (.CLK(clknet_leaf_165_clk),
    .D(booth_b56_m31),
    .Q(pp_row87_17));
 sky130_fd_sc_hd__dfxtp_1 _0714_ (.CLK(clknet_leaf_165_clk),
    .D(booth_b58_m29),
    .Q(pp_row87_18));
 sky130_fd_sc_hd__dfxtp_1 _0715_ (.CLK(clknet_leaf_165_clk),
    .D(booth_b60_m27),
    .Q(pp_row87_19));
 sky130_fd_sc_hd__dfxtp_1 _0716_ (.CLK(clknet_leaf_165_clk),
    .D(booth_b62_m25),
    .Q(pp_row87_20));
 sky130_fd_sc_hd__dfxtp_1 _0717_ (.CLK(clknet_leaf_179_clk),
    .D(booth_b64_m23),
    .Q(pp_row87_21));
 sky130_fd_sc_hd__dfxtp_1 _0718_ (.CLK(clknet_leaf_184_clk),
    .D(net242),
    .Q(pp_row87_22));
 sky130_fd_sc_hd__dfxtp_1 _0719_ (.CLK(clknet_leaf_134_clk),
    .D(booth_b24_m64),
    .Q(pp_row88_1));
 sky130_fd_sc_hd__dfxtp_1 _0720_ (.CLK(clknet_leaf_161_clk),
    .D(booth_b26_m62),
    .Q(pp_row88_2));
 sky130_fd_sc_hd__dfxtp_1 _0721_ (.CLK(clknet_leaf_132_clk),
    .D(booth_b56_m62),
    .Q(pp_row118_2));
 sky130_fd_sc_hd__dfxtp_1 _0722_ (.CLK(clknet_leaf_181_clk),
    .D(net158),
    .Q(pp_row126_3));
 sky130_fd_sc_hd__dfxtp_1 _0723_ (.CLK(clknet_leaf_135_clk),
    .D(booth_b28_m60),
    .Q(pp_row88_3));
 sky130_fd_sc_hd__dfxtp_1 _0724_ (.CLK(clknet_leaf_135_clk),
    .D(booth_b30_m58),
    .Q(pp_row88_4));
 sky130_fd_sc_hd__dfxtp_1 _0725_ (.CLK(clknet_leaf_135_clk),
    .D(booth_b32_m56),
    .Q(pp_row88_5));
 sky130_fd_sc_hd__dfxtp_1 _0726_ (.CLK(clknet_leaf_161_clk),
    .D(booth_b34_m54),
    .Q(pp_row88_6));
 sky130_fd_sc_hd__dfxtp_1 _0727_ (.CLK(clknet_leaf_161_clk),
    .D(booth_b36_m52),
    .Q(pp_row88_7));
 sky130_fd_sc_hd__dfxtp_1 _0728_ (.CLK(clknet_leaf_161_clk),
    .D(booth_b38_m50),
    .Q(pp_row88_8));
 sky130_fd_sc_hd__dfxtp_1 _0729_ (.CLK(clknet_leaf_135_clk),
    .D(booth_b40_m48),
    .Q(pp_row88_9));
 sky130_fd_sc_hd__dfxtp_1 _0730_ (.CLK(clknet_leaf_135_clk),
    .D(booth_b42_m46),
    .Q(pp_row88_10));
 sky130_fd_sc_hd__dfxtp_1 _0731_ (.CLK(clknet_leaf_135_clk),
    .D(booth_b44_m44),
    .Q(pp_row88_11));
 sky130_fd_sc_hd__dfxtp_1 _0732_ (.CLK(clknet_leaf_163_clk),
    .D(booth_b46_m42),
    .Q(pp_row88_12));
 sky130_fd_sc_hd__dfxtp_1 _0733_ (.CLK(clknet_leaf_132_clk),
    .D(booth_b58_m60),
    .Q(pp_row118_3));
 sky130_fd_sc_hd__dfxtp_1 _0734_ (.CLK(clknet_leaf_163_clk),
    .D(booth_b48_m40),
    .Q(pp_row88_13));
 sky130_fd_sc_hd__dfxtp_1 _0735_ (.CLK(clknet_leaf_162_clk),
    .D(booth_b50_m38),
    .Q(pp_row88_14));
 sky130_fd_sc_hd__dfxtp_1 _0736_ (.CLK(clknet_leaf_134_clk),
    .D(booth_b52_m36),
    .Q(pp_row88_15));
 sky130_fd_sc_hd__dfxtp_1 _0737_ (.CLK(clknet_leaf_134_clk),
    .D(booth_b54_m34),
    .Q(pp_row88_16));
 sky130_fd_sc_hd__dfxtp_1 _0738_ (.CLK(clknet_leaf_163_clk),
    .D(booth_b56_m32),
    .Q(pp_row88_17));
 sky130_fd_sc_hd__dfxtp_1 _0739_ (.CLK(clknet_leaf_163_clk),
    .D(booth_b58_m30),
    .Q(pp_row88_18));
 sky130_fd_sc_hd__dfxtp_1 _0740_ (.CLK(clknet_leaf_163_clk),
    .D(booth_b60_m28),
    .Q(pp_row88_19));
 sky130_fd_sc_hd__dfxtp_1 _0741_ (.CLK(clknet_leaf_171_clk),
    .D(booth_b62_m26),
    .Q(pp_row88_20));
 sky130_fd_sc_hd__dfxtp_1 _0742_ (.CLK(clknet_leaf_166_clk),
    .D(booth_b64_m24),
    .Q(pp_row88_21));
 sky130_fd_sc_hd__dfxtp_1 _0743_ (.CLK(clknet_leaf_184_clk),
    .D(net243),
    .Q(pp_row88_22));
 sky130_fd_sc_hd__dfxtp_1 _0744_ (.CLK(clknet_leaf_131_clk),
    .D(booth_b60_m58),
    .Q(pp_row118_4));
 sky130_fd_sc_hd__dfxtp_1 _0745_ (.CLK(clknet_leaf_143_clk),
    .D(\notsign$5314 ),
    .Q(pp_row89_0));
 sky130_fd_sc_hd__dfxtp_1 _0746_ (.CLK(clknet_leaf_142_clk),
    .D(booth_b26_m63),
    .Q(pp_row89_1));
 sky130_fd_sc_hd__dfxtp_1 _0747_ (.CLK(clknet_leaf_143_clk),
    .D(booth_b28_m61),
    .Q(pp_row89_2));
 sky130_fd_sc_hd__dfxtp_1 _0748_ (.CLK(clknet_leaf_160_clk),
    .D(booth_b30_m59),
    .Q(pp_row89_3));
 sky130_fd_sc_hd__dfxtp_1 _0749_ (.CLK(clknet_leaf_160_clk),
    .D(booth_b32_m57),
    .Q(pp_row89_4));
 sky130_fd_sc_hd__dfxtp_1 _0750_ (.CLK(clknet_leaf_160_clk),
    .D(booth_b34_m55),
    .Q(pp_row89_5));
 sky130_fd_sc_hd__dfxtp_1 _0751_ (.CLK(clknet_leaf_160_clk),
    .D(booth_b36_m53),
    .Q(pp_row89_6));
 sky130_fd_sc_hd__dfxtp_1 _0752_ (.CLK(clknet_leaf_160_clk),
    .D(booth_b38_m51),
    .Q(pp_row89_7));
 sky130_fd_sc_hd__dfxtp_1 _0753_ (.CLK(clknet_leaf_160_clk),
    .D(booth_b40_m49),
    .Q(pp_row89_8));
 sky130_fd_sc_hd__dfxtp_1 _0754_ (.CLK(clknet_leaf_160_clk),
    .D(booth_b42_m47),
    .Q(pp_row89_9));
 sky130_fd_sc_hd__dfxtp_1 _0755_ (.CLK(clknet_leaf_132_clk),
    .D(booth_b62_m56),
    .Q(pp_row118_5));
 sky130_fd_sc_hd__dfxtp_1 _0756_ (.CLK(clknet_leaf_161_clk),
    .D(booth_b44_m45),
    .Q(pp_row89_10));
 sky130_fd_sc_hd__dfxtp_1 _0757_ (.CLK(clknet_leaf_160_clk),
    .D(booth_b46_m43),
    .Q(pp_row89_11));
 sky130_fd_sc_hd__dfxtp_1 _0758_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b48_m41),
    .Q(pp_row89_12));
 sky130_fd_sc_hd__dfxtp_1 _0759_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b50_m39),
    .Q(pp_row89_13));
 sky130_fd_sc_hd__dfxtp_1 _0760_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b52_m37),
    .Q(pp_row89_14));
 sky130_fd_sc_hd__dfxtp_1 _0761_ (.CLK(clknet_leaf_161_clk),
    .D(booth_b54_m35),
    .Q(pp_row89_15));
 sky130_fd_sc_hd__dfxtp_1 _0762_ (.CLK(clknet_leaf_161_clk),
    .D(booth_b56_m33),
    .Q(pp_row89_16));
 sky130_fd_sc_hd__dfxtp_1 _0763_ (.CLK(clknet_leaf_161_clk),
    .D(booth_b58_m31),
    .Q(pp_row89_17));
 sky130_fd_sc_hd__dfxtp_1 _0764_ (.CLK(clknet_leaf_152_clk),
    .D(booth_b60_m29),
    .Q(pp_row89_18));
 sky130_fd_sc_hd__dfxtp_1 _0765_ (.CLK(clknet_leaf_152_clk),
    .D(booth_b62_m27),
    .Q(pp_row89_19));
 sky130_fd_sc_hd__dfxtp_1 _0766_ (.CLK(clknet_leaf_128_clk),
    .D(booth_b64_m54),
    .Q(pp_row118_6));
 sky130_fd_sc_hd__dfxtp_1 _0767_ (.CLK(clknet_leaf_152_clk),
    .D(booth_b64_m25),
    .Q(pp_row89_20));
 sky130_fd_sc_hd__dfxtp_2 _0768_ (.CLK(clknet_leaf_194_clk),
    .D(net244),
    .Q(pp_row89_21));
 sky130_fd_sc_hd__dfxtp_1 _0769_ (.CLK(clknet_leaf_138_clk),
    .D(booth_b26_m64),
    .Q(pp_row90_1));
 sky130_fd_sc_hd__dfxtp_1 _0770_ (.CLK(clknet_leaf_138_clk),
    .D(booth_b28_m62),
    .Q(pp_row90_2));
 sky130_fd_sc_hd__dfxtp_1 _0771_ (.CLK(clknet_leaf_144_clk),
    .D(booth_b30_m60),
    .Q(pp_row90_3));
 sky130_fd_sc_hd__dfxtp_1 _0772_ (.CLK(clknet_leaf_144_clk),
    .D(booth_b32_m58),
    .Q(pp_row90_4));
 sky130_fd_sc_hd__dfxtp_1 _0773_ (.CLK(clknet_leaf_144_clk),
    .D(booth_b34_m56),
    .Q(pp_row90_5));
 sky130_fd_sc_hd__dfxtp_1 _0774_ (.CLK(clknet_leaf_141_clk),
    .D(booth_b36_m54),
    .Q(pp_row90_6));
 sky130_fd_sc_hd__dfxtp_1 _0775_ (.CLK(clknet_leaf_141_clk),
    .D(booth_b38_m52),
    .Q(pp_row90_7));
 sky130_fd_sc_hd__dfxtp_1 _0776_ (.CLK(clknet_leaf_141_clk),
    .D(booth_b40_m50),
    .Q(pp_row90_8));
 sky130_fd_sc_hd__dfxtp_2 _0777_ (.CLK(clknet_leaf_181_clk),
    .D(net149),
    .Q(pp_row118_7));
 sky130_fd_sc_hd__dfxtp_1 _0778_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b42_m48),
    .Q(pp_row90_9));
 sky130_fd_sc_hd__dfxtp_1 _0779_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b44_m46),
    .Q(pp_row90_10));
 sky130_fd_sc_hd__dfxtp_1 _0780_ (.CLK(clknet_leaf_140_clk),
    .D(booth_b46_m44),
    .Q(pp_row90_11));
 sky130_fd_sc_hd__dfxtp_1 _0781_ (.CLK(clknet_leaf_140_clk),
    .D(booth_b48_m42),
    .Q(pp_row90_12));
 sky130_fd_sc_hd__dfxtp_1 _0782_ (.CLK(clknet_leaf_140_clk),
    .D(booth_b50_m40),
    .Q(pp_row90_13));
 sky130_fd_sc_hd__dfxtp_1 _0783_ (.CLK(clknet_leaf_140_clk),
    .D(booth_b52_m38),
    .Q(pp_row90_14));
 sky130_fd_sc_hd__dfxtp_1 _0784_ (.CLK(clknet_leaf_138_clk),
    .D(booth_b54_m36),
    .Q(pp_row90_15));
 sky130_fd_sc_hd__dfxtp_1 _0785_ (.CLK(clknet_leaf_138_clk),
    .D(booth_b56_m34),
    .Q(pp_row90_16));
 sky130_fd_sc_hd__dfxtp_1 _0786_ (.CLK(clknet_leaf_140_clk),
    .D(booth_b58_m32),
    .Q(pp_row90_17));
 sky130_fd_sc_hd__dfxtp_1 _0787_ (.CLK(clknet_leaf_139_clk),
    .D(booth_b60_m30),
    .Q(pp_row90_18));
 sky130_fd_sc_hd__dfxtp_1 _0788_ (.CLK(clknet_leaf_132_clk),
    .D(\notsign$6364 ),
    .Q(pp_row119_0));
 sky130_fd_sc_hd__dfxtp_1 _0789_ (.CLK(clknet_leaf_138_clk),
    .D(booth_b62_m28),
    .Q(pp_row90_19));
 sky130_fd_sc_hd__dfxtp_1 _0790_ (.CLK(clknet_leaf_139_clk),
    .D(booth_b64_m26),
    .Q(pp_row90_20));
 sky130_fd_sc_hd__dfxtp_2 _0791_ (.CLK(clknet_leaf_194_clk),
    .D(net246),
    .Q(pp_row90_21));
 sky130_fd_sc_hd__dfxtp_1 _0792_ (.CLK(clknet_leaf_93_clk),
    .D(\notsign$5384 ),
    .Q(pp_row91_0));
 sky130_fd_sc_hd__dfxtp_1 _0793_ (.CLK(clknet_leaf_93_clk),
    .D(booth_b28_m63),
    .Q(pp_row91_1));
 sky130_fd_sc_hd__dfxtp_1 _0794_ (.CLK(clknet_leaf_93_clk),
    .D(booth_b30_m61),
    .Q(pp_row91_2));
 sky130_fd_sc_hd__dfxtp_1 _0795_ (.CLK(clknet_leaf_139_clk),
    .D(booth_b32_m59),
    .Q(pp_row91_3));
 sky130_fd_sc_hd__dfxtp_1 _0796_ (.CLK(clknet_leaf_140_clk),
    .D(booth_b34_m57),
    .Q(pp_row91_4));
 sky130_fd_sc_hd__dfxtp_1 _0797_ (.CLK(clknet_leaf_139_clk),
    .D(booth_b36_m55),
    .Q(pp_row91_5));
 sky130_fd_sc_hd__dfxtp_1 _0798_ (.CLK(clknet_leaf_123_clk),
    .D(booth_b38_m53),
    .Q(pp_row91_6));
 sky130_fd_sc_hd__dfxtp_1 _0799_ (.CLK(clknet_leaf_132_clk),
    .D(booth_b56_m63),
    .Q(pp_row119_1));
 sky130_fd_sc_hd__dfxtp_1 _0800_ (.CLK(clknet_leaf_123_clk),
    .D(booth_b40_m51),
    .Q(pp_row91_7));
 sky130_fd_sc_hd__dfxtp_1 _0801_ (.CLK(clknet_leaf_139_clk),
    .D(booth_b42_m49),
    .Q(pp_row91_8));
 sky130_fd_sc_hd__dfxtp_1 _0802_ (.CLK(clknet_leaf_94_clk),
    .D(booth_b44_m47),
    .Q(pp_row91_9));
 sky130_fd_sc_hd__dfxtp_1 _0803_ (.CLK(clknet_leaf_94_clk),
    .D(booth_b46_m45),
    .Q(pp_row91_10));
 sky130_fd_sc_hd__dfxtp_1 _0804_ (.CLK(clknet_leaf_94_clk),
    .D(booth_b48_m43),
    .Q(pp_row91_11));
 sky130_fd_sc_hd__dfxtp_1 _0805_ (.CLK(clknet_leaf_94_clk),
    .D(booth_b50_m41),
    .Q(pp_row91_12));
 sky130_fd_sc_hd__dfxtp_1 _0806_ (.CLK(clknet_leaf_106_clk),
    .D(booth_b52_m39),
    .Q(pp_row91_13));
 sky130_fd_sc_hd__dfxtp_1 _0807_ (.CLK(clknet_leaf_94_clk),
    .D(booth_b54_m37),
    .Q(pp_row91_14));
 sky130_fd_sc_hd__dfxtp_1 _0808_ (.CLK(clknet_leaf_101_clk),
    .D(booth_b56_m35),
    .Q(pp_row91_15));
 sky130_fd_sc_hd__dfxtp_1 _0809_ (.CLK(clknet_leaf_97_clk),
    .D(booth_b58_m33),
    .Q(pp_row91_16));
 sky130_fd_sc_hd__dfxtp_1 _0810_ (.CLK(clknet_leaf_132_clk),
    .D(booth_b58_m61),
    .Q(pp_row119_2));
 sky130_fd_sc_hd__dfxtp_1 _0811_ (.CLK(clknet_leaf_97_clk),
    .D(booth_b60_m31),
    .Q(pp_row91_17));
 sky130_fd_sc_hd__dfxtp_1 _0812_ (.CLK(clknet_leaf_93_clk),
    .D(booth_b62_m29),
    .Q(pp_row91_18));
 sky130_fd_sc_hd__dfxtp_1 _0813_ (.CLK(clknet_leaf_94_clk),
    .D(booth_b64_m27),
    .Q(pp_row91_19));
 sky130_fd_sc_hd__dfxtp_2 _0814_ (.CLK(clknet_leaf_194_clk),
    .D(net247),
    .Q(pp_row91_20));
 sky130_fd_sc_hd__dfxtp_1 _0815_ (.CLK(clknet_leaf_139_clk),
    .D(booth_b28_m64),
    .Q(pp_row92_1));
 sky130_fd_sc_hd__dfxtp_1 _0816_ (.CLK(clknet_leaf_93_clk),
    .D(booth_b30_m62),
    .Q(pp_row92_2));
 sky130_fd_sc_hd__dfxtp_1 _0817_ (.CLK(clknet_leaf_111_clk),
    .D(booth_b32_m60),
    .Q(pp_row92_3));
 sky130_fd_sc_hd__dfxtp_1 _0818_ (.CLK(clknet_leaf_109_clk),
    .D(booth_b34_m58),
    .Q(pp_row92_4));
 sky130_fd_sc_hd__dfxtp_1 _0819_ (.CLK(clknet_leaf_111_clk),
    .D(booth_b36_m56),
    .Q(pp_row92_5));
 sky130_fd_sc_hd__dfxtp_1 _0820_ (.CLK(clknet_leaf_106_clk),
    .D(booth_b38_m54),
    .Q(pp_row92_6));
 sky130_fd_sc_hd__dfxtp_1 _0821_ (.CLK(clknet_leaf_164_clk),
    .D(booth_b60_m59),
    .Q(pp_row119_3));
 sky130_fd_sc_hd__dfxtp_1 _0822_ (.CLK(clknet_leaf_106_clk),
    .D(booth_b40_m52),
    .Q(pp_row92_7));
 sky130_fd_sc_hd__dfxtp_1 _0823_ (.CLK(clknet_leaf_108_clk),
    .D(booth_b42_m50),
    .Q(pp_row92_8));
 sky130_fd_sc_hd__dfxtp_1 _0824_ (.CLK(clknet_leaf_109_clk),
    .D(booth_b44_m48),
    .Q(pp_row92_9));
 sky130_fd_sc_hd__dfxtp_1 _0825_ (.CLK(clknet_leaf_109_clk),
    .D(booth_b46_m46),
    .Q(pp_row92_10));
 sky130_fd_sc_hd__dfxtp_1 _0826_ (.CLK(clknet_leaf_108_clk),
    .D(booth_b48_m44),
    .Q(pp_row92_11));
 sky130_fd_sc_hd__dfxtp_1 _0827_ (.CLK(clknet_leaf_108_clk),
    .D(booth_b50_m42),
    .Q(pp_row92_12));
 sky130_fd_sc_hd__dfxtp_1 _0828_ (.CLK(clknet_leaf_108_clk),
    .D(booth_b52_m40),
    .Q(pp_row92_13));
 sky130_fd_sc_hd__dfxtp_1 _0829_ (.CLK(clknet_leaf_108_clk),
    .D(booth_b54_m38),
    .Q(pp_row92_14));
 sky130_fd_sc_hd__dfxtp_1 _0830_ (.CLK(clknet_leaf_108_clk),
    .D(booth_b56_m36),
    .Q(pp_row92_15));
 sky130_fd_sc_hd__dfxtp_1 _0831_ (.CLK(clknet_leaf_107_clk),
    .D(booth_b58_m34),
    .Q(pp_row92_16));
 sky130_fd_sc_hd__dfxtp_1 _0832_ (.CLK(clknet_leaf_132_clk),
    .D(booth_b62_m57),
    .Q(pp_row119_4));
 sky130_fd_sc_hd__dfxtp_1 _0833_ (.CLK(clknet_leaf_180_clk),
    .D(\notsign$6644 ),
    .Q(pp_row127_0));
 sky130_fd_sc_hd__dfxtp_1 _0834_ (.CLK(clknet_leaf_106_clk),
    .D(booth_b60_m32),
    .Q(pp_row92_17));
 sky130_fd_sc_hd__dfxtp_1 _0835_ (.CLK(clknet_leaf_107_clk),
    .D(booth_b62_m30),
    .Q(pp_row92_18));
 sky130_fd_sc_hd__dfxtp_1 _0836_ (.CLK(clknet_leaf_106_clk),
    .D(booth_b64_m28),
    .Q(pp_row92_19));
 sky130_fd_sc_hd__dfxtp_2 _0837_ (.CLK(clknet_leaf_194_clk),
    .D(net248),
    .Q(pp_row92_20));
 sky130_fd_sc_hd__dfxtp_1 _0838_ (.CLK(clknet_leaf_105_clk),
    .D(\notsign$5454 ),
    .Q(pp_row93_0));
 sky130_fd_sc_hd__dfxtp_1 _0839_ (.CLK(clknet_leaf_105_clk),
    .D(booth_b30_m63),
    .Q(pp_row93_1));
 sky130_fd_sc_hd__dfxtp_1 _0840_ (.CLK(clknet_leaf_105_clk),
    .D(booth_b32_m61),
    .Q(pp_row93_2));
 sky130_fd_sc_hd__dfxtp_1 _0841_ (.CLK(clknet_leaf_102_clk),
    .D(booth_b34_m59),
    .Q(pp_row93_3));
 sky130_fd_sc_hd__dfxtp_1 _0842_ (.CLK(clknet_leaf_106_clk),
    .D(booth_b36_m57),
    .Q(pp_row93_4));
 sky130_fd_sc_hd__dfxtp_1 _0843_ (.CLK(clknet_leaf_106_clk),
    .D(booth_b38_m55),
    .Q(pp_row93_5));
 sky130_fd_sc_hd__dfxtp_1 _0844_ (.CLK(clknet_leaf_129_clk),
    .D(booth_b64_m55),
    .Q(pp_row119_5));
 sky130_fd_sc_hd__dfxtp_1 _0845_ (.CLK(clknet_leaf_105_clk),
    .D(booth_b40_m53),
    .Q(pp_row93_6));
 sky130_fd_sc_hd__dfxtp_1 _0846_ (.CLK(clknet_leaf_105_clk),
    .D(booth_b42_m51),
    .Q(pp_row93_7));
 sky130_fd_sc_hd__dfxtp_1 _0847_ (.CLK(clknet_leaf_105_clk),
    .D(booth_b44_m49),
    .Q(pp_row93_8));
 sky130_fd_sc_hd__dfxtp_1 _0848_ (.CLK(clknet_leaf_109_clk),
    .D(booth_b46_m47),
    .Q(pp_row93_9));
 sky130_fd_sc_hd__dfxtp_1 _0849_ (.CLK(clknet_leaf_109_clk),
    .D(booth_b48_m45),
    .Q(pp_row93_10));
 sky130_fd_sc_hd__dfxtp_1 _0850_ (.CLK(clknet_leaf_109_clk),
    .D(booth_b50_m43),
    .Q(pp_row93_11));
 sky130_fd_sc_hd__dfxtp_1 _0851_ (.CLK(clknet_leaf_144_clk),
    .D(booth_b52_m41),
    .Q(pp_row93_12));
 sky130_fd_sc_hd__dfxtp_1 _0852_ (.CLK(clknet_leaf_144_clk),
    .D(booth_b54_m39),
    .Q(pp_row93_13));
 sky130_fd_sc_hd__dfxtp_1 _0853_ (.CLK(clknet_leaf_144_clk),
    .D(booth_b56_m37),
    .Q(pp_row93_14));
 sky130_fd_sc_hd__dfxtp_1 _0854_ (.CLK(clknet_leaf_142_clk),
    .D(booth_b58_m35),
    .Q(pp_row93_15));
 sky130_fd_sc_hd__dfxtp_2 _0855_ (.CLK(clknet_leaf_181_clk),
    .D(net150),
    .Q(pp_row119_6));
 sky130_fd_sc_hd__dfxtp_1 _0856_ (.CLK(clknet_leaf_142_clk),
    .D(booth_b60_m33),
    .Q(pp_row93_16));
 sky130_fd_sc_hd__dfxtp_1 _0857_ (.CLK(clknet_leaf_142_clk),
    .D(booth_b62_m31),
    .Q(pp_row93_17));
 sky130_fd_sc_hd__dfxtp_1 _0858_ (.CLK(clknet_leaf_140_clk),
    .D(booth_b64_m29),
    .Q(pp_row93_18));
 sky130_fd_sc_hd__dfxtp_2 _0859_ (.CLK(clknet_leaf_194_clk),
    .D(net249),
    .Q(pp_row93_19));
 sky130_fd_sc_hd__dfxtp_1 _0860_ (.CLK(clknet_leaf_102_clk),
    .D(booth_b30_m64),
    .Q(pp_row94_1));
 sky130_fd_sc_hd__dfxtp_1 _0861_ (.CLK(clknet_leaf_102_clk),
    .D(booth_b32_m62),
    .Q(pp_row94_2));
 sky130_fd_sc_hd__dfxtp_1 _0862_ (.CLK(clknet_leaf_105_clk),
    .D(booth_b34_m60),
    .Q(pp_row94_3));
 sky130_fd_sc_hd__dfxtp_1 _0863_ (.CLK(clknet_leaf_105_clk),
    .D(booth_b36_m58),
    .Q(pp_row94_4));
 sky130_fd_sc_hd__dfxtp_1 _0864_ (.CLK(clknet_leaf_111_clk),
    .D(booth_b38_m56),
    .Q(pp_row94_5));
 sky130_fd_sc_hd__dfxtp_1 _0865_ (.CLK(clknet_leaf_111_clk),
    .D(booth_b40_m54),
    .Q(pp_row94_6));
 sky130_fd_sc_hd__dfxtp_1 _0866_ (.CLK(clknet_leaf_134_clk),
    .D(booth_b56_m64),
    .Q(pp_row120_1));
 sky130_fd_sc_hd__dfxtp_1 _0867_ (.CLK(clknet_leaf_111_clk),
    .D(booth_b42_m52),
    .Q(pp_row94_7));
 sky130_fd_sc_hd__dfxtp_1 _0868_ (.CLK(clknet_leaf_111_clk),
    .D(booth_b44_m50),
    .Q(pp_row94_8));
 sky130_fd_sc_hd__dfxtp_1 _0869_ (.CLK(clknet_leaf_104_clk),
    .D(booth_b46_m48),
    .Q(pp_row94_9));
 sky130_fd_sc_hd__dfxtp_1 _0870_ (.CLK(clknet_leaf_104_clk),
    .D(booth_b48_m46),
    .Q(pp_row94_10));
 sky130_fd_sc_hd__dfxtp_1 _0871_ (.CLK(clknet_leaf_141_clk),
    .D(booth_b50_m44),
    .Q(pp_row94_11));
 sky130_fd_sc_hd__dfxtp_1 _0872_ (.CLK(clknet_leaf_141_clk),
    .D(booth_b52_m42),
    .Q(pp_row94_12));
 sky130_fd_sc_hd__dfxtp_1 _0873_ (.CLK(clknet_leaf_141_clk),
    .D(booth_b54_m40),
    .Q(pp_row94_13));
 sky130_fd_sc_hd__dfxtp_1 _0874_ (.CLK(clknet_leaf_93_clk),
    .D(booth_b56_m38),
    .Q(pp_row94_14));
 sky130_fd_sc_hd__dfxtp_1 _0875_ (.CLK(clknet_leaf_93_clk),
    .D(booth_b58_m36),
    .Q(pp_row94_15));
 sky130_fd_sc_hd__dfxtp_1 _0876_ (.CLK(clknet_leaf_93_clk),
    .D(booth_b60_m34),
    .Q(pp_row94_16));
 sky130_fd_sc_hd__dfxtp_1 _0877_ (.CLK(clknet_leaf_133_clk),
    .D(booth_b58_m62),
    .Q(pp_row120_2));
 sky130_fd_sc_hd__dfxtp_1 _0878_ (.CLK(clknet_leaf_93_clk),
    .D(booth_b62_m32),
    .Q(pp_row94_17));
 sky130_fd_sc_hd__dfxtp_1 _0879_ (.CLK(clknet_leaf_93_clk),
    .D(booth_b64_m30),
    .Q(pp_row94_18));
 sky130_fd_sc_hd__dfxtp_2 _0880_ (.CLK(clknet_leaf_194_clk),
    .D(net250),
    .Q(pp_row94_19));
 sky130_fd_sc_hd__dfxtp_1 _0881_ (.CLK(clknet_leaf_111_clk),
    .D(\notsign$5524 ),
    .Q(pp_row95_0));
 sky130_fd_sc_hd__dfxtp_1 _0882_ (.CLK(clknet_leaf_110_clk),
    .D(booth_b32_m63),
    .Q(pp_row95_1));
 sky130_fd_sc_hd__dfxtp_1 _0883_ (.CLK(clknet_leaf_110_clk),
    .D(booth_b34_m61),
    .Q(pp_row95_2));
 sky130_fd_sc_hd__dfxtp_1 _0884_ (.CLK(clknet_leaf_100_clk),
    .D(booth_b36_m59),
    .Q(pp_row95_3));
 sky130_fd_sc_hd__dfxtp_1 _0885_ (.CLK(clknet_leaf_100_clk),
    .D(booth_b38_m57),
    .Q(pp_row95_4));
 sky130_fd_sc_hd__dfxtp_1 _0886_ (.CLK(clknet_leaf_100_clk),
    .D(booth_b40_m55),
    .Q(pp_row95_5));
 sky130_fd_sc_hd__dfxtp_1 _0887_ (.CLK(clknet_leaf_100_clk),
    .D(booth_b42_m53),
    .Q(pp_row95_6));
 sky130_fd_sc_hd__dfxtp_1 _0888_ (.CLK(clknet_leaf_130_clk),
    .D(booth_b60_m60),
    .Q(pp_row120_3));
 sky130_fd_sc_hd__dfxtp_1 _0889_ (.CLK(clknet_leaf_100_clk),
    .D(booth_b44_m51),
    .Q(pp_row95_7));
 sky130_fd_sc_hd__dfxtp_1 _0890_ (.CLK(clknet_leaf_100_clk),
    .D(booth_b46_m49),
    .Q(pp_row95_8));
 sky130_fd_sc_hd__dfxtp_1 _0891_ (.CLK(clknet_leaf_100_clk),
    .D(booth_b48_m47),
    .Q(pp_row95_9));
 sky130_fd_sc_hd__dfxtp_1 _0892_ (.CLK(clknet_leaf_100_clk),
    .D(booth_b50_m45),
    .Q(pp_row95_10));
 sky130_fd_sc_hd__dfxtp_1 _0893_ (.CLK(clknet_leaf_101_clk),
    .D(booth_b52_m43),
    .Q(pp_row95_11));
 sky130_fd_sc_hd__dfxtp_1 _0894_ (.CLK(clknet_leaf_100_clk),
    .D(booth_b54_m41),
    .Q(pp_row95_12));
 sky130_fd_sc_hd__dfxtp_1 _0895_ (.CLK(clknet_leaf_100_clk),
    .D(booth_b56_m39),
    .Q(pp_row95_13));
 sky130_fd_sc_hd__dfxtp_1 _0896_ (.CLK(clknet_leaf_100_clk),
    .D(booth_b58_m37),
    .Q(pp_row95_14));
 sky130_fd_sc_hd__dfxtp_1 _0897_ (.CLK(clknet_leaf_101_clk),
    .D(booth_b60_m35),
    .Q(pp_row95_15));
 sky130_fd_sc_hd__dfxtp_1 _0898_ (.CLK(clknet_leaf_101_clk),
    .D(booth_b62_m33),
    .Q(pp_row95_16));
 sky130_fd_sc_hd__dfxtp_1 _0899_ (.CLK(clknet_leaf_130_clk),
    .D(booth_b62_m58),
    .Q(pp_row120_4));
 sky130_fd_sc_hd__dfxtp_1 _0900_ (.CLK(clknet_leaf_101_clk),
    .D(booth_b64_m31),
    .Q(pp_row95_17));
 sky130_fd_sc_hd__dfxtp_4 _0901_ (.CLK(clknet_leaf_194_clk),
    .D(net251),
    .Q(pp_row95_18));
 sky130_fd_sc_hd__dfxtp_1 _0902_ (.CLK(clknet_leaf_102_clk),
    .D(booth_b32_m64),
    .Q(pp_row96_1));
 sky130_fd_sc_hd__dfxtp_1 _0903_ (.CLK(clknet_leaf_103_clk),
    .D(booth_b34_m62),
    .Q(pp_row96_2));
 sky130_fd_sc_hd__dfxtp_1 _0904_ (.CLK(clknet_leaf_103_clk),
    .D(booth_b36_m60),
    .Q(pp_row96_3));
 sky130_fd_sc_hd__dfxtp_1 _0905_ (.CLK(clknet_leaf_103_clk),
    .D(booth_b38_m58),
    .Q(pp_row96_4));
 sky130_fd_sc_hd__dfxtp_1 _0906_ (.CLK(clknet_leaf_103_clk),
    .D(booth_b40_m56),
    .Q(pp_row96_5));
 sky130_fd_sc_hd__dfxtp_1 _0907_ (.CLK(clknet_leaf_103_clk),
    .D(booth_b42_m54),
    .Q(pp_row96_6));
 sky130_fd_sc_hd__dfxtp_1 _0908_ (.CLK(clknet_leaf_103_clk),
    .D(booth_b44_m52),
    .Q(pp_row96_7));
 sky130_fd_sc_hd__dfxtp_1 _0909_ (.CLK(clknet_leaf_104_clk),
    .D(booth_b46_m50),
    .Q(pp_row96_8));
 sky130_fd_sc_hd__dfxtp_1 _0910_ (.CLK(clknet_leaf_133_clk),
    .D(booth_b64_m56),
    .Q(pp_row120_5));
 sky130_fd_sc_hd__dfxtp_1 _0911_ (.CLK(clknet_leaf_104_clk),
    .D(booth_b48_m48),
    .Q(pp_row96_9));
 sky130_fd_sc_hd__dfxtp_1 _0912_ (.CLK(clknet_leaf_104_clk),
    .D(booth_b50_m46),
    .Q(pp_row96_10));
 sky130_fd_sc_hd__dfxtp_1 _0913_ (.CLK(clknet_leaf_104_clk),
    .D(booth_b52_m44),
    .Q(pp_row96_11));
 sky130_fd_sc_hd__dfxtp_1 _0914_ (.CLK(clknet_leaf_104_clk),
    .D(booth_b54_m42),
    .Q(pp_row96_12));
 sky130_fd_sc_hd__dfxtp_1 _0915_ (.CLK(clknet_leaf_104_clk),
    .D(booth_b56_m40),
    .Q(pp_row96_13));
 sky130_fd_sc_hd__dfxtp_1 _0916_ (.CLK(clknet_leaf_103_clk),
    .D(booth_b58_m38),
    .Q(pp_row96_14));
 sky130_fd_sc_hd__dfxtp_1 _0917_ (.CLK(clknet_leaf_103_clk),
    .D(booth_b60_m36),
    .Q(pp_row96_15));
 sky130_fd_sc_hd__dfxtp_1 _0918_ (.CLK(clknet_leaf_104_clk),
    .D(booth_b62_m34),
    .Q(pp_row96_16));
 sky130_fd_sc_hd__dfxtp_1 _0919_ (.CLK(clknet_leaf_111_clk),
    .D(booth_b64_m32),
    .Q(pp_row96_17));
 sky130_fd_sc_hd__dfxtp_4 _0920_ (.CLK(clknet_leaf_185_clk),
    .D(net252),
    .Q(pp_row96_18));
 sky130_fd_sc_hd__dfxtp_2 _0921_ (.CLK(clknet_leaf_181_clk),
    .D(net152),
    .Q(pp_row120_6));
 sky130_fd_sc_hd__dfxtp_1 _0922_ (.CLK(clknet_leaf_112_clk),
    .D(\notsign$5594 ),
    .Q(pp_row97_0));
 sky130_fd_sc_hd__dfxtp_1 _0923_ (.CLK(clknet_leaf_112_clk),
    .D(booth_b34_m63),
    .Q(pp_row97_1));
 sky130_fd_sc_hd__dfxtp_1 _0924_ (.CLK(clknet_leaf_113_clk),
    .D(booth_b36_m61),
    .Q(pp_row97_2));
 sky130_fd_sc_hd__dfxtp_1 _0925_ (.CLK(clknet_leaf_112_clk),
    .D(booth_b38_m59),
    .Q(pp_row97_3));
 sky130_fd_sc_hd__dfxtp_1 _0926_ (.CLK(clknet_leaf_112_clk),
    .D(booth_b40_m57),
    .Q(pp_row97_4));
 sky130_fd_sc_hd__dfxtp_1 _0927_ (.CLK(clknet_leaf_112_clk),
    .D(booth_b42_m55),
    .Q(pp_row97_5));
 sky130_fd_sc_hd__dfxtp_1 _0928_ (.CLK(clknet_leaf_112_clk),
    .D(booth_b44_m53),
    .Q(pp_row97_6));
 sky130_fd_sc_hd__dfxtp_1 _0929_ (.CLK(clknet_leaf_112_clk),
    .D(booth_b46_m51),
    .Q(pp_row97_7));
 sky130_fd_sc_hd__dfxtp_1 _0930_ (.CLK(clknet_leaf_111_clk),
    .D(booth_b48_m49),
    .Q(pp_row97_8));
 sky130_fd_sc_hd__dfxtp_1 _0931_ (.CLK(clknet_leaf_112_clk),
    .D(booth_b50_m47),
    .Q(pp_row97_9));
 sky130_fd_sc_hd__dfxtp_1 _0932_ (.CLK(clknet_leaf_130_clk),
    .D(\notsign$6434 ),
    .Q(pp_row121_0));
 sky130_fd_sc_hd__dfxtp_1 _0933_ (.CLK(clknet_leaf_112_clk),
    .D(booth_b52_m45),
    .Q(pp_row97_10));
 sky130_fd_sc_hd__dfxtp_1 _0934_ (.CLK(clknet_leaf_112_clk),
    .D(booth_b54_m43),
    .Q(pp_row97_11));
 sky130_fd_sc_hd__dfxtp_1 _0935_ (.CLK(clknet_leaf_104_clk),
    .D(booth_b56_m41),
    .Q(pp_row97_12));
 sky130_fd_sc_hd__dfxtp_1 _0936_ (.CLK(clknet_leaf_104_clk),
    .D(booth_b58_m39),
    .Q(pp_row97_13));
 sky130_fd_sc_hd__dfxtp_1 _0937_ (.CLK(clknet_leaf_104_clk),
    .D(booth_b60_m37),
    .Q(pp_row97_14));
 sky130_fd_sc_hd__dfxtp_1 _0938_ (.CLK(clknet_leaf_113_clk),
    .D(booth_b62_m35),
    .Q(pp_row97_15));
 sky130_fd_sc_hd__dfxtp_1 _0939_ (.CLK(clknet_leaf_114_clk),
    .D(booth_b64_m33),
    .Q(pp_row97_16));
 sky130_fd_sc_hd__dfxtp_4 _0940_ (.CLK(clknet_leaf_184_clk),
    .D(net253),
    .Q(pp_row97_17));
 sky130_fd_sc_hd__dfxtp_1 _0941_ (.CLK(clknet_leaf_113_clk),
    .D(booth_b34_m64),
    .Q(pp_row98_1));
 sky130_fd_sc_hd__dfxtp_1 _0942_ (.CLK(clknet_leaf_113_clk),
    .D(booth_b36_m62),
    .Q(pp_row98_2));
 sky130_fd_sc_hd__dfxtp_1 _0943_ (.CLK(clknet_leaf_130_clk),
    .D(booth_b58_m63),
    .Q(pp_row121_1));
 sky130_fd_sc_hd__dfxtp_1 _0944_ (.CLK(clknet_leaf_180_clk),
    .D(booth_b64_m63),
    .Q(pp_row127_1));
 sky130_fd_sc_hd__dfxtp_1 _0945_ (.CLK(clknet_leaf_113_clk),
    .D(booth_b38_m60),
    .Q(pp_row98_3));
 sky130_fd_sc_hd__dfxtp_1 _0946_ (.CLK(clknet_leaf_113_clk),
    .D(booth_b40_m58),
    .Q(pp_row98_4));
 sky130_fd_sc_hd__dfxtp_1 _0947_ (.CLK(clknet_leaf_113_clk),
    .D(booth_b42_m56),
    .Q(pp_row98_5));
 sky130_fd_sc_hd__dfxtp_1 _0948_ (.CLK(clknet_leaf_113_clk),
    .D(booth_b44_m54),
    .Q(pp_row98_6));
 sky130_fd_sc_hd__dfxtp_1 _0949_ (.CLK(clknet_leaf_113_clk),
    .D(booth_b46_m52),
    .Q(pp_row98_7));
 sky130_fd_sc_hd__dfxtp_1 _0950_ (.CLK(clknet_leaf_114_clk),
    .D(booth_b48_m50),
    .Q(pp_row98_8));
 sky130_fd_sc_hd__dfxtp_1 _0951_ (.CLK(clknet_leaf_114_clk),
    .D(booth_b50_m48),
    .Q(pp_row98_9));
 sky130_fd_sc_hd__dfxtp_1 _0952_ (.CLK(clknet_leaf_114_clk),
    .D(booth_b52_m46),
    .Q(pp_row98_10));
 sky130_fd_sc_hd__dfxtp_1 _0953_ (.CLK(clknet_leaf_114_clk),
    .D(booth_b54_m44),
    .Q(pp_row98_11));
 sky130_fd_sc_hd__dfxtp_1 _0954_ (.CLK(clknet_leaf_116_clk),
    .D(booth_b56_m42),
    .Q(pp_row98_12));
 sky130_fd_sc_hd__dfxtp_1 _0955_ (.CLK(clknet_leaf_131_clk),
    .D(booth_b60_m61),
    .Q(pp_row121_2));
 sky130_fd_sc_hd__dfxtp_1 _0956_ (.CLK(clknet_leaf_116_clk),
    .D(booth_b58_m40),
    .Q(pp_row98_13));
 sky130_fd_sc_hd__dfxtp_1 _0957_ (.CLK(clknet_leaf_114_clk),
    .D(booth_b60_m38),
    .Q(pp_row98_14));
 sky130_fd_sc_hd__dfxtp_1 _0958_ (.CLK(clknet_leaf_114_clk),
    .D(booth_b62_m36),
    .Q(pp_row98_15));
 sky130_fd_sc_hd__dfxtp_1 _0959_ (.CLK(clknet_leaf_114_clk),
    .D(booth_b64_m34),
    .Q(pp_row98_16));
 sky130_fd_sc_hd__dfxtp_4 _0960_ (.CLK(clknet_leaf_185_clk),
    .D(net254),
    .Q(pp_row98_17));
 sky130_fd_sc_hd__dfxtp_1 _0961_ (.CLK(clknet_leaf_114_clk),
    .D(\notsign$5664 ),
    .Q(pp_row99_0));
 sky130_fd_sc_hd__dfxtp_1 _0962_ (.CLK(clknet_leaf_114_clk),
    .D(booth_b36_m63),
    .Q(pp_row99_1));
 sky130_fd_sc_hd__dfxtp_1 _0963_ (.CLK(clknet_leaf_114_clk),
    .D(booth_b38_m61),
    .Q(pp_row99_2));
 sky130_fd_sc_hd__dfxtp_1 _0964_ (.CLK(clknet_leaf_116_clk),
    .D(booth_b40_m59),
    .Q(pp_row99_3));
 sky130_fd_sc_hd__dfxtp_1 _0965_ (.CLK(clknet_leaf_116_clk),
    .D(booth_b42_m57),
    .Q(pp_row99_4));
 sky130_fd_sc_hd__dfxtp_1 _0966_ (.CLK(clknet_leaf_180_clk),
    .D(booth_b62_m59),
    .Q(pp_row121_3));
 sky130_fd_sc_hd__dfxtp_1 _0967_ (.CLK(clknet_leaf_116_clk),
    .D(booth_b44_m55),
    .Q(pp_row99_5));
 sky130_fd_sc_hd__dfxtp_1 _0968_ (.CLK(clknet_leaf_116_clk),
    .D(booth_b46_m53),
    .Q(pp_row99_6));
 sky130_fd_sc_hd__dfxtp_1 _0969_ (.CLK(clknet_leaf_116_clk),
    .D(booth_b48_m51),
    .Q(pp_row99_7));
 sky130_fd_sc_hd__dfxtp_1 _0970_ (.CLK(clknet_leaf_116_clk),
    .D(booth_b50_m49),
    .Q(pp_row99_8));
 sky130_fd_sc_hd__dfxtp_1 _0971_ (.CLK(clknet_leaf_117_clk),
    .D(booth_b52_m47),
    .Q(pp_row99_9));
 sky130_fd_sc_hd__dfxtp_1 _0972_ (.CLK(clknet_leaf_117_clk),
    .D(booth_b54_m45),
    .Q(pp_row99_10));
 sky130_fd_sc_hd__dfxtp_1 _0973_ (.CLK(clknet_leaf_117_clk),
    .D(booth_b56_m43),
    .Q(pp_row99_11));
 sky130_fd_sc_hd__dfxtp_1 _0974_ (.CLK(clknet_leaf_116_clk),
    .D(booth_b58_m41),
    .Q(pp_row99_12));
 sky130_fd_sc_hd__dfxtp_1 _0975_ (.CLK(clknet_leaf_116_clk),
    .D(booth_b60_m39),
    .Q(pp_row99_13));
 sky130_fd_sc_hd__dfxtp_1 _0976_ (.CLK(clknet_leaf_116_clk),
    .D(booth_b62_m37),
    .Q(pp_row99_14));
 sky130_fd_sc_hd__dfxtp_1 _0977_ (.CLK(clknet_leaf_180_clk),
    .D(booth_b64_m57),
    .Q(pp_row121_4));
 sky130_fd_sc_hd__dfxtp_1 _0978_ (.CLK(clknet_leaf_113_clk),
    .D(booth_b64_m35),
    .Q(pp_row99_15));
 sky130_fd_sc_hd__dfxtp_4 _0979_ (.CLK(clknet_leaf_184_clk),
    .D(net255),
    .Q(pp_row99_16));
 sky130_fd_sc_hd__dfxtp_1 _0980_ (.CLK(clknet_leaf_114_clk),
    .D(booth_b36_m64),
    .Q(pp_row100_1));
 sky130_fd_sc_hd__dfxtp_1 _0981_ (.CLK(clknet_leaf_114_clk),
    .D(booth_b38_m62),
    .Q(pp_row100_2));
 sky130_fd_sc_hd__dfxtp_1 _0982_ (.CLK(clknet_leaf_115_clk),
    .D(booth_b40_m60),
    .Q(pp_row100_3));
 sky130_fd_sc_hd__dfxtp_1 _0983_ (.CLK(clknet_leaf_118_clk),
    .D(booth_b42_m58),
    .Q(pp_row100_4));
 sky130_fd_sc_hd__dfxtp_1 _0984_ (.CLK(clknet_leaf_115_clk),
    .D(booth_b44_m56),
    .Q(pp_row100_5));
 sky130_fd_sc_hd__dfxtp_1 _0985_ (.CLK(clknet_leaf_117_clk),
    .D(booth_b46_m54),
    .Q(pp_row100_6));
 sky130_fd_sc_hd__dfxtp_1 _0986_ (.CLK(clknet_leaf_115_clk),
    .D(booth_b48_m52),
    .Q(pp_row100_7));
 sky130_fd_sc_hd__dfxtp_1 _0987_ (.CLK(clknet_leaf_115_clk),
    .D(booth_b50_m50),
    .Q(pp_row100_8));
 sky130_fd_sc_hd__dfxtp_1 _0988_ (.CLK(clknet_leaf_181_clk),
    .D(net153),
    .Q(pp_row121_5));
 sky130_fd_sc_hd__dfxtp_1 _0989_ (.CLK(clknet_leaf_118_clk),
    .D(booth_b52_m48),
    .Q(pp_row100_9));
 sky130_fd_sc_hd__dfxtp_1 _0990_ (.CLK(clknet_leaf_118_clk),
    .D(booth_b54_m46),
    .Q(pp_row100_10));
 sky130_fd_sc_hd__dfxtp_1 _0991_ (.CLK(clknet_leaf_118_clk),
    .D(booth_b56_m44),
    .Q(pp_row100_11));
 sky130_fd_sc_hd__dfxtp_1 _0992_ (.CLK(clknet_leaf_116_clk),
    .D(booth_b58_m42),
    .Q(pp_row100_12));
 sky130_fd_sc_hd__dfxtp_1 _0993_ (.CLK(clknet_leaf_116_clk),
    .D(booth_b60_m40),
    .Q(pp_row100_13));
 sky130_fd_sc_hd__dfxtp_1 _0994_ (.CLK(clknet_leaf_121_clk),
    .D(booth_b62_m38),
    .Q(pp_row100_14));
 sky130_fd_sc_hd__dfxtp_1 _0995_ (.CLK(clknet_leaf_110_clk),
    .D(booth_b64_m36),
    .Q(pp_row100_15));
 sky130_fd_sc_hd__dfxtp_4 _0996_ (.CLK(clknet_leaf_184_clk),
    .D(net130),
    .Q(pp_row100_16));
 sky130_fd_sc_hd__dfxtp_1 _0997_ (.CLK(clknet_leaf_119_clk),
    .D(\notsign$5734 ),
    .Q(pp_row101_0));
 sky130_fd_sc_hd__dfxtp_1 _0998_ (.CLK(clknet_leaf_118_clk),
    .D(booth_b38_m63),
    .Q(pp_row101_1));
 sky130_fd_sc_hd__dfxtp_1 _0999_ (.CLK(clknet_leaf_164_clk),
    .D(booth_b58_m64),
    .Q(pp_row122_1));
 sky130_fd_sc_hd__dfxtp_1 _1000_ (.CLK(clknet_leaf_119_clk),
    .D(booth_b40_m61),
    .Q(pp_row101_2));
 sky130_fd_sc_hd__dfxtp_1 _1001_ (.CLK(clknet_leaf_119_clk),
    .D(booth_b42_m59),
    .Q(pp_row101_3));
 sky130_fd_sc_hd__dfxtp_1 _1002_ (.CLK(clknet_leaf_118_clk),
    .D(booth_b44_m57),
    .Q(pp_row101_4));
 sky130_fd_sc_hd__dfxtp_1 _1003_ (.CLK(clknet_leaf_118_clk),
    .D(booth_b46_m55),
    .Q(pp_row101_5));
 sky130_fd_sc_hd__dfxtp_1 _1004_ (.CLK(clknet_leaf_117_clk),
    .D(booth_b48_m53),
    .Q(pp_row101_6));
 sky130_fd_sc_hd__dfxtp_1 _1005_ (.CLK(clknet_leaf_118_clk),
    .D(booth_b50_m51),
    .Q(pp_row101_7));
 sky130_fd_sc_hd__dfxtp_1 _1006_ (.CLK(clknet_leaf_117_clk),
    .D(booth_b52_m49),
    .Q(pp_row101_8));
 sky130_fd_sc_hd__dfxtp_1 _1007_ (.CLK(clknet_leaf_119_clk),
    .D(booth_b54_m47),
    .Q(pp_row101_9));
 sky130_fd_sc_hd__dfxtp_1 _1008_ (.CLK(clknet_leaf_117_clk),
    .D(booth_b56_m45),
    .Q(pp_row101_10));
 sky130_fd_sc_hd__dfxtp_1 _1009_ (.CLK(clknet_leaf_119_clk),
    .D(booth_b58_m43),
    .Q(pp_row101_11));
 sky130_fd_sc_hd__dfxtp_1 _1010_ (.CLK(clknet_leaf_129_clk),
    .D(booth_b60_m62),
    .Q(pp_row122_2));
 sky130_fd_sc_hd__dfxtp_1 _1011_ (.CLK(clknet_leaf_115_clk),
    .D(booth_b60_m41),
    .Q(pp_row101_12));
 sky130_fd_sc_hd__dfxtp_1 _1012_ (.CLK(clknet_leaf_115_clk),
    .D(booth_b62_m39),
    .Q(pp_row101_13));
 sky130_fd_sc_hd__dfxtp_1 _1013_ (.CLK(clknet_leaf_115_clk),
    .D(booth_b64_m37),
    .Q(pp_row101_14));
 sky130_fd_sc_hd__dfxtp_4 _1014_ (.CLK(clknet_leaf_182_clk),
    .D(net131),
    .Q(pp_row101_15));
 sky130_fd_sc_hd__dfxtp_1 _1015_ (.CLK(clknet_leaf_120_clk),
    .D(booth_b38_m64),
    .Q(pp_row102_1));
 sky130_fd_sc_hd__dfxtp_1 _1016_ (.CLK(clknet_leaf_120_clk),
    .D(booth_b40_m62),
    .Q(pp_row102_2));
 sky130_fd_sc_hd__dfxtp_1 _1017_ (.CLK(clknet_leaf_60_clk),
    .D(booth_b0_m0),
    .Q(pp_row0_0));
 sky130_fd_sc_hd__dfxtp_4 _1018_ (.CLK(clknet_leaf_60_clk),
    .D(net1574),
    .Q(pp_row0_1));
 sky130_fd_sc_hd__dfxtp_2 _1019_ (.CLK(clknet_leaf_249_clk),
    .D(net129),
    .Q(pp_row0_2));
 sky130_fd_sc_hd__dfxtp_1 _1020_ (.CLK(clknet_leaf_60_clk),
    .D(booth_b0_m1),
    .Q(pp_row1_0));
 sky130_fd_sc_hd__dfxtp_2 _1021_ (.CLK(clknet_leaf_249_clk),
    .D(net168),
    .Q(pp_row1_1));
 sky130_fd_sc_hd__dfxtp_1 _1022_ (.CLK(clknet_leaf_60_clk),
    .D(booth_b0_m2),
    .Q(pp_row2_0));
 sky130_fd_sc_hd__dfxtp_1 _1023_ (.CLK(clknet_leaf_60_clk),
    .D(booth_b2_m0),
    .Q(pp_row2_1));
 sky130_fd_sc_hd__dfxtp_1 _1024_ (.CLK(clknet_leaf_60_clk),
    .D(net1391),
    .Q(pp_row2_2));
 sky130_fd_sc_hd__dfxtp_4 _1025_ (.CLK(clknet_leaf_249_clk),
    .D(net179),
    .Q(pp_row2_3));
 sky130_fd_sc_hd__dfxtp_1 _1026_ (.CLK(clknet_leaf_61_clk),
    .D(booth_b0_m3),
    .Q(pp_row3_0));
 sky130_fd_sc_hd__dfxtp_1 _1027_ (.CLK(clknet_leaf_120_clk),
    .D(booth_b42_m60),
    .Q(pp_row102_3));
 sky130_fd_sc_hd__dfxtp_1 _1028_ (.CLK(clknet_leaf_61_clk),
    .D(booth_b2_m1),
    .Q(pp_row3_1));
 sky130_fd_sc_hd__dfxtp_4 _1029_ (.CLK(clknet_leaf_248_clk),
    .D(net190),
    .Q(pp_row3_2));
 sky130_fd_sc_hd__dfxtp_1 _1030_ (.CLK(clknet_leaf_61_clk),
    .D(booth_b0_m4),
    .Q(pp_row4_0));
 sky130_fd_sc_hd__dfxtp_1 _1031_ (.CLK(clknet_leaf_61_clk),
    .D(booth_b2_m2),
    .Q(pp_row4_1));
 sky130_fd_sc_hd__dfxtp_1 _1032_ (.CLK(clknet_leaf_60_clk),
    .D(booth_b4_m0),
    .Q(pp_row4_2));
 sky130_fd_sc_hd__dfxtp_1 _1033_ (.CLK(clknet_leaf_60_clk),
    .D(net1278),
    .Q(pp_row4_3));
 sky130_fd_sc_hd__dfxtp_4 _1034_ (.CLK(clknet_leaf_248_clk),
    .D(net201),
    .Q(pp_row4_4));
 sky130_fd_sc_hd__dfxtp_1 _1035_ (.CLK(clknet_leaf_61_clk),
    .D(booth_b0_m5),
    .Q(pp_row5_0));
 sky130_fd_sc_hd__dfxtp_1 _1036_ (.CLK(clknet_leaf_61_clk),
    .D(booth_b2_m3),
    .Q(pp_row5_1));
 sky130_fd_sc_hd__dfxtp_1 _1037_ (.CLK(clknet_leaf_60_clk),
    .D(booth_b4_m1),
    .Q(pp_row5_2));
 sky130_fd_sc_hd__dfxtp_1 _1038_ (.CLK(clknet_leaf_120_clk),
    .D(booth_b44_m58),
    .Q(pp_row102_4));
 sky130_fd_sc_hd__dfxtp_4 _1039_ (.CLK(clknet_leaf_248_clk),
    .D(net212),
    .Q(pp_row5_3));
 sky130_fd_sc_hd__dfxtp_1 _1040_ (.CLK(clknet_leaf_57_clk),
    .D(booth_b0_m6),
    .Q(pp_row6_0));
 sky130_fd_sc_hd__dfxtp_1 _1041_ (.CLK(clknet_leaf_57_clk),
    .D(booth_b2_m4),
    .Q(pp_row6_1));
 sky130_fd_sc_hd__dfxtp_1 _1042_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b4_m2),
    .Q(pp_row6_2));
 sky130_fd_sc_hd__dfxtp_1 _1043_ (.CLK(clknet_leaf_56_clk),
    .D(booth_b6_m0),
    .Q(pp_row6_3));
 sky130_fd_sc_hd__dfxtp_1 _1044_ (.CLK(clknet_leaf_56_clk),
    .D(net1249),
    .Q(pp_row6_4));
 sky130_fd_sc_hd__dfxtp_4 _1045_ (.CLK(clknet_leaf_248_clk),
    .D(net223),
    .Q(pp_row6_5));
 sky130_fd_sc_hd__dfxtp_1 _1046_ (.CLK(clknet_leaf_61_clk),
    .D(booth_b0_m7),
    .Q(pp_row7_0));
 sky130_fd_sc_hd__dfxtp_1 _1047_ (.CLK(clknet_leaf_61_clk),
    .D(booth_b2_m5),
    .Q(pp_row7_1));
 sky130_fd_sc_hd__dfxtp_1 _1048_ (.CLK(clknet_leaf_57_clk),
    .D(booth_b4_m3),
    .Q(pp_row7_2));
 sky130_fd_sc_hd__dfxtp_1 _1049_ (.CLK(clknet_leaf_120_clk),
    .D(booth_b46_m56),
    .Q(pp_row102_5));
 sky130_fd_sc_hd__dfxtp_1 _1050_ (.CLK(clknet_leaf_57_clk),
    .D(booth_b6_m1),
    .Q(pp_row7_3));
 sky130_fd_sc_hd__dfxtp_2 _1051_ (.CLK(clknet_leaf_248_clk),
    .D(net234),
    .Q(pp_row7_4));
 sky130_fd_sc_hd__dfxtp_1 _1052_ (.CLK(clknet_leaf_53_clk),
    .D(booth_b0_m8),
    .Q(pp_row8_0));
 sky130_fd_sc_hd__dfxtp_1 _1053_ (.CLK(clknet_leaf_53_clk),
    .D(booth_b2_m6),
    .Q(pp_row8_1));
 sky130_fd_sc_hd__dfxtp_1 _1054_ (.CLK(clknet_leaf_56_clk),
    .D(booth_b4_m4),
    .Q(pp_row8_2));
 sky130_fd_sc_hd__dfxtp_1 _1055_ (.CLK(clknet_leaf_58_clk),
    .D(booth_b6_m2),
    .Q(pp_row8_3));
 sky130_fd_sc_hd__dfxtp_1 _1056_ (.CLK(clknet_leaf_56_clk),
    .D(booth_b8_m0),
    .Q(pp_row8_4));
 sky130_fd_sc_hd__dfxtp_1 _1057_ (.CLK(clknet_leaf_58_clk),
    .D(net1240),
    .Q(pp_row8_5));
 sky130_fd_sc_hd__dfxtp_2 _1058_ (.CLK(clknet_leaf_248_clk),
    .D(net245),
    .Q(pp_row8_6));
 sky130_fd_sc_hd__dfxtp_1 _1059_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b0_m9),
    .Q(pp_row9_0));
 sky130_fd_sc_hd__dfxtp_1 _1060_ (.CLK(clknet_leaf_120_clk),
    .D(booth_b48_m54),
    .Q(pp_row102_6));
 sky130_fd_sc_hd__dfxtp_1 _1061_ (.CLK(clknet_leaf_129_clk),
    .D(booth_b62_m60),
    .Q(pp_row122_3));
 sky130_fd_sc_hd__dfxtp_1 _1062_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b2_m7),
    .Q(pp_row9_1));
 sky130_fd_sc_hd__dfxtp_1 _1063_ (.CLK(clknet_leaf_60_clk),
    .D(booth_b4_m5),
    .Q(pp_row9_2));
 sky130_fd_sc_hd__dfxtp_1 _1064_ (.CLK(clknet_leaf_59_clk),
    .D(booth_b6_m3),
    .Q(pp_row9_3));
 sky130_fd_sc_hd__dfxtp_1 _1065_ (.CLK(clknet_leaf_59_clk),
    .D(booth_b8_m1),
    .Q(pp_row9_4));
 sky130_fd_sc_hd__dfxtp_2 _1066_ (.CLK(clknet_leaf_248_clk),
    .D(net256),
    .Q(pp_row9_5));
 sky130_fd_sc_hd__dfxtp_1 _1067_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b0_m10),
    .Q(pp_row10_0));
 sky130_fd_sc_hd__dfxtp_1 _1068_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b2_m8),
    .Q(pp_row10_1));
 sky130_fd_sc_hd__dfxtp_1 _1069_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b4_m6),
    .Q(pp_row10_2));
 sky130_fd_sc_hd__dfxtp_1 _1070_ (.CLK(clknet_leaf_52_clk),
    .D(booth_b6_m4),
    .Q(pp_row10_3));
 sky130_fd_sc_hd__dfxtp_1 _1071_ (.CLK(clknet_leaf_52_clk),
    .D(booth_b8_m2),
    .Q(pp_row10_4));
 sky130_fd_sc_hd__dfxtp_1 _1072_ (.CLK(clknet_leaf_120_clk),
    .D(booth_b50_m52),
    .Q(pp_row102_7));
 sky130_fd_sc_hd__dfxtp_1 _1073_ (.CLK(clknet_leaf_52_clk),
    .D(booth_b10_m0),
    .Q(pp_row10_5));
 sky130_fd_sc_hd__dfxtp_1 _1074_ (.CLK(clknet_leaf_53_clk),
    .D(net1415),
    .Q(pp_row10_6));
 sky130_fd_sc_hd__dfxtp_2 _1075_ (.CLK(clknet_leaf_248_clk),
    .D(net140),
    .Q(pp_row10_7));
 sky130_fd_sc_hd__dfxtp_1 _1076_ (.CLK(clknet_leaf_52_clk),
    .D(booth_b0_m11),
    .Q(pp_row11_0));
 sky130_fd_sc_hd__dfxtp_1 _1077_ (.CLK(clknet_leaf_52_clk),
    .D(booth_b2_m9),
    .Q(pp_row11_1));
 sky130_fd_sc_hd__dfxtp_1 _1078_ (.CLK(clknet_leaf_52_clk),
    .D(booth_b4_m7),
    .Q(pp_row11_2));
 sky130_fd_sc_hd__dfxtp_1 _1079_ (.CLK(clknet_leaf_52_clk),
    .D(booth_b6_m5),
    .Q(pp_row11_3));
 sky130_fd_sc_hd__dfxtp_1 _1080_ (.CLK(clknet_leaf_52_clk),
    .D(booth_b8_m3),
    .Q(pp_row11_4));
 sky130_fd_sc_hd__dfxtp_1 _1081_ (.CLK(clknet_leaf_53_clk),
    .D(booth_b10_m1),
    .Q(pp_row11_5));
 sky130_fd_sc_hd__dfxtp_2 _1082_ (.CLK(clknet_leaf_248_clk),
    .D(net151),
    .Q(pp_row11_6));
 sky130_fd_sc_hd__dfxtp_1 _1083_ (.CLK(clknet_leaf_120_clk),
    .D(booth_b52_m50),
    .Q(pp_row102_8));
 sky130_fd_sc_hd__dfxtp_1 _1084_ (.CLK(clknet_leaf_58_clk),
    .D(booth_b0_m12),
    .Q(pp_row12_0));
 sky130_fd_sc_hd__dfxtp_1 _1085_ (.CLK(clknet_leaf_58_clk),
    .D(booth_b2_m10),
    .Q(pp_row12_1));
 sky130_fd_sc_hd__dfxtp_1 _1086_ (.CLK(clknet_leaf_58_clk),
    .D(booth_b4_m8),
    .Q(pp_row12_2));
 sky130_fd_sc_hd__dfxtp_1 _1087_ (.CLK(clknet_leaf_58_clk),
    .D(booth_b6_m6),
    .Q(pp_row12_3));
 sky130_fd_sc_hd__dfxtp_1 _1088_ (.CLK(clknet_leaf_58_clk),
    .D(booth_b8_m4),
    .Q(pp_row12_4));
 sky130_fd_sc_hd__dfxtp_1 _1089_ (.CLK(clknet_leaf_59_clk),
    .D(booth_b10_m2),
    .Q(pp_row12_5));
 sky130_fd_sc_hd__dfxtp_1 _1090_ (.CLK(clknet_leaf_58_clk),
    .D(booth_b12_m0),
    .Q(pp_row12_6));
 sky130_fd_sc_hd__dfxtp_1 _1091_ (.CLK(clknet_leaf_59_clk),
    .D(net1313),
    .Q(pp_row12_7));
 sky130_fd_sc_hd__dfxtp_2 _1092_ (.CLK(clknet_leaf_248_clk),
    .D(net160),
    .Q(pp_row12_8));
 sky130_fd_sc_hd__dfxtp_1 _1093_ (.CLK(clknet_leaf_59_clk),
    .D(booth_b0_m13),
    .Q(pp_row13_0));
 sky130_fd_sc_hd__dfxtp_1 _1094_ (.CLK(clknet_leaf_121_clk),
    .D(booth_b54_m48),
    .Q(pp_row102_9));
 sky130_fd_sc_hd__dfxtp_1 _1095_ (.CLK(clknet_leaf_59_clk),
    .D(booth_b2_m11),
    .Q(pp_row13_1));
 sky130_fd_sc_hd__dfxtp_1 _1096_ (.CLK(clknet_leaf_60_clk),
    .D(booth_b4_m9),
    .Q(pp_row13_2));
 sky130_fd_sc_hd__dfxtp_1 _1097_ (.CLK(clknet_leaf_59_clk),
    .D(booth_b6_m7),
    .Q(pp_row13_3));
 sky130_fd_sc_hd__dfxtp_1 _1098_ (.CLK(clknet_leaf_59_clk),
    .D(booth_b8_m5),
    .Q(pp_row13_4));
 sky130_fd_sc_hd__dfxtp_1 _1099_ (.CLK(clknet_leaf_52_clk),
    .D(booth_b10_m3),
    .Q(pp_row13_5));
 sky130_fd_sc_hd__dfxtp_1 _1100_ (.CLK(clknet_leaf_52_clk),
    .D(booth_b12_m1),
    .Q(pp_row13_6));
 sky130_fd_sc_hd__dfxtp_2 _1101_ (.CLK(clknet_leaf_248_clk),
    .D(net161),
    .Q(pp_row13_7));
 sky130_fd_sc_hd__dfxtp_1 _1102_ (.CLK(clknet_leaf_14_clk),
    .D(booth_b0_m14),
    .Q(pp_row14_0));
 sky130_fd_sc_hd__dfxtp_1 _1103_ (.CLK(clknet_leaf_14_clk),
    .D(booth_b2_m12),
    .Q(pp_row14_1));
 sky130_fd_sc_hd__dfxtp_1 _1104_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b4_m10),
    .Q(pp_row14_2));
 sky130_fd_sc_hd__dfxtp_1 _1105_ (.CLK(clknet_leaf_121_clk),
    .D(booth_b56_m46),
    .Q(pp_row102_10));
 sky130_fd_sc_hd__dfxtp_1 _1106_ (.CLK(clknet_leaf_14_clk),
    .D(booth_b6_m8),
    .Q(pp_row14_3));
 sky130_fd_sc_hd__dfxtp_1 _1107_ (.CLK(clknet_leaf_14_clk),
    .D(booth_b8_m6),
    .Q(pp_row14_4));
 sky130_fd_sc_hd__dfxtp_1 _1108_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b10_m4),
    .Q(pp_row14_5));
 sky130_fd_sc_hd__dfxtp_1 _1109_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b12_m2),
    .Q(pp_row14_6));
 sky130_fd_sc_hd__dfxtp_1 _1110_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b14_m0),
    .Q(pp_row14_7));
 sky130_fd_sc_hd__dfxtp_1 _1111_ (.CLK(clknet_leaf_15_clk),
    .D(net1185),
    .Q(pp_row14_8));
 sky130_fd_sc_hd__dfxtp_2 _1112_ (.CLK(clknet_leaf_248_clk),
    .D(net162),
    .Q(pp_row14_9));
 sky130_fd_sc_hd__dfxtp_1 _1113_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b0_m15),
    .Q(pp_row15_0));
 sky130_fd_sc_hd__dfxtp_1 _1114_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b2_m13),
    .Q(pp_row15_1));
 sky130_fd_sc_hd__dfxtp_1 _1115_ (.CLK(clknet_leaf_47_clk),
    .D(booth_b4_m11),
    .Q(pp_row15_2));
 sky130_fd_sc_hd__dfxtp_1 _1116_ (.CLK(clknet_leaf_121_clk),
    .D(booth_b58_m44),
    .Q(pp_row102_11));
 sky130_fd_sc_hd__dfxtp_1 _1117_ (.CLK(clknet_leaf_47_clk),
    .D(booth_b6_m9),
    .Q(pp_row15_3));
 sky130_fd_sc_hd__dfxtp_1 _1118_ (.CLK(clknet_leaf_14_clk),
    .D(booth_b8_m7),
    .Q(pp_row15_4));
 sky130_fd_sc_hd__dfxtp_1 _1119_ (.CLK(clknet_leaf_48_clk),
    .D(booth_b10_m5),
    .Q(pp_row15_5));
 sky130_fd_sc_hd__dfxtp_1 _1120_ (.CLK(clknet_leaf_48_clk),
    .D(booth_b12_m3),
    .Q(pp_row15_6));
 sky130_fd_sc_hd__dfxtp_1 _1121_ (.CLK(clknet_leaf_48_clk),
    .D(booth_b14_m1),
    .Q(pp_row15_7));
 sky130_fd_sc_hd__dfxtp_2 _1122_ (.CLK(clknet_leaf_248_clk),
    .D(net163),
    .Q(pp_row15_8));
 sky130_fd_sc_hd__dfxtp_1 _1123_ (.CLK(clknet_leaf_11_clk),
    .D(booth_b0_m16),
    .Q(pp_row16_0));
 sky130_fd_sc_hd__dfxtp_1 _1124_ (.CLK(clknet_leaf_11_clk),
    .D(booth_b2_m14),
    .Q(pp_row16_1));
 sky130_fd_sc_hd__dfxtp_1 _1125_ (.CLK(clknet_leaf_11_clk),
    .D(booth_b4_m12),
    .Q(pp_row16_2));
 sky130_fd_sc_hd__dfxtp_1 _1126_ (.CLK(clknet_leaf_12_clk),
    .D(booth_b6_m10),
    .Q(pp_row16_3));
 sky130_fd_sc_hd__dfxtp_1 _1127_ (.CLK(clknet_leaf_119_clk),
    .D(booth_b60_m42),
    .Q(pp_row102_12));
 sky130_fd_sc_hd__dfxtp_1 _1128_ (.CLK(clknet_leaf_12_clk),
    .D(booth_b8_m8),
    .Q(pp_row16_4));
 sky130_fd_sc_hd__dfxtp_1 _1129_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b10_m6),
    .Q(pp_row16_5));
 sky130_fd_sc_hd__dfxtp_1 _1130_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b12_m4),
    .Q(pp_row16_6));
 sky130_fd_sc_hd__dfxtp_1 _1131_ (.CLK(clknet_leaf_11_clk),
    .D(booth_b14_m2),
    .Q(pp_row16_7));
 sky130_fd_sc_hd__dfxtp_1 _1132_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b16_m0),
    .Q(pp_row16_8));
 sky130_fd_sc_hd__dfxtp_1 _1133_ (.CLK(clknet_leaf_13_clk),
    .D(net1008),
    .Q(pp_row16_9));
 sky130_fd_sc_hd__dfxtp_1 _1134_ (.CLK(clknet_leaf_247_clk),
    .D(net164),
    .Q(pp_row16_10));
 sky130_fd_sc_hd__dfxtp_1 _1135_ (.CLK(clknet_leaf_16_clk),
    .D(booth_b0_m17),
    .Q(pp_row17_0));
 sky130_fd_sc_hd__dfxtp_1 _1136_ (.CLK(clknet_leaf_16_clk),
    .D(booth_b2_m15),
    .Q(pp_row17_1));
 sky130_fd_sc_hd__dfxtp_1 _1137_ (.CLK(clknet_leaf_16_clk),
    .D(booth_b4_m13),
    .Q(pp_row17_2));
 sky130_fd_sc_hd__dfxtp_1 _1138_ (.CLK(clknet_leaf_119_clk),
    .D(booth_b62_m40),
    .Q(pp_row102_13));
 sky130_fd_sc_hd__dfxtp_1 _1139_ (.CLK(clknet_leaf_16_clk),
    .D(booth_b6_m11),
    .Q(pp_row17_3));
 sky130_fd_sc_hd__dfxtp_1 _1140_ (.CLK(clknet_leaf_15_clk),
    .D(booth_b8_m9),
    .Q(pp_row17_4));
 sky130_fd_sc_hd__dfxtp_1 _1141_ (.CLK(clknet_leaf_11_clk),
    .D(booth_b10_m7),
    .Q(pp_row17_5));
 sky130_fd_sc_hd__dfxtp_1 _1142_ (.CLK(clknet_leaf_11_clk),
    .D(booth_b12_m5),
    .Q(pp_row17_6));
 sky130_fd_sc_hd__dfxtp_1 _1143_ (.CLK(clknet_leaf_11_clk),
    .D(booth_b14_m3),
    .Q(pp_row17_7));
 sky130_fd_sc_hd__dfxtp_1 _1144_ (.CLK(clknet_leaf_11_clk),
    .D(booth_b16_m1),
    .Q(pp_row17_8));
 sky130_fd_sc_hd__dfxtp_2 _1145_ (.CLK(clknet_leaf_245_clk),
    .D(net165),
    .Q(pp_row17_9));
 sky130_fd_sc_hd__dfxtp_1 _1146_ (.CLK(clknet_leaf_15_clk),
    .D(booth_b0_m18),
    .Q(pp_row18_0));
 sky130_fd_sc_hd__dfxtp_1 _1147_ (.CLK(clknet_leaf_15_clk),
    .D(booth_b2_m16),
    .Q(pp_row18_1));
 sky130_fd_sc_hd__dfxtp_1 _1148_ (.CLK(clknet_leaf_15_clk),
    .D(booth_b4_m14),
    .Q(pp_row18_2));
 sky130_fd_sc_hd__dfxtp_1 _1149_ (.CLK(clknet_leaf_119_clk),
    .D(booth_b64_m38),
    .Q(pp_row102_14));
 sky130_fd_sc_hd__dfxtp_1 _1150_ (.CLK(clknet_leaf_14_clk),
    .D(booth_b6_m12),
    .Q(pp_row18_3));
 sky130_fd_sc_hd__dfxtp_1 _1151_ (.CLK(clknet_leaf_15_clk),
    .D(booth_b8_m10),
    .Q(pp_row18_4));
 sky130_fd_sc_hd__dfxtp_1 _1152_ (.CLK(clknet_leaf_15_clk),
    .D(booth_b10_m8),
    .Q(pp_row18_5));
 sky130_fd_sc_hd__dfxtp_1 _1153_ (.CLK(clknet_leaf_15_clk),
    .D(booth_b12_m6),
    .Q(pp_row18_6));
 sky130_fd_sc_hd__dfxtp_1 _1154_ (.CLK(clknet_leaf_47_clk),
    .D(booth_b14_m4),
    .Q(pp_row18_7));
 sky130_fd_sc_hd__dfxtp_1 _1155_ (.CLK(clknet_leaf_15_clk),
    .D(booth_b16_m2),
    .Q(pp_row18_8));
 sky130_fd_sc_hd__dfxtp_1 _1156_ (.CLK(clknet_leaf_15_clk),
    .D(booth_b18_m0),
    .Q(pp_row18_9));
 sky130_fd_sc_hd__dfxtp_1 _1157_ (.CLK(clknet_leaf_15_clk),
    .D(net1664),
    .Q(pp_row18_10));
 sky130_fd_sc_hd__dfxtp_2 _1158_ (.CLK(clknet_leaf_245_clk),
    .D(net166),
    .Q(pp_row18_11));
 sky130_fd_sc_hd__dfxtp_1 _1159_ (.CLK(clknet_leaf_46_clk),
    .D(booth_b0_m19),
    .Q(pp_row19_0));
 sky130_fd_sc_hd__dfxtp_4 _1160_ (.CLK(clknet_leaf_182_clk),
    .D(net132),
    .Q(pp_row102_15));
 sky130_fd_sc_hd__dfxtp_1 _1161_ (.CLK(clknet_leaf_46_clk),
    .D(booth_b2_m17),
    .Q(pp_row19_1));
 sky130_fd_sc_hd__dfxtp_1 _1162_ (.CLK(clknet_leaf_46_clk),
    .D(booth_b4_m15),
    .Q(pp_row19_2));
 sky130_fd_sc_hd__dfxtp_1 _1163_ (.CLK(clknet_leaf_50_clk),
    .D(booth_b6_m13),
    .Q(pp_row19_3));
 sky130_fd_sc_hd__dfxtp_1 _1164_ (.CLK(clknet_leaf_50_clk),
    .D(booth_b8_m11),
    .Q(pp_row19_4));
 sky130_fd_sc_hd__dfxtp_1 _1165_ (.CLK(clknet_leaf_50_clk),
    .D(booth_b10_m9),
    .Q(pp_row19_5));
 sky130_fd_sc_hd__dfxtp_1 _1166_ (.CLK(clknet_leaf_46_clk),
    .D(booth_b12_m7),
    .Q(pp_row19_6));
 sky130_fd_sc_hd__dfxtp_1 _1167_ (.CLK(clknet_leaf_45_clk),
    .D(booth_b14_m5),
    .Q(pp_row19_7));
 sky130_fd_sc_hd__dfxtp_1 _1168_ (.CLK(clknet_leaf_46_clk),
    .D(booth_b16_m3),
    .Q(pp_row19_8));
 sky130_fd_sc_hd__dfxtp_1 _1169_ (.CLK(clknet_leaf_47_clk),
    .D(booth_b18_m1),
    .Q(pp_row19_9));
 sky130_fd_sc_hd__dfxtp_2 _1170_ (.CLK(clknet_leaf_247_clk),
    .D(net167),
    .Q(pp_row19_10));
 sky130_fd_sc_hd__dfxtp_1 _1171_ (.CLK(clknet_leaf_125_clk),
    .D(\notsign$5804 ),
    .Q(pp_row103_0));
 sky130_fd_sc_hd__dfxtp_1 _1172_ (.CLK(clknet_leaf_129_clk),
    .D(booth_b64_m58),
    .Q(pp_row122_4));
 sky130_fd_sc_hd__dfxtp_1 _1173_ (.CLK(clknet_leaf_46_clk),
    .D(booth_b0_m20),
    .Q(pp_row20_0));
 sky130_fd_sc_hd__dfxtp_1 _1174_ (.CLK(clknet_leaf_46_clk),
    .D(booth_b2_m18),
    .Q(pp_row20_1));
 sky130_fd_sc_hd__dfxtp_1 _1175_ (.CLK(clknet_leaf_45_clk),
    .D(booth_b4_m16),
    .Q(pp_row20_2));
 sky130_fd_sc_hd__dfxtp_1 _1176_ (.CLK(clknet_leaf_50_clk),
    .D(booth_b6_m14),
    .Q(pp_row20_3));
 sky130_fd_sc_hd__dfxtp_1 _1177_ (.CLK(clknet_leaf_50_clk),
    .D(booth_b8_m12),
    .Q(pp_row20_4));
 sky130_fd_sc_hd__dfxtp_1 _1178_ (.CLK(clknet_leaf_50_clk),
    .D(booth_b10_m10),
    .Q(pp_row20_5));
 sky130_fd_sc_hd__dfxtp_1 _1179_ (.CLK(clknet_leaf_49_clk),
    .D(booth_b12_m8),
    .Q(pp_row20_6));
 sky130_fd_sc_hd__dfxtp_1 _1180_ (.CLK(clknet_leaf_49_clk),
    .D(booth_b14_m6),
    .Q(pp_row20_7));
 sky130_fd_sc_hd__dfxtp_1 _1181_ (.CLK(clknet_leaf_49_clk),
    .D(booth_b16_m4),
    .Q(pp_row20_8));
 sky130_fd_sc_hd__dfxtp_1 _1182_ (.CLK(clknet_leaf_53_clk),
    .D(booth_b18_m2),
    .Q(pp_row20_9));
 sky130_fd_sc_hd__dfxtp_1 _1183_ (.CLK(clknet_leaf_124_clk),
    .D(booth_b40_m63),
    .Q(pp_row103_1));
 sky130_fd_sc_hd__dfxtp_1 _1184_ (.CLK(clknet_leaf_53_clk),
    .D(booth_b20_m0),
    .Q(pp_row20_10));
 sky130_fd_sc_hd__dfxtp_1 _1185_ (.CLK(clknet_leaf_46_clk),
    .D(net1487),
    .Q(pp_row20_11));
 sky130_fd_sc_hd__dfxtp_2 _1186_ (.CLK(clknet_leaf_244_clk),
    .D(net169),
    .Q(pp_row20_12));
 sky130_fd_sc_hd__dfxtp_1 _1187_ (.CLK(clknet_leaf_49_clk),
    .D(booth_b0_m21),
    .Q(pp_row21_0));
 sky130_fd_sc_hd__dfxtp_1 _1188_ (.CLK(clknet_leaf_49_clk),
    .D(booth_b2_m19),
    .Q(pp_row21_1));
 sky130_fd_sc_hd__dfxtp_1 _1189_ (.CLK(clknet_leaf_49_clk),
    .D(booth_b4_m17),
    .Q(pp_row21_2));
 sky130_fd_sc_hd__dfxtp_1 _1190_ (.CLK(clknet_leaf_59_clk),
    .D(booth_b6_m15),
    .Q(pp_row21_3));
 sky130_fd_sc_hd__dfxtp_1 _1191_ (.CLK(clknet_leaf_59_clk),
    .D(booth_b8_m13),
    .Q(pp_row21_4));
 sky130_fd_sc_hd__dfxtp_1 _1192_ (.CLK(clknet_leaf_52_clk),
    .D(booth_b10_m11),
    .Q(pp_row21_5));
 sky130_fd_sc_hd__dfxtp_1 _1193_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b12_m9),
    .Q(pp_row21_6));
 sky130_fd_sc_hd__dfxtp_1 _1194_ (.CLK(clknet_leaf_124_clk),
    .D(booth_b42_m61),
    .Q(pp_row103_2));
 sky130_fd_sc_hd__dfxtp_1 _1195_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b14_m7),
    .Q(pp_row21_7));
 sky130_fd_sc_hd__dfxtp_1 _1196_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b16_m5),
    .Q(pp_row21_8));
 sky130_fd_sc_hd__dfxtp_1 _1197_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b18_m3),
    .Q(pp_row21_9));
 sky130_fd_sc_hd__dfxtp_1 _1198_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b20_m1),
    .Q(pp_row21_10));
 sky130_fd_sc_hd__dfxtp_2 _1199_ (.CLK(clknet_leaf_245_clk),
    .D(net170),
    .Q(pp_row21_11));
 sky130_fd_sc_hd__dfxtp_1 _1200_ (.CLK(clknet_leaf_49_clk),
    .D(booth_b0_m22),
    .Q(pp_row22_0));
 sky130_fd_sc_hd__dfxtp_1 _1201_ (.CLK(clknet_leaf_49_clk),
    .D(booth_b2_m20),
    .Q(pp_row22_1));
 sky130_fd_sc_hd__dfxtp_1 _1202_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b4_m18),
    .Q(pp_row22_2));
 sky130_fd_sc_hd__dfxtp_1 _1203_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b6_m16),
    .Q(pp_row22_3));
 sky130_fd_sc_hd__dfxtp_1 _1204_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b8_m14),
    .Q(pp_row22_4));
 sky130_fd_sc_hd__dfxtp_1 _1205_ (.CLK(clknet_leaf_143_clk),
    .D(booth_b44_m59),
    .Q(pp_row103_3));
 sky130_fd_sc_hd__dfxtp_1 _1206_ (.CLK(clknet_leaf_47_clk),
    .D(booth_b10_m12),
    .Q(pp_row22_5));
 sky130_fd_sc_hd__dfxtp_1 _1207_ (.CLK(clknet_leaf_47_clk),
    .D(booth_b12_m10),
    .Q(pp_row22_6));
 sky130_fd_sc_hd__dfxtp_1 _1208_ (.CLK(clknet_leaf_47_clk),
    .D(booth_b14_m8),
    .Q(pp_row22_7));
 sky130_fd_sc_hd__dfxtp_1 _1209_ (.CLK(clknet_leaf_49_clk),
    .D(booth_b16_m6),
    .Q(pp_row22_8));
 sky130_fd_sc_hd__dfxtp_1 _1210_ (.CLK(clknet_leaf_49_clk),
    .D(booth_b18_m4),
    .Q(pp_row22_9));
 sky130_fd_sc_hd__dfxtp_1 _1211_ (.CLK(clknet_leaf_49_clk),
    .D(booth_b20_m2),
    .Q(pp_row22_10));
 sky130_fd_sc_hd__dfxtp_1 _1212_ (.CLK(clknet_leaf_49_clk),
    .D(booth_b22_m0),
    .Q(pp_row22_11));
 sky130_fd_sc_hd__dfxtp_1 _1213_ (.CLK(clknet_leaf_49_clk),
    .D(net1478),
    .Q(pp_row22_12));
 sky130_fd_sc_hd__dfxtp_2 _1214_ (.CLK(clknet_leaf_245_clk),
    .D(net171),
    .Q(pp_row22_13));
 sky130_fd_sc_hd__dfxtp_1 _1215_ (.CLK(clknet_leaf_47_clk),
    .D(booth_b0_m23),
    .Q(pp_row23_0));
 sky130_fd_sc_hd__dfxtp_1 _1216_ (.CLK(clknet_leaf_143_clk),
    .D(booth_b46_m57),
    .Q(pp_row103_4));
 sky130_fd_sc_hd__dfxtp_1 _1217_ (.CLK(clknet_leaf_47_clk),
    .D(booth_b2_m21),
    .Q(pp_row23_1));
 sky130_fd_sc_hd__dfxtp_1 _1218_ (.CLK(clknet_leaf_48_clk),
    .D(booth_b4_m19),
    .Q(pp_row23_2));
 sky130_fd_sc_hd__dfxtp_1 _1219_ (.CLK(clknet_leaf_48_clk),
    .D(booth_b6_m17),
    .Q(pp_row23_3));
 sky130_fd_sc_hd__dfxtp_1 _1220_ (.CLK(clknet_leaf_48_clk),
    .D(booth_b8_m15),
    .Q(pp_row23_4));
 sky130_fd_sc_hd__dfxtp_1 _1221_ (.CLK(clknet_leaf_48_clk),
    .D(booth_b10_m13),
    .Q(pp_row23_5));
 sky130_fd_sc_hd__dfxtp_1 _1222_ (.CLK(clknet_leaf_48_clk),
    .D(booth_b12_m11),
    .Q(pp_row23_6));
 sky130_fd_sc_hd__dfxtp_1 _1223_ (.CLK(clknet_leaf_48_clk),
    .D(booth_b14_m9),
    .Q(pp_row23_7));
 sky130_fd_sc_hd__dfxtp_1 _1224_ (.CLK(clknet_leaf_48_clk),
    .D(booth_b16_m7),
    .Q(pp_row23_8));
 sky130_fd_sc_hd__dfxtp_1 _1225_ (.CLK(clknet_leaf_48_clk),
    .D(booth_b18_m5),
    .Q(pp_row23_9));
 sky130_fd_sc_hd__dfxtp_1 _1226_ (.CLK(clknet_leaf_48_clk),
    .D(booth_b20_m3),
    .Q(pp_row23_10));
 sky130_fd_sc_hd__dfxtp_1 _1227_ (.CLK(clknet_leaf_143_clk),
    .D(booth_b48_m55),
    .Q(pp_row103_5));
 sky130_fd_sc_hd__dfxtp_1 _1228_ (.CLK(clknet_leaf_49_clk),
    .D(booth_b22_m1),
    .Q(pp_row23_11));
 sky130_fd_sc_hd__dfxtp_2 _1229_ (.CLK(clknet_leaf_244_clk),
    .D(net172),
    .Q(pp_row23_12));
 sky130_fd_sc_hd__dfxtp_1 _1230_ (.CLK(clknet_leaf_12_clk),
    .D(booth_b0_m24),
    .Q(pp_row24_0));
 sky130_fd_sc_hd__dfxtp_1 _1231_ (.CLK(clknet_leaf_12_clk),
    .D(booth_b2_m22),
    .Q(pp_row24_1));
 sky130_fd_sc_hd__dfxtp_1 _1232_ (.CLK(clknet_leaf_12_clk),
    .D(booth_b4_m20),
    .Q(pp_row24_2));
 sky130_fd_sc_hd__dfxtp_1 _1233_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b6_m18),
    .Q(pp_row24_3));
 sky130_fd_sc_hd__dfxtp_1 _1234_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b8_m16),
    .Q(pp_row24_4));
 sky130_fd_sc_hd__dfxtp_1 _1235_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b10_m14),
    .Q(pp_row24_5));
 sky130_fd_sc_hd__dfxtp_1 _1236_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b12_m12),
    .Q(pp_row24_6));
 sky130_fd_sc_hd__dfxtp_1 _1237_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b14_m10),
    .Q(pp_row24_7));
 sky130_fd_sc_hd__dfxtp_1 _1238_ (.CLK(clknet_leaf_109_clk),
    .D(booth_b50_m53),
    .Q(pp_row103_6));
 sky130_fd_sc_hd__dfxtp_1 _1239_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b16_m8),
    .Q(pp_row24_8));
 sky130_fd_sc_hd__dfxtp_1 _1240_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b18_m6),
    .Q(pp_row24_9));
 sky130_fd_sc_hd__dfxtp_1 _1241_ (.CLK(clknet_leaf_13_clk),
    .D(booth_b20_m4),
    .Q(pp_row24_10));
 sky130_fd_sc_hd__dfxtp_1 _1242_ (.CLK(clknet_leaf_15_clk),
    .D(booth_b22_m2),
    .Q(pp_row24_11));
 sky130_fd_sc_hd__dfxtp_1 _1243_ (.CLK(clknet_leaf_15_clk),
    .D(booth_b24_m0),
    .Q(pp_row24_12));
 sky130_fd_sc_hd__dfxtp_1 _1244_ (.CLK(clknet_leaf_14_clk),
    .D(net1467),
    .Q(pp_row24_13));
 sky130_fd_sc_hd__dfxtp_2 _1245_ (.CLK(clknet_leaf_244_clk),
    .D(net173),
    .Q(pp_row24_14));
 sky130_fd_sc_hd__dfxtp_1 _1246_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b0_m25),
    .Q(pp_row25_0));
 sky130_fd_sc_hd__dfxtp_1 _1247_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b2_m23),
    .Q(pp_row25_1));
 sky130_fd_sc_hd__dfxtp_1 _1248_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b4_m21),
    .Q(pp_row25_2));
 sky130_fd_sc_hd__dfxtp_1 _1249_ (.CLK(clknet_leaf_111_clk),
    .D(booth_b52_m51),
    .Q(pp_row103_7));
 sky130_fd_sc_hd__dfxtp_1 _1250_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b6_m19),
    .Q(pp_row25_3));
 sky130_fd_sc_hd__dfxtp_1 _1251_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b8_m17),
    .Q(pp_row25_4));
 sky130_fd_sc_hd__dfxtp_1 _1252_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b10_m15),
    .Q(pp_row25_5));
 sky130_fd_sc_hd__dfxtp_1 _1253_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b12_m13),
    .Q(pp_row25_6));
 sky130_fd_sc_hd__dfxtp_1 _1254_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b14_m11),
    .Q(pp_row25_7));
 sky130_fd_sc_hd__dfxtp_1 _1255_ (.CLK(clknet_leaf_11_clk),
    .D(booth_b16_m9),
    .Q(pp_row25_8));
 sky130_fd_sc_hd__dfxtp_1 _1256_ (.CLK(clknet_leaf_11_clk),
    .D(booth_b18_m7),
    .Q(pp_row25_9));
 sky130_fd_sc_hd__dfxtp_1 _1257_ (.CLK(clknet_leaf_11_clk),
    .D(booth_b20_m5),
    .Q(pp_row25_10));
 sky130_fd_sc_hd__dfxtp_1 _1258_ (.CLK(clknet_leaf_9_clk),
    .D(booth_b22_m3),
    .Q(pp_row25_11));
 sky130_fd_sc_hd__dfxtp_1 _1259_ (.CLK(clknet_leaf_9_clk),
    .D(booth_b24_m1),
    .Q(pp_row25_12));
 sky130_fd_sc_hd__dfxtp_1 _1260_ (.CLK(clknet_leaf_109_clk),
    .D(booth_b54_m49),
    .Q(pp_row103_8));
 sky130_fd_sc_hd__dfxtp_1 _1261_ (.CLK(clknet_leaf_248_clk),
    .D(net174),
    .Q(pp_row25_13));
 sky130_fd_sc_hd__dfxtp_1 _1262_ (.CLK(clknet_leaf_2_clk),
    .D(booth_b0_m26),
    .Q(pp_row26_0));
 sky130_fd_sc_hd__dfxtp_1 _1263_ (.CLK(clknet_leaf_2_clk),
    .D(booth_b2_m24),
    .Q(pp_row26_1));
 sky130_fd_sc_hd__dfxtp_1 _1264_ (.CLK(clknet_leaf_2_clk),
    .D(booth_b4_m22),
    .Q(pp_row26_2));
 sky130_fd_sc_hd__dfxtp_1 _1265_ (.CLK(clknet_leaf_2_clk),
    .D(booth_b6_m20),
    .Q(pp_row26_3));
 sky130_fd_sc_hd__dfxtp_1 _1266_ (.CLK(clknet_leaf_2_clk),
    .D(booth_b8_m18),
    .Q(pp_row26_4));
 sky130_fd_sc_hd__dfxtp_1 _1267_ (.CLK(clknet_leaf_2_clk),
    .D(booth_b10_m16),
    .Q(pp_row26_5));
 sky130_fd_sc_hd__dfxtp_1 _1268_ (.CLK(clknet_leaf_1_clk),
    .D(booth_b12_m14),
    .Q(pp_row26_6));
 sky130_fd_sc_hd__dfxtp_1 _1269_ (.CLK(clknet_leaf_1_clk),
    .D(booth_b14_m12),
    .Q(pp_row26_7));
 sky130_fd_sc_hd__dfxtp_1 _1270_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b16_m10),
    .Q(pp_row26_8));
 sky130_fd_sc_hd__dfxtp_1 _1271_ (.CLK(clknet_leaf_120_clk),
    .D(booth_b56_m47),
    .Q(pp_row103_9));
 sky130_fd_sc_hd__dfxtp_1 _1272_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b18_m8),
    .Q(pp_row26_9));
 sky130_fd_sc_hd__dfxtp_1 _1273_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b20_m6),
    .Q(pp_row26_10));
 sky130_fd_sc_hd__dfxtp_1 _1274_ (.CLK(clknet_leaf_11_clk),
    .D(booth_b22_m4),
    .Q(pp_row26_11));
 sky130_fd_sc_hd__dfxtp_1 _1275_ (.CLK(clknet_leaf_11_clk),
    .D(booth_b24_m2),
    .Q(pp_row26_12));
 sky130_fd_sc_hd__dfxtp_1 _1276_ (.CLK(clknet_leaf_8_clk),
    .D(booth_b26_m0),
    .Q(pp_row26_13));
 sky130_fd_sc_hd__dfxtp_1 _1277_ (.CLK(clknet_leaf_9_clk),
    .D(net1458),
    .Q(pp_row26_14));
 sky130_fd_sc_hd__dfxtp_2 _1278_ (.CLK(clknet_leaf_244_clk),
    .D(net175),
    .Q(pp_row26_15));
 sky130_fd_sc_hd__dfxtp_1 _1279_ (.CLK(clknet_leaf_251_clk),
    .D(booth_b0_m27),
    .Q(pp_row27_0));
 sky130_fd_sc_hd__dfxtp_1 _1280_ (.CLK(clknet_leaf_250_clk),
    .D(booth_b2_m25),
    .Q(pp_row27_1));
 sky130_fd_sc_hd__dfxtp_1 _1281_ (.CLK(clknet_leaf_250_clk),
    .D(booth_b4_m23),
    .Q(pp_row27_2));
 sky130_fd_sc_hd__dfxtp_1 _1282_ (.CLK(clknet_leaf_120_clk),
    .D(booth_b58_m45),
    .Q(pp_row103_10));
 sky130_fd_sc_hd__dfxtp_2 _1283_ (.CLK(clknet_leaf_181_clk),
    .D(net154),
    .Q(pp_row122_5));
 sky130_fd_sc_hd__dfxtp_1 _1284_ (.CLK(clknet_leaf_1_clk),
    .D(booth_b6_m21),
    .Q(pp_row27_3));
 sky130_fd_sc_hd__dfxtp_1 _1285_ (.CLK(clknet_leaf_1_clk),
    .D(booth_b8_m19),
    .Q(pp_row27_4));
 sky130_fd_sc_hd__dfxtp_1 _1286_ (.CLK(clknet_leaf_1_clk),
    .D(booth_b10_m17),
    .Q(pp_row27_5));
 sky130_fd_sc_hd__dfxtp_1 _1287_ (.CLK(clknet_leaf_1_clk),
    .D(booth_b12_m15),
    .Q(pp_row27_6));
 sky130_fd_sc_hd__dfxtp_1 _1288_ (.CLK(clknet_leaf_1_clk),
    .D(booth_b14_m13),
    .Q(pp_row27_7));
 sky130_fd_sc_hd__dfxtp_1 _1289_ (.CLK(clknet_leaf_2_clk),
    .D(booth_b16_m11),
    .Q(pp_row27_8));
 sky130_fd_sc_hd__dfxtp_1 _1290_ (.CLK(clknet_leaf_2_clk),
    .D(booth_b18_m9),
    .Q(pp_row27_9));
 sky130_fd_sc_hd__dfxtp_1 _1291_ (.CLK(clknet_leaf_2_clk),
    .D(booth_b20_m7),
    .Q(pp_row27_10));
 sky130_fd_sc_hd__dfxtp_1 _1292_ (.CLK(clknet_leaf_3_clk),
    .D(booth_b22_m5),
    .Q(pp_row27_11));
 sky130_fd_sc_hd__dfxtp_1 _1293_ (.CLK(clknet_leaf_3_clk),
    .D(booth_b24_m3),
    .Q(pp_row27_12));
 sky130_fd_sc_hd__dfxtp_1 _1294_ (.CLK(clknet_leaf_119_clk),
    .D(booth_b60_m43),
    .Q(pp_row103_11));
 sky130_fd_sc_hd__dfxtp_1 _1295_ (.CLK(clknet_leaf_3_clk),
    .D(booth_b26_m1),
    .Q(pp_row27_13));
 sky130_fd_sc_hd__dfxtp_1 _1296_ (.CLK(clknet_leaf_248_clk),
    .D(net176),
    .Q(pp_row27_14));
 sky130_fd_sc_hd__dfxtp_1 _1297_ (.CLK(clknet_leaf_251_clk),
    .D(booth_b0_m28),
    .Q(pp_row28_0));
 sky130_fd_sc_hd__dfxtp_1 _1298_ (.CLK(clknet_leaf_251_clk),
    .D(booth_b2_m26),
    .Q(pp_row28_1));
 sky130_fd_sc_hd__dfxtp_1 _1299_ (.CLK(clknet_leaf_250_clk),
    .D(booth_b4_m24),
    .Q(pp_row28_2));
 sky130_fd_sc_hd__dfxtp_1 _1300_ (.CLK(clknet_leaf_250_clk),
    .D(booth_b6_m22),
    .Q(pp_row28_3));
 sky130_fd_sc_hd__dfxtp_1 _1301_ (.CLK(clknet_leaf_250_clk),
    .D(booth_b8_m20),
    .Q(pp_row28_4));
 sky130_fd_sc_hd__dfxtp_1 _1302_ (.CLK(clknet_leaf_250_clk),
    .D(booth_b10_m18),
    .Q(pp_row28_5));
 sky130_fd_sc_hd__dfxtp_1 _1303_ (.CLK(clknet_leaf_1_clk),
    .D(booth_b12_m16),
    .Q(pp_row28_6));
 sky130_fd_sc_hd__dfxtp_1 _1304_ (.CLK(clknet_leaf_1_clk),
    .D(booth_b14_m14),
    .Q(pp_row28_7));
 sky130_fd_sc_hd__dfxtp_1 _1305_ (.CLK(clknet_leaf_122_clk),
    .D(booth_b62_m41),
    .Q(pp_row103_12));
 sky130_fd_sc_hd__dfxtp_1 _1306_ (.CLK(clknet_leaf_1_clk),
    .D(booth_b16_m12),
    .Q(pp_row28_8));
 sky130_fd_sc_hd__dfxtp_1 _1307_ (.CLK(clknet_leaf_1_clk),
    .D(booth_b18_m10),
    .Q(pp_row28_9));
 sky130_fd_sc_hd__dfxtp_1 _1308_ (.CLK(clknet_leaf_1_clk),
    .D(booth_b20_m8),
    .Q(pp_row28_10));
 sky130_fd_sc_hd__dfxtp_1 _1309_ (.CLK(clknet_leaf_3_clk),
    .D(booth_b22_m6),
    .Q(pp_row28_11));
 sky130_fd_sc_hd__dfxtp_1 _1310_ (.CLK(clknet_leaf_2_clk),
    .D(booth_b24_m4),
    .Q(pp_row28_12));
 sky130_fd_sc_hd__dfxtp_1 _1311_ (.CLK(clknet_leaf_3_clk),
    .D(booth_b26_m2),
    .Q(pp_row28_13));
 sky130_fd_sc_hd__dfxtp_1 _1312_ (.CLK(clknet_leaf_246_clk),
    .D(booth_b28_m0),
    .Q(pp_row28_14));
 sky130_fd_sc_hd__dfxtp_1 _1313_ (.CLK(clknet_leaf_246_clk),
    .D(net1448),
    .Q(pp_row28_15));
 sky130_fd_sc_hd__dfxtp_1 _1314_ (.CLK(clknet_leaf_244_clk),
    .D(net177),
    .Q(pp_row28_16));
 sky130_fd_sc_hd__dfxtp_1 _1315_ (.CLK(clknet_leaf_246_clk),
    .D(booth_b0_m29),
    .Q(pp_row29_0));
 sky130_fd_sc_hd__dfxtp_1 _1316_ (.CLK(clknet_leaf_122_clk),
    .D(booth_b64_m39),
    .Q(pp_row103_13));
 sky130_fd_sc_hd__dfxtp_1 _1317_ (.CLK(clknet_leaf_247_clk),
    .D(booth_b2_m27),
    .Q(pp_row29_1));
 sky130_fd_sc_hd__dfxtp_1 _1318_ (.CLK(clknet_leaf_247_clk),
    .D(booth_b4_m25),
    .Q(pp_row29_2));
 sky130_fd_sc_hd__dfxtp_1 _1319_ (.CLK(clknet_leaf_250_clk),
    .D(booth_b6_m23),
    .Q(pp_row29_3));
 sky130_fd_sc_hd__dfxtp_1 _1320_ (.CLK(clknet_leaf_250_clk),
    .D(booth_b8_m21),
    .Q(pp_row29_4));
 sky130_fd_sc_hd__dfxtp_1 _1321_ (.CLK(clknet_leaf_0_clk),
    .D(booth_b10_m19),
    .Q(pp_row29_5));
 sky130_fd_sc_hd__dfxtp_1 _1322_ (.CLK(clknet_leaf_0_clk),
    .D(booth_b12_m17),
    .Q(pp_row29_6));
 sky130_fd_sc_hd__dfxtp_1 _1323_ (.CLK(clknet_leaf_1_clk),
    .D(booth_b14_m15),
    .Q(pp_row29_7));
 sky130_fd_sc_hd__dfxtp_1 _1324_ (.CLK(clknet_leaf_250_clk),
    .D(booth_b16_m13),
    .Q(pp_row29_8));
 sky130_fd_sc_hd__dfxtp_1 _1325_ (.CLK(clknet_leaf_1_clk),
    .D(booth_b18_m11),
    .Q(pp_row29_9));
 sky130_fd_sc_hd__dfxtp_1 _1326_ (.CLK(clknet_leaf_1_clk),
    .D(booth_b20_m9),
    .Q(pp_row29_10));
 sky130_fd_sc_hd__dfxtp_2 _1327_ (.CLK(clknet_leaf_184_clk),
    .D(net133),
    .Q(pp_row103_14));
 sky130_fd_sc_hd__dfxtp_1 _1328_ (.CLK(clknet_leaf_4_clk),
    .D(booth_b22_m7),
    .Q(pp_row29_11));
 sky130_fd_sc_hd__dfxtp_1 _1329_ (.CLK(clknet_leaf_4_clk),
    .D(booth_b24_m5),
    .Q(pp_row29_12));
 sky130_fd_sc_hd__dfxtp_1 _1330_ (.CLK(clknet_leaf_4_clk),
    .D(booth_b26_m3),
    .Q(pp_row29_13));
 sky130_fd_sc_hd__dfxtp_1 _1331_ (.CLK(clknet_leaf_246_clk),
    .D(booth_b28_m1),
    .Q(pp_row29_14));
 sky130_fd_sc_hd__dfxtp_1 _1332_ (.CLK(clknet_leaf_244_clk),
    .D(net178),
    .Q(pp_row29_15));
 sky130_fd_sc_hd__dfxtp_1 _1333_ (.CLK(clknet_leaf_0_clk),
    .D(booth_b0_m30),
    .Q(pp_row30_0));
 sky130_fd_sc_hd__dfxtp_1 _1334_ (.CLK(clknet_leaf_0_clk),
    .D(booth_b2_m28),
    .Q(pp_row30_1));
 sky130_fd_sc_hd__dfxtp_1 _1335_ (.CLK(clknet_leaf_0_clk),
    .D(booth_b4_m26),
    .Q(pp_row30_2));
 sky130_fd_sc_hd__dfxtp_1 _1336_ (.CLK(clknet_leaf_247_clk),
    .D(booth_b6_m24),
    .Q(pp_row30_3));
 sky130_fd_sc_hd__dfxtp_1 _1337_ (.CLK(clknet_leaf_0_clk),
    .D(booth_b8_m22),
    .Q(pp_row30_4));
 sky130_fd_sc_hd__dfxtp_1 _1338_ (.CLK(clknet_leaf_123_clk),
    .D(booth_b40_m64),
    .Q(pp_row104_1));
 sky130_fd_sc_hd__dfxtp_1 _1339_ (.CLK(clknet_leaf_0_clk),
    .D(booth_b10_m20),
    .Q(pp_row30_5));
 sky130_fd_sc_hd__dfxtp_1 _1340_ (.CLK(clknet_leaf_0_clk),
    .D(booth_b12_m18),
    .Q(pp_row30_6));
 sky130_fd_sc_hd__dfxtp_1 _1341_ (.CLK(clknet_leaf_0_clk),
    .D(booth_b14_m16),
    .Q(pp_row30_7));
 sky130_fd_sc_hd__dfxtp_1 _1342_ (.CLK(clknet_leaf_0_clk),
    .D(booth_b16_m14),
    .Q(pp_row30_8));
 sky130_fd_sc_hd__dfxtp_1 _1343_ (.CLK(clknet_leaf_3_clk),
    .D(booth_b18_m12),
    .Q(pp_row30_9));
 sky130_fd_sc_hd__dfxtp_1 _1344_ (.CLK(clknet_leaf_3_clk),
    .D(booth_b20_m10),
    .Q(pp_row30_10));
 sky130_fd_sc_hd__dfxtp_1 _1345_ (.CLK(clknet_leaf_3_clk),
    .D(booth_b22_m8),
    .Q(pp_row30_11));
 sky130_fd_sc_hd__dfxtp_1 _1346_ (.CLK(clknet_leaf_3_clk),
    .D(booth_b24_m6),
    .Q(pp_row30_12));
 sky130_fd_sc_hd__dfxtp_1 _1347_ (.CLK(clknet_leaf_3_clk),
    .D(booth_b26_m4),
    .Q(pp_row30_13));
 sky130_fd_sc_hd__dfxtp_1 _1348_ (.CLK(clknet_leaf_241_clk),
    .D(booth_b28_m2),
    .Q(pp_row30_14));
 sky130_fd_sc_hd__dfxtp_1 _1349_ (.CLK(clknet_leaf_123_clk),
    .D(booth_b42_m62),
    .Q(pp_row104_2));
 sky130_fd_sc_hd__dfxtp_1 _1350_ (.CLK(clknet_leaf_246_clk),
    .D(booth_b30_m0),
    .Q(pp_row30_15));
 sky130_fd_sc_hd__dfxtp_1 _1351_ (.CLK(clknet_leaf_241_clk),
    .D(net1439),
    .Q(pp_row30_16));
 sky130_fd_sc_hd__dfxtp_1 _1352_ (.CLK(clknet_leaf_244_clk),
    .D(net180),
    .Q(pp_row30_17));
 sky130_fd_sc_hd__dfxtp_1 _1353_ (.CLK(clknet_leaf_4_clk),
    .D(booth_b0_m31),
    .Q(pp_row31_0));
 sky130_fd_sc_hd__dfxtp_1 _1354_ (.CLK(clknet_leaf_4_clk),
    .D(booth_b2_m29),
    .Q(pp_row31_1));
 sky130_fd_sc_hd__dfxtp_1 _1355_ (.CLK(clknet_leaf_3_clk),
    .D(booth_b4_m27),
    .Q(pp_row31_2));
 sky130_fd_sc_hd__dfxtp_1 _1356_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b6_m25),
    .Q(pp_row31_3));
 sky130_fd_sc_hd__dfxtp_1 _1357_ (.CLK(clknet_leaf_2_clk),
    .D(booth_b8_m23),
    .Q(pp_row31_4));
 sky130_fd_sc_hd__dfxtp_1 _1358_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b10_m21),
    .Q(pp_row31_5));
 sky130_fd_sc_hd__dfxtp_1 _1359_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b12_m19),
    .Q(pp_row31_6));
 sky130_fd_sc_hd__dfxtp_1 _1360_ (.CLK(clknet_leaf_110_clk),
    .D(booth_b44_m60),
    .Q(pp_row104_3));
 sky130_fd_sc_hd__dfxtp_1 _1361_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b14_m17),
    .Q(pp_row31_7));
 sky130_fd_sc_hd__dfxtp_1 _1362_ (.CLK(clknet_leaf_10_clk),
    .D(booth_b16_m15),
    .Q(pp_row31_8));
 sky130_fd_sc_hd__dfxtp_1 _1363_ (.CLK(clknet_leaf_9_clk),
    .D(booth_b18_m13),
    .Q(pp_row31_9));
 sky130_fd_sc_hd__dfxtp_1 _1364_ (.CLK(clknet_leaf_9_clk),
    .D(booth_b20_m11),
    .Q(pp_row31_10));
 sky130_fd_sc_hd__dfxtp_1 _1365_ (.CLK(clknet_leaf_9_clk),
    .D(booth_b22_m9),
    .Q(pp_row31_11));
 sky130_fd_sc_hd__dfxtp_1 _1366_ (.CLK(clknet_leaf_3_clk),
    .D(booth_b24_m7),
    .Q(pp_row31_12));
 sky130_fd_sc_hd__dfxtp_1 _1367_ (.CLK(clknet_leaf_3_clk),
    .D(booth_b26_m5),
    .Q(pp_row31_13));
 sky130_fd_sc_hd__dfxtp_1 _1368_ (.CLK(clknet_leaf_4_clk),
    .D(booth_b28_m3),
    .Q(pp_row31_14));
 sky130_fd_sc_hd__dfxtp_1 _1369_ (.CLK(clknet_leaf_4_clk),
    .D(booth_b30_m1),
    .Q(pp_row31_15));
 sky130_fd_sc_hd__dfxtp_1 _1370_ (.CLK(clknet_leaf_244_clk),
    .D(net181),
    .Q(pp_row31_16));
 sky130_fd_sc_hd__dfxtp_1 _1371_ (.CLK(clknet_leaf_110_clk),
    .D(booth_b46_m58),
    .Q(pp_row104_4));
 sky130_fd_sc_hd__dfxtp_1 _1372_ (.CLK(clknet_leaf_7_clk),
    .D(booth_b0_m32),
    .Q(pp_row32_0));
 sky130_fd_sc_hd__dfxtp_1 _1373_ (.CLK(clknet_leaf_7_clk),
    .D(booth_b2_m30),
    .Q(pp_row32_1));
 sky130_fd_sc_hd__dfxtp_1 _1374_ (.CLK(clknet_leaf_9_clk),
    .D(booth_b4_m28),
    .Q(pp_row32_2));
 sky130_fd_sc_hd__dfxtp_1 _1375_ (.CLK(clknet_leaf_7_clk),
    .D(booth_b6_m26),
    .Q(pp_row32_3));
 sky130_fd_sc_hd__dfxtp_1 _1376_ (.CLK(clknet_leaf_7_clk),
    .D(booth_b8_m24),
    .Q(pp_row32_4));
 sky130_fd_sc_hd__dfxtp_1 _1377_ (.CLK(clknet_leaf_7_clk),
    .D(booth_b10_m22),
    .Q(pp_row32_5));
 sky130_fd_sc_hd__dfxtp_1 _1378_ (.CLK(clknet_leaf_43_clk),
    .D(booth_b12_m20),
    .Q(pp_row32_6));
 sky130_fd_sc_hd__dfxtp_1 _1379_ (.CLK(clknet_leaf_35_clk),
    .D(booth_b14_m18),
    .Q(pp_row32_7));
 sky130_fd_sc_hd__dfxtp_1 _1380_ (.CLK(clknet_leaf_42_clk),
    .D(booth_b16_m16),
    .Q(pp_row32_8));
 sky130_fd_sc_hd__dfxtp_1 _1381_ (.CLK(clknet_leaf_43_clk),
    .D(booth_b18_m14),
    .Q(pp_row32_9));
 sky130_fd_sc_hd__dfxtp_1 _1382_ (.CLK(clknet_leaf_110_clk),
    .D(booth_b48_m56),
    .Q(pp_row104_5));
 sky130_fd_sc_hd__dfxtp_1 _1383_ (.CLK(clknet_leaf_44_clk),
    .D(booth_b20_m12),
    .Q(pp_row32_10));
 sky130_fd_sc_hd__dfxtp_1 _1384_ (.CLK(clknet_leaf_44_clk),
    .D(booth_b22_m10),
    .Q(pp_row32_11));
 sky130_fd_sc_hd__dfxtp_1 _1385_ (.CLK(clknet_leaf_42_clk),
    .D(booth_b24_m8),
    .Q(pp_row32_12));
 sky130_fd_sc_hd__dfxtp_1 _1386_ (.CLK(clknet_leaf_42_clk),
    .D(booth_b26_m6),
    .Q(pp_row32_13));
 sky130_fd_sc_hd__dfxtp_1 _1387_ (.CLK(clknet_leaf_42_clk),
    .D(booth_b28_m4),
    .Q(pp_row32_14));
 sky130_fd_sc_hd__dfxtp_1 _1388_ (.CLK(clknet_leaf_45_clk),
    .D(booth_b30_m2),
    .Q(pp_row32_15));
 sky130_fd_sc_hd__dfxtp_1 _1389_ (.CLK(clknet_leaf_45_clk),
    .D(booth_b32_m0),
    .Q(pp_row32_16));
 sky130_fd_sc_hd__dfxtp_1 _1390_ (.CLK(clknet_leaf_5_clk),
    .D(net1430),
    .Q(pp_row32_17));
 sky130_fd_sc_hd__dfxtp_1 _1391_ (.CLK(clknet_leaf_244_clk),
    .D(net182),
    .Q(pp_row32_18));
 sky130_fd_sc_hd__dfxtp_1 _1392_ (.CLK(clknet_leaf_54_clk),
    .D(booth_b0_m33),
    .Q(pp_row33_0));
 sky130_fd_sc_hd__dfxtp_1 _1393_ (.CLK(clknet_leaf_110_clk),
    .D(booth_b50_m54),
    .Q(pp_row104_6));
 sky130_fd_sc_hd__dfxtp_1 _1394_ (.CLK(clknet_leaf_164_clk),
    .D(\notsign$6504 ),
    .Q(pp_row123_0));
 sky130_fd_sc_hd__dfxtp_1 _1395_ (.CLK(clknet_leaf_181_clk),
    .D(net159),
    .Q(pp_row127_2));
 sky130_fd_sc_hd__dfxtp_1 _1396_ (.CLK(clknet_leaf_54_clk),
    .D(booth_b2_m31),
    .Q(pp_row33_1));
 sky130_fd_sc_hd__dfxtp_1 _1397_ (.CLK(clknet_leaf_54_clk),
    .D(booth_b4_m29),
    .Q(pp_row33_2));
 sky130_fd_sc_hd__dfxtp_1 _1398_ (.CLK(clknet_leaf_54_clk),
    .D(booth_b6_m27),
    .Q(pp_row33_3));
 sky130_fd_sc_hd__dfxtp_1 _1399_ (.CLK(clknet_leaf_54_clk),
    .D(booth_b8_m25),
    .Q(pp_row33_4));
 sky130_fd_sc_hd__dfxtp_1 _1400_ (.CLK(clknet_leaf_53_clk),
    .D(booth_b10_m23),
    .Q(pp_row33_5));
 sky130_fd_sc_hd__dfxtp_1 _1401_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b12_m21),
    .Q(pp_row33_6));
 sky130_fd_sc_hd__dfxtp_1 _1402_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b14_m19),
    .Q(pp_row33_7));
 sky130_fd_sc_hd__dfxtp_1 _1403_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b16_m17),
    .Q(pp_row33_8));
 sky130_fd_sc_hd__dfxtp_1 _1404_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b18_m15),
    .Q(pp_row33_9));
 sky130_fd_sc_hd__dfxtp_1 _1405_ (.CLK(clknet_leaf_51_clk),
    .D(booth_b20_m13),
    .Q(pp_row33_10));
 sky130_fd_sc_hd__dfxtp_1 _1406_ (.CLK(clknet_leaf_109_clk),
    .D(booth_b52_m52),
    .Q(pp_row104_7));
 sky130_fd_sc_hd__dfxtp_1 _1407_ (.CLK(clknet_leaf_54_clk),
    .D(booth_b22_m11),
    .Q(pp_row33_11));
 sky130_fd_sc_hd__dfxtp_1 _1408_ (.CLK(clknet_leaf_57_clk),
    .D(booth_b24_m9),
    .Q(pp_row33_12));
 sky130_fd_sc_hd__dfxtp_1 _1409_ (.CLK(clknet_leaf_57_clk),
    .D(booth_b26_m7),
    .Q(pp_row33_13));
 sky130_fd_sc_hd__dfxtp_1 _1410_ (.CLK(clknet_leaf_58_clk),
    .D(booth_b28_m5),
    .Q(pp_row33_14));
 sky130_fd_sc_hd__dfxtp_1 _1411_ (.CLK(clknet_leaf_41_clk),
    .D(booth_b30_m3),
    .Q(pp_row33_15));
 sky130_fd_sc_hd__dfxtp_1 _1412_ (.CLK(clknet_leaf_41_clk),
    .D(booth_b32_m1),
    .Q(pp_row33_16));
 sky130_fd_sc_hd__dfxtp_1 _1413_ (.CLK(clknet_leaf_244_clk),
    .D(net183),
    .Q(pp_row33_17));
 sky130_fd_sc_hd__dfxtp_1 _1414_ (.CLK(clknet_leaf_40_clk),
    .D(booth_b0_m34),
    .Q(pp_row34_0));
 sky130_fd_sc_hd__dfxtp_1 _1415_ (.CLK(clknet_leaf_40_clk),
    .D(booth_b2_m32),
    .Q(pp_row34_1));
 sky130_fd_sc_hd__dfxtp_1 _1416_ (.CLK(clknet_leaf_56_clk),
    .D(booth_b4_m30),
    .Q(pp_row34_2));
 sky130_fd_sc_hd__dfxtp_1 _1417_ (.CLK(clknet_leaf_121_clk),
    .D(booth_b54_m50),
    .Q(pp_row104_8));
 sky130_fd_sc_hd__dfxtp_1 _1418_ (.CLK(clknet_leaf_56_clk),
    .D(booth_b6_m28),
    .Q(pp_row34_3));
 sky130_fd_sc_hd__dfxtp_1 _1419_ (.CLK(clknet_leaf_56_clk),
    .D(booth_b8_m26),
    .Q(pp_row34_4));
 sky130_fd_sc_hd__dfxtp_1 _1420_ (.CLK(clknet_leaf_54_clk),
    .D(booth_b10_m24),
    .Q(pp_row34_5));
 sky130_fd_sc_hd__dfxtp_1 _1421_ (.CLK(clknet_leaf_54_clk),
    .D(booth_b12_m22),
    .Q(pp_row34_6));
 sky130_fd_sc_hd__dfxtp_1 _1422_ (.CLK(clknet_leaf_55_clk),
    .D(booth_b14_m20),
    .Q(pp_row34_7));
 sky130_fd_sc_hd__dfxtp_1 _1423_ (.CLK(clknet_leaf_56_clk),
    .D(booth_b16_m18),
    .Q(pp_row34_8));
 sky130_fd_sc_hd__dfxtp_1 _1424_ (.CLK(clknet_leaf_56_clk),
    .D(booth_b18_m16),
    .Q(pp_row34_9));
 sky130_fd_sc_hd__dfxtp_1 _1425_ (.CLK(clknet_leaf_56_clk),
    .D(booth_b20_m14),
    .Q(pp_row34_10));
 sky130_fd_sc_hd__dfxtp_1 _1426_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b22_m12),
    .Q(pp_row34_11));
 sky130_fd_sc_hd__dfxtp_1 _1427_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b24_m10),
    .Q(pp_row34_12));
 sky130_fd_sc_hd__dfxtp_1 _1428_ (.CLK(clknet_leaf_121_clk),
    .D(booth_b56_m48),
    .Q(pp_row104_9));
 sky130_fd_sc_hd__dfxtp_1 _1429_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b26_m8),
    .Q(pp_row34_13));
 sky130_fd_sc_hd__dfxtp_1 _1430_ (.CLK(clknet_leaf_63_clk),
    .D(booth_b28_m6),
    .Q(pp_row34_14));
 sky130_fd_sc_hd__dfxtp_1 _1431_ (.CLK(clknet_leaf_63_clk),
    .D(booth_b30_m4),
    .Q(pp_row34_15));
 sky130_fd_sc_hd__dfxtp_1 _1432_ (.CLK(clknet_leaf_63_clk),
    .D(booth_b32_m2),
    .Q(pp_row34_16));
 sky130_fd_sc_hd__dfxtp_1 _1433_ (.CLK(clknet_leaf_40_clk),
    .D(booth_b34_m0),
    .Q(pp_row34_17));
 sky130_fd_sc_hd__dfxtp_1 _1434_ (.CLK(clknet_leaf_40_clk),
    .D(net1423),
    .Q(pp_row34_18));
 sky130_fd_sc_hd__dfxtp_2 _1435_ (.CLK(clknet_leaf_244_clk),
    .D(net184),
    .Q(pp_row34_19));
 sky130_fd_sc_hd__dfxtp_1 _1436_ (.CLK(clknet_leaf_41_clk),
    .D(booth_b0_m35),
    .Q(pp_row35_0));
 sky130_fd_sc_hd__dfxtp_1 _1437_ (.CLK(clknet_leaf_53_clk),
    .D(booth_b2_m33),
    .Q(pp_row35_1));
 sky130_fd_sc_hd__dfxtp_1 _1438_ (.CLK(clknet_leaf_55_clk),
    .D(booth_b4_m31),
    .Q(pp_row35_2));
 sky130_fd_sc_hd__dfxtp_1 _1439_ (.CLK(clknet_leaf_121_clk),
    .D(booth_b58_m46),
    .Q(pp_row104_10));
 sky130_fd_sc_hd__dfxtp_1 _1440_ (.CLK(clknet_leaf_54_clk),
    .D(booth_b6_m29),
    .Q(pp_row35_3));
 sky130_fd_sc_hd__dfxtp_1 _1441_ (.CLK(clknet_leaf_54_clk),
    .D(booth_b8_m27),
    .Q(pp_row35_4));
 sky130_fd_sc_hd__dfxtp_1 _1442_ (.CLK(clknet_leaf_54_clk),
    .D(booth_b10_m25),
    .Q(pp_row35_5));
 sky130_fd_sc_hd__dfxtp_1 _1443_ (.CLK(clknet_leaf_55_clk),
    .D(booth_b12_m23),
    .Q(pp_row35_6));
 sky130_fd_sc_hd__dfxtp_1 _1444_ (.CLK(clknet_leaf_54_clk),
    .D(booth_b14_m21),
    .Q(pp_row35_7));
 sky130_fd_sc_hd__dfxtp_1 _1445_ (.CLK(clknet_leaf_65_clk),
    .D(booth_b16_m19),
    .Q(pp_row35_8));
 sky130_fd_sc_hd__dfxtp_1 _1446_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b18_m17),
    .Q(pp_row35_9));
 sky130_fd_sc_hd__dfxtp_1 _1447_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b20_m15),
    .Q(pp_row35_10));
 sky130_fd_sc_hd__dfxtp_1 _1448_ (.CLK(clknet_leaf_56_clk),
    .D(booth_b22_m13),
    .Q(pp_row35_11));
 sky130_fd_sc_hd__dfxtp_1 _1449_ (.CLK(clknet_leaf_65_clk),
    .D(booth_b24_m11),
    .Q(pp_row35_12));
 sky130_fd_sc_hd__dfxtp_1 _1450_ (.CLK(clknet_leaf_110_clk),
    .D(booth_b60_m44),
    .Q(pp_row104_11));
 sky130_fd_sc_hd__dfxtp_1 _1451_ (.CLK(clknet_leaf_65_clk),
    .D(booth_b26_m9),
    .Q(pp_row35_13));
 sky130_fd_sc_hd__dfxtp_1 _1452_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b28_m7),
    .Q(pp_row35_14));
 sky130_fd_sc_hd__dfxtp_1 _1453_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b30_m5),
    .Q(pp_row35_15));
 sky130_fd_sc_hd__dfxtp_1 _1454_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b32_m3),
    .Q(pp_row35_16));
 sky130_fd_sc_hd__dfxtp_1 _1455_ (.CLK(clknet_leaf_40_clk),
    .D(booth_b34_m1),
    .Q(pp_row35_17));
 sky130_fd_sc_hd__dfxtp_2 _1456_ (.CLK(clknet_leaf_244_clk),
    .D(net185),
    .Q(pp_row35_18));
 sky130_fd_sc_hd__dfxtp_1 _1457_ (.CLK(clknet_leaf_41_clk),
    .D(booth_b0_m36),
    .Q(pp_row36_0));
 sky130_fd_sc_hd__dfxtp_1 _1458_ (.CLK(clknet_leaf_42_clk),
    .D(booth_b2_m34),
    .Q(pp_row36_1));
 sky130_fd_sc_hd__dfxtp_1 _1459_ (.CLK(clknet_leaf_40_clk),
    .D(booth_b4_m32),
    .Q(pp_row36_2));
 sky130_fd_sc_hd__dfxtp_1 _1460_ (.CLK(clknet_leaf_40_clk),
    .D(booth_b6_m30),
    .Q(pp_row36_3));
 sky130_fd_sc_hd__dfxtp_1 _1461_ (.CLK(clknet_leaf_110_clk),
    .D(booth_b62_m42),
    .Q(pp_row104_12));
 sky130_fd_sc_hd__dfxtp_1 _1462_ (.CLK(clknet_leaf_41_clk),
    .D(booth_b8_m28),
    .Q(pp_row36_4));
 sky130_fd_sc_hd__dfxtp_1 _1463_ (.CLK(clknet_leaf_40_clk),
    .D(booth_b10_m26),
    .Q(pp_row36_5));
 sky130_fd_sc_hd__dfxtp_1 _1464_ (.CLK(clknet_leaf_40_clk),
    .D(booth_b12_m24),
    .Q(pp_row36_6));
 sky130_fd_sc_hd__dfxtp_1 _1465_ (.CLK(clknet_leaf_39_clk),
    .D(booth_b14_m22),
    .Q(pp_row36_7));
 sky130_fd_sc_hd__dfxtp_1 _1466_ (.CLK(clknet_leaf_40_clk),
    .D(booth_b16_m20),
    .Q(pp_row36_8));
 sky130_fd_sc_hd__dfxtp_1 _1467_ (.CLK(clknet_leaf_40_clk),
    .D(booth_b18_m18),
    .Q(pp_row36_9));
 sky130_fd_sc_hd__dfxtp_1 _1468_ (.CLK(clknet_leaf_40_clk),
    .D(booth_b20_m16),
    .Q(pp_row36_10));
 sky130_fd_sc_hd__dfxtp_1 _1469_ (.CLK(clknet_leaf_39_clk),
    .D(booth_b22_m14),
    .Q(pp_row36_11));
 sky130_fd_sc_hd__dfxtp_1 _1470_ (.CLK(clknet_leaf_39_clk),
    .D(booth_b24_m12),
    .Q(pp_row36_12));
 sky130_fd_sc_hd__dfxtp_1 _1471_ (.CLK(clknet_leaf_39_clk),
    .D(booth_b26_m10),
    .Q(pp_row36_13));
 sky130_fd_sc_hd__dfxtp_1 _1472_ (.CLK(clknet_leaf_110_clk),
    .D(booth_b64_m40),
    .Q(pp_row104_13));
 sky130_fd_sc_hd__dfxtp_1 _1473_ (.CLK(clknet_leaf_39_clk),
    .D(booth_b28_m8),
    .Q(pp_row36_14));
 sky130_fd_sc_hd__dfxtp_1 _1474_ (.CLK(clknet_leaf_39_clk),
    .D(booth_b30_m6),
    .Q(pp_row36_15));
 sky130_fd_sc_hd__dfxtp_1 _1475_ (.CLK(clknet_leaf_39_clk),
    .D(booth_b32_m4),
    .Q(pp_row36_16));
 sky130_fd_sc_hd__dfxtp_1 _1476_ (.CLK(clknet_leaf_38_clk),
    .D(booth_b34_m2),
    .Q(pp_row36_17));
 sky130_fd_sc_hd__dfxtp_1 _1477_ (.CLK(clknet_leaf_38_clk),
    .D(booth_b36_m0),
    .Q(pp_row36_18));
 sky130_fd_sc_hd__dfxtp_1 _1478_ (.CLK(clknet_leaf_38_clk),
    .D(net1406),
    .Q(pp_row36_19));
 sky130_fd_sc_hd__dfxtp_2 _1479_ (.CLK(clknet_leaf_236_clk),
    .D(net186),
    .Q(pp_row36_20));
 sky130_fd_sc_hd__dfxtp_1 _1480_ (.CLK(clknet_leaf_241_clk),
    .D(booth_b0_m37),
    .Q(pp_row37_0));
 sky130_fd_sc_hd__dfxtp_1 _1481_ (.CLK(clknet_leaf_246_clk),
    .D(booth_b2_m35),
    .Q(pp_row37_1));
 sky130_fd_sc_hd__dfxtp_1 _1482_ (.CLK(clknet_leaf_241_clk),
    .D(booth_b4_m33),
    .Q(pp_row37_2));
 sky130_fd_sc_hd__dfxtp_2 _1483_ (.CLK(clknet_leaf_184_clk),
    .D(net134),
    .Q(pp_row104_14));
 sky130_fd_sc_hd__dfxtp_1 _1484_ (.CLK(clknet_leaf_45_clk),
    .D(booth_b6_m31),
    .Q(pp_row37_3));
 sky130_fd_sc_hd__dfxtp_1 _1485_ (.CLK(clknet_leaf_45_clk),
    .D(booth_b8_m29),
    .Q(pp_row37_4));
 sky130_fd_sc_hd__dfxtp_1 _1486_ (.CLK(clknet_leaf_43_clk),
    .D(booth_b10_m27),
    .Q(pp_row37_5));
 sky130_fd_sc_hd__dfxtp_1 _1487_ (.CLK(clknet_leaf_34_clk),
    .D(booth_b12_m25),
    .Q(pp_row37_6));
 sky130_fd_sc_hd__dfxtp_1 _1488_ (.CLK(clknet_leaf_43_clk),
    .D(booth_b14_m23),
    .Q(pp_row37_7));
 sky130_fd_sc_hd__dfxtp_1 _1489_ (.CLK(clknet_leaf_43_clk),
    .D(booth_b16_m21),
    .Q(pp_row37_8));
 sky130_fd_sc_hd__dfxtp_1 _1490_ (.CLK(clknet_leaf_44_clk),
    .D(booth_b18_m19),
    .Q(pp_row37_9));
 sky130_fd_sc_hd__dfxtp_1 _1491_ (.CLK(clknet_leaf_18_clk),
    .D(booth_b20_m17),
    .Q(pp_row37_10));
 sky130_fd_sc_hd__dfxtp_1 _1492_ (.CLK(clknet_leaf_45_clk),
    .D(booth_b22_m15),
    .Q(pp_row37_11));
 sky130_fd_sc_hd__dfxtp_1 _1493_ (.CLK(clknet_leaf_45_clk),
    .D(booth_b24_m13),
    .Q(pp_row37_12));
 sky130_fd_sc_hd__dfxtp_1 _1494_ (.CLK(clknet_leaf_122_clk),
    .D(\notsign$5874 ),
    .Q(pp_row105_0));
 sky130_fd_sc_hd__dfxtp_1 _1495_ (.CLK(clknet_leaf_45_clk),
    .D(booth_b26_m11),
    .Q(pp_row37_13));
 sky130_fd_sc_hd__dfxtp_1 _1496_ (.CLK(clknet_leaf_45_clk),
    .D(booth_b28_m9),
    .Q(pp_row37_14));
 sky130_fd_sc_hd__dfxtp_1 _1497_ (.CLK(clknet_leaf_45_clk),
    .D(booth_b30_m7),
    .Q(pp_row37_15));
 sky130_fd_sc_hd__dfxtp_1 _1498_ (.CLK(clknet_leaf_45_clk),
    .D(booth_b32_m5),
    .Q(pp_row37_16));
 sky130_fd_sc_hd__dfxtp_1 _1499_ (.CLK(clknet_leaf_41_clk),
    .D(booth_b34_m3),
    .Q(pp_row37_17));
 sky130_fd_sc_hd__dfxtp_1 _1500_ (.CLK(clknet_leaf_45_clk),
    .D(booth_b36_m1),
    .Q(pp_row37_18));
 sky130_fd_sc_hd__dfxtp_2 _1501_ (.CLK(clknet_leaf_244_clk),
    .D(net187),
    .Q(pp_row37_19));
 sky130_fd_sc_hd__dfxtp_1 _1502_ (.CLK(clknet_leaf_20_clk),
    .D(booth_b0_m38),
    .Q(pp_row38_0));
 sky130_fd_sc_hd__dfxtp_1 _1503_ (.CLK(clknet_leaf_17_clk),
    .D(booth_b2_m36),
    .Q(pp_row38_1));
 sky130_fd_sc_hd__dfxtp_1 _1504_ (.CLK(clknet_leaf_20_clk),
    .D(booth_b4_m34),
    .Q(pp_row38_2));
 sky130_fd_sc_hd__dfxtp_1 _1505_ (.CLK(clknet_leaf_122_clk),
    .D(booth_b42_m63),
    .Q(pp_row105_1));
 sky130_fd_sc_hd__dfxtp_1 _1506_ (.CLK(clknet_leaf_164_clk),
    .D(booth_b60_m63),
    .Q(pp_row123_1));
 sky130_fd_sc_hd__dfxtp_1 _1507_ (.CLK(clknet_leaf_16_clk),
    .D(booth_b6_m32),
    .Q(pp_row38_3));
 sky130_fd_sc_hd__dfxtp_1 _1508_ (.CLK(clknet_leaf_16_clk),
    .D(booth_b8_m30),
    .Q(pp_row38_4));
 sky130_fd_sc_hd__dfxtp_1 _1509_ (.CLK(clknet_leaf_17_clk),
    .D(booth_b10_m28),
    .Q(pp_row38_5));
 sky130_fd_sc_hd__dfxtp_1 _1510_ (.CLK(clknet_leaf_44_clk),
    .D(booth_b12_m26),
    .Q(pp_row38_6));
 sky130_fd_sc_hd__dfxtp_1 _1511_ (.CLK(clknet_leaf_44_clk),
    .D(booth_b14_m24),
    .Q(pp_row38_7));
 sky130_fd_sc_hd__dfxtp_1 _1512_ (.CLK(clknet_leaf_44_clk),
    .D(booth_b16_m22),
    .Q(pp_row38_8));
 sky130_fd_sc_hd__dfxtp_1 _1513_ (.CLK(clknet_leaf_44_clk),
    .D(booth_b18_m20),
    .Q(pp_row38_9));
 sky130_fd_sc_hd__dfxtp_1 _1514_ (.CLK(clknet_leaf_17_clk),
    .D(booth_b20_m18),
    .Q(pp_row38_10));
 sky130_fd_sc_hd__dfxtp_1 _1515_ (.CLK(clknet_leaf_17_clk),
    .D(booth_b22_m16),
    .Q(pp_row38_11));
 sky130_fd_sc_hd__dfxtp_1 _1516_ (.CLK(clknet_leaf_17_clk),
    .D(booth_b24_m14),
    .Q(pp_row38_12));
 sky130_fd_sc_hd__dfxtp_1 _1517_ (.CLK(clknet_leaf_121_clk),
    .D(booth_b44_m61),
    .Q(pp_row105_2));
 sky130_fd_sc_hd__dfxtp_1 _1518_ (.CLK(clknet_leaf_17_clk),
    .D(booth_b26_m12),
    .Q(pp_row38_13));
 sky130_fd_sc_hd__dfxtp_1 _1519_ (.CLK(clknet_leaf_246_clk),
    .D(booth_b28_m10),
    .Q(pp_row38_14));
 sky130_fd_sc_hd__dfxtp_1 _1520_ (.CLK(clknet_leaf_246_clk),
    .D(booth_b30_m8),
    .Q(pp_row38_15));
 sky130_fd_sc_hd__dfxtp_1 _1521_ (.CLK(clknet_leaf_246_clk),
    .D(booth_b32_m6),
    .Q(pp_row38_16));
 sky130_fd_sc_hd__dfxtp_1 _1522_ (.CLK(clknet_leaf_242_clk),
    .D(booth_b34_m4),
    .Q(pp_row38_17));
 sky130_fd_sc_hd__dfxtp_1 _1523_ (.CLK(clknet_leaf_242_clk),
    .D(booth_b36_m2),
    .Q(pp_row38_18));
 sky130_fd_sc_hd__dfxtp_1 _1524_ (.CLK(clknet_leaf_242_clk),
    .D(booth_b38_m0),
    .Q(pp_row38_19));
 sky130_fd_sc_hd__dfxtp_1 _1525_ (.CLK(clknet_leaf_241_clk),
    .D(net1394),
    .Q(pp_row38_20));
 sky130_fd_sc_hd__dfxtp_1 _1526_ (.CLK(clknet_leaf_236_clk),
    .D(net188),
    .Q(pp_row38_21));
 sky130_fd_sc_hd__dfxtp_1 _1527_ (.CLK(clknet_leaf_18_clk),
    .D(booth_b0_m39),
    .Q(pp_row39_0));
 sky130_fd_sc_hd__dfxtp_1 _1528_ (.CLK(clknet_leaf_121_clk),
    .D(booth_b46_m59),
    .Q(pp_row105_3));
 sky130_fd_sc_hd__dfxtp_1 _1529_ (.CLK(clknet_leaf_18_clk),
    .D(booth_b2_m37),
    .Q(pp_row39_1));
 sky130_fd_sc_hd__dfxtp_1 _1530_ (.CLK(clknet_leaf_17_clk),
    .D(booth_b4_m35),
    .Q(pp_row39_2));
 sky130_fd_sc_hd__dfxtp_1 _1531_ (.CLK(clknet_leaf_44_clk),
    .D(booth_b6_m33),
    .Q(pp_row39_3));
 sky130_fd_sc_hd__dfxtp_1 _1532_ (.CLK(clknet_leaf_44_clk),
    .D(booth_b8_m31),
    .Q(pp_row39_4));
 sky130_fd_sc_hd__dfxtp_1 _1533_ (.CLK(clknet_leaf_44_clk),
    .D(booth_b10_m29),
    .Q(pp_row39_5));
 sky130_fd_sc_hd__dfxtp_1 _1534_ (.CLK(clknet_leaf_16_clk),
    .D(booth_b12_m27),
    .Q(pp_row39_6));
 sky130_fd_sc_hd__dfxtp_1 _1535_ (.CLK(clknet_leaf_16_clk),
    .D(booth_b14_m25),
    .Q(pp_row39_7));
 sky130_fd_sc_hd__dfxtp_1 _1536_ (.CLK(clknet_leaf_8_clk),
    .D(booth_b16_m23),
    .Q(pp_row39_8));
 sky130_fd_sc_hd__dfxtp_1 _1537_ (.CLK(clknet_leaf_7_clk),
    .D(booth_b18_m21),
    .Q(pp_row39_9));
 sky130_fd_sc_hd__dfxtp_1 _1538_ (.CLK(clknet_leaf_8_clk),
    .D(booth_b20_m19),
    .Q(pp_row39_10));
 sky130_fd_sc_hd__dfxtp_1 _1539_ (.CLK(clknet_leaf_121_clk),
    .D(booth_b48_m57),
    .Q(pp_row105_4));
 sky130_fd_sc_hd__dfxtp_1 _1540_ (.CLK(clknet_leaf_12_clk),
    .D(booth_b22_m17),
    .Q(pp_row39_11));
 sky130_fd_sc_hd__dfxtp_1 _1541_ (.CLK(clknet_leaf_8_clk),
    .D(booth_b24_m15),
    .Q(pp_row39_12));
 sky130_fd_sc_hd__dfxtp_1 _1542_ (.CLK(clknet_leaf_12_clk),
    .D(booth_b26_m13),
    .Q(pp_row39_13));
 sky130_fd_sc_hd__dfxtp_1 _1543_ (.CLK(clknet_leaf_16_clk),
    .D(booth_b28_m11),
    .Q(pp_row39_14));
 sky130_fd_sc_hd__dfxtp_1 _1544_ (.CLK(clknet_leaf_16_clk),
    .D(booth_b30_m9),
    .Q(pp_row39_15));
 sky130_fd_sc_hd__dfxtp_1 _1545_ (.CLK(clknet_leaf_17_clk),
    .D(booth_b32_m7),
    .Q(pp_row39_16));
 sky130_fd_sc_hd__dfxtp_1 _1546_ (.CLK(clknet_leaf_20_clk),
    .D(booth_b34_m5),
    .Q(pp_row39_17));
 sky130_fd_sc_hd__dfxtp_1 _1547_ (.CLK(clknet_leaf_19_clk),
    .D(booth_b36_m3),
    .Q(pp_row39_18));
 sky130_fd_sc_hd__dfxtp_1 _1548_ (.CLK(clknet_leaf_19_clk),
    .D(booth_b38_m1),
    .Q(pp_row39_19));
 sky130_fd_sc_hd__dfxtp_2 _1549_ (.CLK(clknet_leaf_236_clk),
    .D(net189),
    .Q(pp_row39_20));
 sky130_fd_sc_hd__dfxtp_1 _1550_ (.CLK(clknet_leaf_121_clk),
    .D(booth_b50_m55),
    .Q(pp_row105_5));
 sky130_fd_sc_hd__dfxtp_1 _1551_ (.CLK(clknet_leaf_240_clk),
    .D(booth_b0_m40),
    .Q(pp_row40_0));
 sky130_fd_sc_hd__dfxtp_1 _1552_ (.CLK(clknet_leaf_5_clk),
    .D(booth_b2_m38),
    .Q(pp_row40_1));
 sky130_fd_sc_hd__dfxtp_1 _1553_ (.CLK(clknet_leaf_5_clk),
    .D(booth_b4_m36),
    .Q(pp_row40_2));
 sky130_fd_sc_hd__dfxtp_1 _1554_ (.CLK(clknet_leaf_6_clk),
    .D(booth_b6_m34),
    .Q(pp_row40_3));
 sky130_fd_sc_hd__dfxtp_1 _1555_ (.CLK(clknet_leaf_7_clk),
    .D(booth_b8_m32),
    .Q(pp_row40_4));
 sky130_fd_sc_hd__dfxtp_1 _1556_ (.CLK(clknet_leaf_9_clk),
    .D(booth_b10_m30),
    .Q(pp_row40_5));
 sky130_fd_sc_hd__dfxtp_1 _1557_ (.CLK(clknet_leaf_9_clk),
    .D(booth_b12_m28),
    .Q(pp_row40_6));
 sky130_fd_sc_hd__dfxtp_1 _1558_ (.CLK(clknet_leaf_7_clk),
    .D(booth_b14_m26),
    .Q(pp_row40_7));
 sky130_fd_sc_hd__dfxtp_1 _1559_ (.CLK(clknet_leaf_7_clk),
    .D(booth_b16_m24),
    .Q(pp_row40_8));
 sky130_fd_sc_hd__dfxtp_1 _1560_ (.CLK(clknet_leaf_7_clk),
    .D(booth_b18_m22),
    .Q(pp_row40_9));
 sky130_fd_sc_hd__dfxtp_1 _1561_ (.CLK(clknet_leaf_108_clk),
    .D(booth_b52_m53),
    .Q(pp_row105_6));
 sky130_fd_sc_hd__dfxtp_1 _1562_ (.CLK(clknet_leaf_7_clk),
    .D(booth_b20_m20),
    .Q(pp_row40_10));
 sky130_fd_sc_hd__dfxtp_1 _1563_ (.CLK(clknet_leaf_7_clk),
    .D(booth_b22_m18),
    .Q(pp_row40_11));
 sky130_fd_sc_hd__dfxtp_1 _1564_ (.CLK(clknet_leaf_8_clk),
    .D(booth_b24_m16),
    .Q(pp_row40_12));
 sky130_fd_sc_hd__dfxtp_1 _1565_ (.CLK(clknet_leaf_8_clk),
    .D(booth_b26_m14),
    .Q(pp_row40_13));
 sky130_fd_sc_hd__dfxtp_1 _1566_ (.CLK(clknet_leaf_7_clk),
    .D(booth_b28_m12),
    .Q(pp_row40_14));
 sky130_fd_sc_hd__dfxtp_1 _1567_ (.CLK(clknet_leaf_7_clk),
    .D(booth_b30_m10),
    .Q(pp_row40_15));
 sky130_fd_sc_hd__dfxtp_1 _1568_ (.CLK(clknet_leaf_7_clk),
    .D(booth_b32_m8),
    .Q(pp_row40_16));
 sky130_fd_sc_hd__dfxtp_1 _1569_ (.CLK(clknet_leaf_20_clk),
    .D(booth_b34_m6),
    .Q(pp_row40_17));
 sky130_fd_sc_hd__dfxtp_1 _1570_ (.CLK(clknet_leaf_19_clk),
    .D(booth_b36_m4),
    .Q(pp_row40_18));
 sky130_fd_sc_hd__dfxtp_1 _1571_ (.CLK(clknet_leaf_20_clk),
    .D(booth_b38_m2),
    .Q(pp_row40_19));
 sky130_fd_sc_hd__dfxtp_1 _1572_ (.CLK(clknet_leaf_108_clk),
    .D(booth_b54_m51),
    .Q(pp_row105_7));
 sky130_fd_sc_hd__dfxtp_1 _1573_ (.CLK(clknet_leaf_21_clk),
    .D(booth_b40_m0),
    .Q(pp_row40_20));
 sky130_fd_sc_hd__dfxtp_1 _1574_ (.CLK(clknet_leaf_21_clk),
    .D(net1376),
    .Q(pp_row40_21));
 sky130_fd_sc_hd__dfxtp_1 _1575_ (.CLK(clknet_leaf_244_clk),
    .D(net191),
    .Q(pp_row40_22));
 sky130_fd_sc_hd__dfxtp_1 _1576_ (.CLK(clknet_leaf_243_clk),
    .D(booth_b0_m41),
    .Q(pp_row41_0));
 sky130_fd_sc_hd__dfxtp_1 _1577_ (.CLK(clknet_leaf_243_clk),
    .D(booth_b2_m39),
    .Q(pp_row41_1));
 sky130_fd_sc_hd__dfxtp_1 _1578_ (.CLK(clknet_leaf_243_clk),
    .D(booth_b4_m37),
    .Q(pp_row41_2));
 sky130_fd_sc_hd__dfxtp_1 _1579_ (.CLK(clknet_leaf_243_clk),
    .D(booth_b6_m35),
    .Q(pp_row41_3));
 sky130_fd_sc_hd__dfxtp_1 _1580_ (.CLK(clknet_leaf_243_clk),
    .D(booth_b8_m33),
    .Q(pp_row41_4));
 sky130_fd_sc_hd__dfxtp_1 _1581_ (.CLK(clknet_leaf_243_clk),
    .D(booth_b10_m31),
    .Q(pp_row41_5));
 sky130_fd_sc_hd__dfxtp_1 _1582_ (.CLK(clknet_leaf_242_clk),
    .D(booth_b12_m29),
    .Q(pp_row41_6));
 sky130_fd_sc_hd__dfxtp_1 _1583_ (.CLK(clknet_leaf_109_clk),
    .D(booth_b56_m49),
    .Q(pp_row105_8));
 sky130_fd_sc_hd__dfxtp_1 _1584_ (.CLK(clknet_leaf_243_clk),
    .D(booth_b14_m27),
    .Q(pp_row41_7));
 sky130_fd_sc_hd__dfxtp_1 _1585_ (.CLK(clknet_leaf_243_clk),
    .D(booth_b16_m25),
    .Q(pp_row41_8));
 sky130_fd_sc_hd__dfxtp_1 _1586_ (.CLK(clknet_leaf_4_clk),
    .D(booth_b18_m23),
    .Q(pp_row41_9));
 sky130_fd_sc_hd__dfxtp_1 _1587_ (.CLK(clknet_leaf_4_clk),
    .D(booth_b20_m21),
    .Q(pp_row41_10));
 sky130_fd_sc_hd__dfxtp_1 _1588_ (.CLK(clknet_leaf_9_clk),
    .D(booth_b22_m19),
    .Q(pp_row41_11));
 sky130_fd_sc_hd__dfxtp_1 _1589_ (.CLK(clknet_leaf_9_clk),
    .D(booth_b24_m17),
    .Q(pp_row41_12));
 sky130_fd_sc_hd__dfxtp_1 _1590_ (.CLK(clknet_leaf_9_clk),
    .D(booth_b26_m15),
    .Q(pp_row41_13));
 sky130_fd_sc_hd__dfxtp_1 _1591_ (.CLK(clknet_leaf_5_clk),
    .D(booth_b28_m13),
    .Q(pp_row41_14));
 sky130_fd_sc_hd__dfxtp_1 _1592_ (.CLK(clknet_leaf_5_clk),
    .D(booth_b30_m11),
    .Q(pp_row41_15));
 sky130_fd_sc_hd__dfxtp_1 _1593_ (.CLK(clknet_leaf_6_clk),
    .D(booth_b32_m9),
    .Q(pp_row41_16));
 sky130_fd_sc_hd__dfxtp_1 _1594_ (.CLK(clknet_leaf_110_clk),
    .D(booth_b58_m47),
    .Q(pp_row105_9));
 sky130_fd_sc_hd__dfxtp_1 _1595_ (.CLK(clknet_leaf_5_clk),
    .D(booth_b34_m7),
    .Q(pp_row41_17));
 sky130_fd_sc_hd__dfxtp_1 _1596_ (.CLK(clknet_leaf_5_clk),
    .D(booth_b36_m5),
    .Q(pp_row41_18));
 sky130_fd_sc_hd__dfxtp_1 _1597_ (.CLK(clknet_leaf_5_clk),
    .D(booth_b38_m3),
    .Q(pp_row41_19));
 sky130_fd_sc_hd__dfxtp_1 _1598_ (.CLK(clknet_leaf_5_clk),
    .D(booth_b40_m1),
    .Q(pp_row41_20));
 sky130_fd_sc_hd__dfxtp_1 _1599_ (.CLK(clknet_leaf_244_clk),
    .D(net192),
    .Q(pp_row41_21));
 sky130_fd_sc_hd__dfxtp_1 _1600_ (.CLK(clknet_leaf_237_clk),
    .D(booth_b0_m42),
    .Q(pp_row42_0));
 sky130_fd_sc_hd__dfxtp_1 _1601_ (.CLK(clknet_leaf_243_clk),
    .D(booth_b2_m40),
    .Q(pp_row42_1));
 sky130_fd_sc_hd__dfxtp_1 _1602_ (.CLK(clknet_leaf_243_clk),
    .D(booth_b4_m38),
    .Q(pp_row42_2));
 sky130_fd_sc_hd__dfxtp_1 _1603_ (.CLK(clknet_leaf_240_clk),
    .D(booth_b6_m36),
    .Q(pp_row42_3));
 sky130_fd_sc_hd__dfxtp_1 _1604_ (.CLK(clknet_leaf_240_clk),
    .D(booth_b8_m34),
    .Q(pp_row42_4));
 sky130_fd_sc_hd__dfxtp_1 _1605_ (.CLK(clknet_leaf_110_clk),
    .D(booth_b60_m45),
    .Q(pp_row105_10));
 sky130_fd_sc_hd__dfxtp_1 _1606_ (.CLK(clknet_leaf_240_clk),
    .D(booth_b10_m32),
    .Q(pp_row42_5));
 sky130_fd_sc_hd__dfxtp_1 _1607_ (.CLK(clknet_leaf_240_clk),
    .D(booth_b12_m30),
    .Q(pp_row42_6));
 sky130_fd_sc_hd__dfxtp_1 _1608_ (.CLK(clknet_leaf_240_clk),
    .D(booth_b14_m28),
    .Q(pp_row42_7));
 sky130_fd_sc_hd__dfxtp_1 _1609_ (.CLK(clknet_leaf_240_clk),
    .D(booth_b16_m26),
    .Q(pp_row42_8));
 sky130_fd_sc_hd__dfxtp_1 _1610_ (.CLK(clknet_leaf_239_clk),
    .D(booth_b18_m24),
    .Q(pp_row42_9));
 sky130_fd_sc_hd__dfxtp_1 _1611_ (.CLK(clknet_leaf_239_clk),
    .D(booth_b20_m22),
    .Q(pp_row42_10));
 sky130_fd_sc_hd__dfxtp_1 _1612_ (.CLK(clknet_leaf_239_clk),
    .D(booth_b22_m20),
    .Q(pp_row42_11));
 sky130_fd_sc_hd__dfxtp_1 _1613_ (.CLK(clknet_leaf_239_clk),
    .D(booth_b24_m18),
    .Q(pp_row42_12));
 sky130_fd_sc_hd__dfxtp_1 _1614_ (.CLK(clknet_leaf_239_clk),
    .D(booth_b26_m16),
    .Q(pp_row42_13));
 sky130_fd_sc_hd__dfxtp_1 _1615_ (.CLK(clknet_leaf_241_clk),
    .D(booth_b28_m14),
    .Q(pp_row42_14));
 sky130_fd_sc_hd__dfxtp_1 _1616_ (.CLK(clknet_leaf_110_clk),
    .D(booth_b62_m43),
    .Q(pp_row105_11));
 sky130_fd_sc_hd__dfxtp_1 _1617_ (.CLK(clknet_leaf_164_clk),
    .D(booth_b62_m61),
    .Q(pp_row123_2));
 sky130_fd_sc_hd__dfxtp_1 _1618_ (.CLK(clknet_leaf_241_clk),
    .D(booth_b30_m12),
    .Q(pp_row42_15));
 sky130_fd_sc_hd__dfxtp_1 _1619_ (.CLK(clknet_leaf_240_clk),
    .D(booth_b32_m10),
    .Q(pp_row42_16));
 sky130_fd_sc_hd__dfxtp_1 _1620_ (.CLK(clknet_leaf_5_clk),
    .D(booth_b34_m8),
    .Q(pp_row42_17));
 sky130_fd_sc_hd__dfxtp_1 _1621_ (.CLK(clknet_leaf_5_clk),
    .D(booth_b36_m6),
    .Q(pp_row42_18));
 sky130_fd_sc_hd__dfxtp_1 _1622_ (.CLK(clknet_leaf_5_clk),
    .D(booth_b38_m4),
    .Q(pp_row42_19));
 sky130_fd_sc_hd__dfxtp_1 _1623_ (.CLK(clknet_leaf_240_clk),
    .D(booth_b40_m2),
    .Q(pp_row42_20));
 sky130_fd_sc_hd__dfxtp_1 _1624_ (.CLK(clknet_leaf_239_clk),
    .D(booth_b42_m0),
    .Q(pp_row42_21));
 sky130_fd_sc_hd__dfxtp_1 _1625_ (.CLK(clknet_leaf_239_clk),
    .D(net1367),
    .Q(pp_row42_22));
 sky130_fd_sc_hd__dfxtp_1 _1626_ (.CLK(clknet_leaf_236_clk),
    .D(net193),
    .Q(pp_row42_23));
 sky130_fd_sc_hd__dfxtp_1 _1627_ (.CLK(clknet_leaf_221_clk),
    .D(booth_b0_m43),
    .Q(pp_row43_0));
 sky130_fd_sc_hd__dfxtp_1 _1628_ (.CLK(clknet_leaf_121_clk),
    .D(booth_b64_m41),
    .Q(pp_row105_12));
 sky130_fd_sc_hd__dfxtp_1 _1629_ (.CLK(clknet_leaf_221_clk),
    .D(booth_b2_m41),
    .Q(pp_row43_1));
 sky130_fd_sc_hd__dfxtp_1 _1630_ (.CLK(clknet_leaf_239_clk),
    .D(booth_b4_m39),
    .Q(pp_row43_2));
 sky130_fd_sc_hd__dfxtp_1 _1631_ (.CLK(clknet_leaf_246_clk),
    .D(booth_b6_m37),
    .Q(pp_row43_3));
 sky130_fd_sc_hd__dfxtp_1 _1632_ (.CLK(clknet_leaf_242_clk),
    .D(booth_b8_m35),
    .Q(pp_row43_4));
 sky130_fd_sc_hd__dfxtp_1 _1633_ (.CLK(clknet_leaf_242_clk),
    .D(booth_b10_m33),
    .Q(pp_row43_5));
 sky130_fd_sc_hd__dfxtp_1 _1634_ (.CLK(clknet_leaf_239_clk),
    .D(booth_b12_m31),
    .Q(pp_row43_6));
 sky130_fd_sc_hd__dfxtp_1 _1635_ (.CLK(clknet_leaf_239_clk),
    .D(booth_b14_m29),
    .Q(pp_row43_7));
 sky130_fd_sc_hd__dfxtp_1 _1636_ (.CLK(clknet_leaf_223_clk),
    .D(booth_b16_m27),
    .Q(pp_row43_8));
 sky130_fd_sc_hd__dfxtp_1 _1637_ (.CLK(clknet_leaf_240_clk),
    .D(booth_b18_m25),
    .Q(pp_row43_9));
 sky130_fd_sc_hd__dfxtp_1 _1638_ (.CLK(clknet_leaf_240_clk),
    .D(booth_b20_m23),
    .Q(pp_row43_10));
 sky130_fd_sc_hd__dfxtp_2 _1639_ (.CLK(clknet_leaf_184_clk),
    .D(net135),
    .Q(pp_row105_13));
 sky130_fd_sc_hd__dfxtp_1 _1640_ (.CLK(clknet_leaf_240_clk),
    .D(booth_b22_m21),
    .Q(pp_row43_11));
 sky130_fd_sc_hd__dfxtp_1 _1641_ (.CLK(clknet_leaf_240_clk),
    .D(booth_b24_m19),
    .Q(pp_row43_12));
 sky130_fd_sc_hd__dfxtp_1 _1642_ (.CLK(clknet_leaf_240_clk),
    .D(booth_b26_m17),
    .Q(pp_row43_13));
 sky130_fd_sc_hd__dfxtp_1 _1643_ (.CLK(clknet_leaf_6_clk),
    .D(booth_b28_m15),
    .Q(pp_row43_14));
 sky130_fd_sc_hd__dfxtp_1 _1644_ (.CLK(clknet_leaf_6_clk),
    .D(booth_b30_m13),
    .Q(pp_row43_15));
 sky130_fd_sc_hd__dfxtp_1 _1645_ (.CLK(clknet_leaf_6_clk),
    .D(booth_b32_m11),
    .Q(pp_row43_16));
 sky130_fd_sc_hd__dfxtp_1 _1646_ (.CLK(clknet_leaf_6_clk),
    .D(booth_b34_m9),
    .Q(pp_row43_17));
 sky130_fd_sc_hd__dfxtp_1 _1647_ (.CLK(clknet_leaf_5_clk),
    .D(booth_b36_m7),
    .Q(pp_row43_18));
 sky130_fd_sc_hd__dfxtp_1 _1648_ (.CLK(clknet_leaf_5_clk),
    .D(booth_b38_m5),
    .Q(pp_row43_19));
 sky130_fd_sc_hd__dfxtp_1 _1649_ (.CLK(clknet_leaf_239_clk),
    .D(booth_b40_m3),
    .Q(pp_row43_20));
 sky130_fd_sc_hd__dfxtp_1 _1650_ (.CLK(clknet_leaf_124_clk),
    .D(booth_b42_m64),
    .Q(pp_row106_1));
 sky130_fd_sc_hd__dfxtp_1 _1651_ (.CLK(clknet_leaf_239_clk),
    .D(booth_b42_m1),
    .Q(pp_row43_21));
 sky130_fd_sc_hd__dfxtp_1 _1652_ (.CLK(clknet_leaf_235_clk),
    .D(net194),
    .Q(pp_row43_22));
 sky130_fd_sc_hd__dfxtp_1 _1653_ (.CLK(clknet_leaf_221_clk),
    .D(booth_b0_m44),
    .Q(pp_row44_0));
 sky130_fd_sc_hd__dfxtp_1 _1654_ (.CLK(clknet_leaf_221_clk),
    .D(booth_b2_m42),
    .Q(pp_row44_1));
 sky130_fd_sc_hd__dfxtp_1 _1655_ (.CLK(clknet_leaf_221_clk),
    .D(booth_b4_m40),
    .Q(pp_row44_2));
 sky130_fd_sc_hd__dfxtp_1 _1656_ (.CLK(clknet_leaf_6_clk),
    .D(booth_b6_m38),
    .Q(pp_row44_3));
 sky130_fd_sc_hd__dfxtp_1 _1657_ (.CLK(clknet_leaf_6_clk),
    .D(booth_b8_m36),
    .Q(pp_row44_4));
 sky130_fd_sc_hd__dfxtp_1 _1658_ (.CLK(clknet_leaf_6_clk),
    .D(booth_b10_m34),
    .Q(pp_row44_5));
 sky130_fd_sc_hd__dfxtp_1 _1659_ (.CLK(clknet_leaf_21_clk),
    .D(booth_b12_m32),
    .Q(pp_row44_6));
 sky130_fd_sc_hd__dfxtp_1 _1660_ (.CLK(clknet_leaf_21_clk),
    .D(booth_b14_m30),
    .Q(pp_row44_7));
 sky130_fd_sc_hd__dfxtp_1 _1661_ (.CLK(clknet_leaf_124_clk),
    .D(booth_b44_m62),
    .Q(pp_row106_2));
 sky130_fd_sc_hd__dfxtp_1 _1662_ (.CLK(clknet_leaf_21_clk),
    .D(booth_b16_m28),
    .Q(pp_row44_8));
 sky130_fd_sc_hd__dfxtp_1 _1663_ (.CLK(clknet_leaf_24_clk),
    .D(booth_b18_m26),
    .Q(pp_row44_9));
 sky130_fd_sc_hd__dfxtp_1 _1664_ (.CLK(clknet_leaf_24_clk),
    .D(booth_b20_m24),
    .Q(pp_row44_10));
 sky130_fd_sc_hd__dfxtp_1 _1665_ (.CLK(clknet_leaf_24_clk),
    .D(booth_b22_m22),
    .Q(pp_row44_11));
 sky130_fd_sc_hd__dfxtp_1 _1666_ (.CLK(clknet_leaf_21_clk),
    .D(booth_b24_m20),
    .Q(pp_row44_12));
 sky130_fd_sc_hd__dfxtp_1 _1667_ (.CLK(clknet_leaf_21_clk),
    .D(booth_b26_m18),
    .Q(pp_row44_13));
 sky130_fd_sc_hd__dfxtp_1 _1668_ (.CLK(clknet_leaf_20_clk),
    .D(booth_b28_m16),
    .Q(pp_row44_14));
 sky130_fd_sc_hd__dfxtp_1 _1669_ (.CLK(clknet_leaf_19_clk),
    .D(booth_b30_m14),
    .Q(pp_row44_15));
 sky130_fd_sc_hd__dfxtp_1 _1670_ (.CLK(clknet_leaf_19_clk),
    .D(booth_b32_m12),
    .Q(pp_row44_16));
 sky130_fd_sc_hd__dfxtp_1 _1671_ (.CLK(clknet_leaf_241_clk),
    .D(booth_b34_m10),
    .Q(pp_row44_17));
 sky130_fd_sc_hd__dfxtp_1 _1672_ (.CLK(clknet_leaf_123_clk),
    .D(booth_b46_m60),
    .Q(pp_row106_3));
 sky130_fd_sc_hd__dfxtp_1 _1673_ (.CLK(clknet_leaf_4_clk),
    .D(booth_b36_m8),
    .Q(pp_row44_18));
 sky130_fd_sc_hd__dfxtp_1 _1674_ (.CLK(clknet_leaf_240_clk),
    .D(booth_b38_m6),
    .Q(pp_row44_19));
 sky130_fd_sc_hd__dfxtp_1 _1675_ (.CLK(clknet_leaf_22_clk),
    .D(booth_b40_m4),
    .Q(pp_row44_20));
 sky130_fd_sc_hd__dfxtp_1 _1676_ (.CLK(clknet_leaf_22_clk),
    .D(booth_b42_m2),
    .Q(pp_row44_21));
 sky130_fd_sc_hd__dfxtp_1 _1677_ (.CLK(clknet_leaf_22_clk),
    .D(booth_b44_m0),
    .Q(pp_row44_22));
 sky130_fd_sc_hd__dfxtp_1 _1678_ (.CLK(clknet_leaf_239_clk),
    .D(net1357),
    .Q(pp_row44_23));
 sky130_fd_sc_hd__dfxtp_1 _1679_ (.CLK(clknet_leaf_235_clk),
    .D(net195),
    .Q(pp_row44_24));
 sky130_fd_sc_hd__dfxtp_1 _1680_ (.CLK(clknet_leaf_24_clk),
    .D(booth_b0_m45),
    .Q(pp_row45_0));
 sky130_fd_sc_hd__dfxtp_1 _1681_ (.CLK(clknet_leaf_24_clk),
    .D(booth_b2_m43),
    .Q(pp_row45_1));
 sky130_fd_sc_hd__dfxtp_1 _1682_ (.CLK(clknet_leaf_24_clk),
    .D(booth_b4_m41),
    .Q(pp_row45_2));
 sky130_fd_sc_hd__dfxtp_1 _1683_ (.CLK(clknet_leaf_123_clk),
    .D(booth_b48_m58),
    .Q(pp_row106_4));
 sky130_fd_sc_hd__dfxtp_1 _1684_ (.CLK(clknet_leaf_19_clk),
    .D(booth_b6_m39),
    .Q(pp_row45_3));
 sky130_fd_sc_hd__dfxtp_1 _1685_ (.CLK(clknet_leaf_19_clk),
    .D(booth_b8_m37),
    .Q(pp_row45_4));
 sky130_fd_sc_hd__dfxtp_1 _1686_ (.CLK(clknet_leaf_19_clk),
    .D(booth_b10_m35),
    .Q(pp_row45_5));
 sky130_fd_sc_hd__dfxtp_1 _1687_ (.CLK(clknet_leaf_25_clk),
    .D(booth_b12_m33),
    .Q(pp_row45_6));
 sky130_fd_sc_hd__dfxtp_1 _1688_ (.CLK(clknet_leaf_18_clk),
    .D(booth_b14_m31),
    .Q(pp_row45_7));
 sky130_fd_sc_hd__dfxtp_1 _1689_ (.CLK(clknet_leaf_18_clk),
    .D(booth_b16_m29),
    .Q(pp_row45_8));
 sky130_fd_sc_hd__dfxtp_1 _1690_ (.CLK(clknet_leaf_19_clk),
    .D(booth_b18_m27),
    .Q(pp_row45_9));
 sky130_fd_sc_hd__dfxtp_1 _1691_ (.CLK(clknet_leaf_19_clk),
    .D(booth_b20_m25),
    .Q(pp_row45_10));
 sky130_fd_sc_hd__dfxtp_1 _1692_ (.CLK(clknet_leaf_19_clk),
    .D(booth_b22_m23),
    .Q(pp_row45_11));
 sky130_fd_sc_hd__dfxtp_1 _1693_ (.CLK(clknet_leaf_18_clk),
    .D(booth_b24_m21),
    .Q(pp_row45_12));
 sky130_fd_sc_hd__dfxtp_1 _1694_ (.CLK(clknet_leaf_123_clk),
    .D(booth_b50_m56),
    .Q(pp_row106_5));
 sky130_fd_sc_hd__dfxtp_1 _1695_ (.CLK(clknet_leaf_18_clk),
    .D(booth_b26_m19),
    .Q(pp_row45_13));
 sky130_fd_sc_hd__dfxtp_1 _1696_ (.CLK(clknet_leaf_18_clk),
    .D(booth_b28_m17),
    .Q(pp_row45_14));
 sky130_fd_sc_hd__dfxtp_1 _1697_ (.CLK(clknet_leaf_19_clk),
    .D(booth_b30_m15),
    .Q(pp_row45_15));
 sky130_fd_sc_hd__dfxtp_1 _1698_ (.CLK(clknet_leaf_19_clk),
    .D(booth_b32_m13),
    .Q(pp_row45_16));
 sky130_fd_sc_hd__dfxtp_1 _1699_ (.CLK(clknet_leaf_23_clk),
    .D(booth_b34_m11),
    .Q(pp_row45_17));
 sky130_fd_sc_hd__dfxtp_1 _1700_ (.CLK(clknet_leaf_22_clk),
    .D(booth_b36_m9),
    .Q(pp_row45_18));
 sky130_fd_sc_hd__dfxtp_1 _1701_ (.CLK(clknet_leaf_22_clk),
    .D(booth_b38_m7),
    .Q(pp_row45_19));
 sky130_fd_sc_hd__dfxtp_1 _1702_ (.CLK(clknet_leaf_23_clk),
    .D(booth_b40_m5),
    .Q(pp_row45_20));
 sky130_fd_sc_hd__dfxtp_1 _1703_ (.CLK(clknet_leaf_23_clk),
    .D(booth_b42_m3),
    .Q(pp_row45_21));
 sky130_fd_sc_hd__dfxtp_1 _1704_ (.CLK(clknet_leaf_23_clk),
    .D(booth_b44_m1),
    .Q(pp_row45_22));
 sky130_fd_sc_hd__dfxtp_1 _1705_ (.CLK(clknet_leaf_123_clk),
    .D(booth_b52_m54),
    .Q(pp_row106_6));
 sky130_fd_sc_hd__dfxtp_1 _1706_ (.CLK(clknet_leaf_236_clk),
    .D(net196),
    .Q(pp_row45_23));
 sky130_fd_sc_hd__dfxtp_1 _1707_ (.CLK(clknet_leaf_236_clk),
    .D(booth_b0_m46),
    .Q(pp_row46_0));
 sky130_fd_sc_hd__dfxtp_1 _1708_ (.CLK(clknet_leaf_236_clk),
    .D(booth_b2_m44),
    .Q(pp_row46_1));
 sky130_fd_sc_hd__dfxtp_1 _1709_ (.CLK(clknet_leaf_236_clk),
    .D(booth_b4_m42),
    .Q(pp_row46_2));
 sky130_fd_sc_hd__dfxtp_1 _1710_ (.CLK(clknet_leaf_236_clk),
    .D(booth_b6_m40),
    .Q(pp_row46_3));
 sky130_fd_sc_hd__dfxtp_1 _1711_ (.CLK(clknet_leaf_237_clk),
    .D(booth_b8_m38),
    .Q(pp_row46_4));
 sky130_fd_sc_hd__dfxtp_1 _1712_ (.CLK(clknet_leaf_236_clk),
    .D(booth_b10_m36),
    .Q(pp_row46_5));
 sky130_fd_sc_hd__dfxtp_1 _1713_ (.CLK(clknet_leaf_237_clk),
    .D(booth_b12_m34),
    .Q(pp_row46_6));
 sky130_fd_sc_hd__dfxtp_1 _1714_ (.CLK(clknet_leaf_237_clk),
    .D(booth_b14_m32),
    .Q(pp_row46_7));
 sky130_fd_sc_hd__dfxtp_1 _1715_ (.CLK(clknet_leaf_237_clk),
    .D(booth_b16_m30),
    .Q(pp_row46_8));
 sky130_fd_sc_hd__dfxtp_1 _1716_ (.CLK(clknet_leaf_138_clk),
    .D(booth_b54_m52),
    .Q(pp_row106_7));
 sky130_fd_sc_hd__dfxtp_1 _1717_ (.CLK(clknet_leaf_21_clk),
    .D(booth_b18_m28),
    .Q(pp_row46_9));
 sky130_fd_sc_hd__dfxtp_1 _1718_ (.CLK(clknet_leaf_21_clk),
    .D(booth_b20_m26),
    .Q(pp_row46_10));
 sky130_fd_sc_hd__dfxtp_1 _1719_ (.CLK(clknet_leaf_21_clk),
    .D(booth_b22_m24),
    .Q(pp_row46_11));
 sky130_fd_sc_hd__dfxtp_1 _1720_ (.CLK(clknet_leaf_22_clk),
    .D(booth_b24_m22),
    .Q(pp_row46_12));
 sky130_fd_sc_hd__dfxtp_1 _1721_ (.CLK(clknet_leaf_22_clk),
    .D(booth_b26_m20),
    .Q(pp_row46_13));
 sky130_fd_sc_hd__dfxtp_1 _1722_ (.CLK(clknet_leaf_22_clk),
    .D(booth_b28_m18),
    .Q(pp_row46_14));
 sky130_fd_sc_hd__dfxtp_1 _1723_ (.CLK(clknet_leaf_21_clk),
    .D(booth_b30_m16),
    .Q(pp_row46_15));
 sky130_fd_sc_hd__dfxtp_1 _1724_ (.CLK(clknet_leaf_22_clk),
    .D(booth_b32_m14),
    .Q(pp_row46_16));
 sky130_fd_sc_hd__dfxtp_1 _1725_ (.CLK(clknet_leaf_21_clk),
    .D(booth_b34_m12),
    .Q(pp_row46_17));
 sky130_fd_sc_hd__dfxtp_1 _1726_ (.CLK(clknet_leaf_23_clk),
    .D(booth_b36_m10),
    .Q(pp_row46_18));
 sky130_fd_sc_hd__dfxtp_1 _1727_ (.CLK(clknet_leaf_123_clk),
    .D(booth_b56_m50),
    .Q(pp_row106_8));
 sky130_fd_sc_hd__dfxtp_1 _1728_ (.CLK(clknet_leaf_164_clk),
    .D(booth_b64_m59),
    .Q(pp_row123_3));
 sky130_fd_sc_hd__dfxtp_1 _1729_ (.CLK(clknet_leaf_21_clk),
    .D(booth_b38_m8),
    .Q(pp_row46_19));
 sky130_fd_sc_hd__dfxtp_1 _1730_ (.CLK(clknet_leaf_24_clk),
    .D(booth_b40_m6),
    .Q(pp_row46_20));
 sky130_fd_sc_hd__dfxtp_1 _1731_ (.CLK(clknet_leaf_24_clk),
    .D(booth_b42_m4),
    .Q(pp_row46_21));
 sky130_fd_sc_hd__dfxtp_1 _1732_ (.CLK(clknet_leaf_24_clk),
    .D(booth_b44_m2),
    .Q(pp_row46_22));
 sky130_fd_sc_hd__dfxtp_1 _1733_ (.CLK(clknet_leaf_24_clk),
    .D(booth_b46_m0),
    .Q(pp_row46_23));
 sky130_fd_sc_hd__dfxtp_1 _1734_ (.CLK(clknet_leaf_23_clk),
    .D(net1348),
    .Q(pp_row46_24));
 sky130_fd_sc_hd__dfxtp_1 _1735_ (.CLK(clknet_leaf_235_clk),
    .D(net197),
    .Q(pp_row46_25));
 sky130_fd_sc_hd__dfxtp_1 _1736_ (.CLK(clknet_leaf_236_clk),
    .D(booth_b0_m47),
    .Q(pp_row47_0));
 sky130_fd_sc_hd__dfxtp_1 _1737_ (.CLK(clknet_leaf_236_clk),
    .D(booth_b2_m45),
    .Q(pp_row47_1));
 sky130_fd_sc_hd__dfxtp_1 _1738_ (.CLK(clknet_leaf_236_clk),
    .D(booth_b4_m43),
    .Q(pp_row47_2));
 sky130_fd_sc_hd__dfxtp_1 _1739_ (.CLK(clknet_leaf_122_clk),
    .D(booth_b58_m48),
    .Q(pp_row106_9));
 sky130_fd_sc_hd__dfxtp_1 _1740_ (.CLK(clknet_leaf_236_clk),
    .D(booth_b6_m41),
    .Q(pp_row47_3));
 sky130_fd_sc_hd__dfxtp_1 _1741_ (.CLK(clknet_leaf_237_clk),
    .D(booth_b8_m39),
    .Q(pp_row47_4));
 sky130_fd_sc_hd__dfxtp_1 _1742_ (.CLK(clknet_leaf_237_clk),
    .D(booth_b10_m37),
    .Q(pp_row47_5));
 sky130_fd_sc_hd__dfxtp_1 _1743_ (.CLK(clknet_leaf_237_clk),
    .D(booth_b12_m35),
    .Q(pp_row47_6));
 sky130_fd_sc_hd__dfxtp_1 _1744_ (.CLK(clknet_leaf_237_clk),
    .D(booth_b14_m33),
    .Q(pp_row47_7));
 sky130_fd_sc_hd__dfxtp_1 _1745_ (.CLK(clknet_leaf_237_clk),
    .D(booth_b16_m31),
    .Q(pp_row47_8));
 sky130_fd_sc_hd__dfxtp_1 _1746_ (.CLK(clknet_leaf_234_clk),
    .D(booth_b18_m29),
    .Q(pp_row47_9));
 sky130_fd_sc_hd__dfxtp_1 _1747_ (.CLK(clknet_leaf_238_clk),
    .D(booth_b20_m27),
    .Q(pp_row47_10));
 sky130_fd_sc_hd__dfxtp_1 _1748_ (.CLK(clknet_leaf_238_clk),
    .D(booth_b22_m25),
    .Q(pp_row47_11));
 sky130_fd_sc_hd__dfxtp_1 _1749_ (.CLK(clknet_leaf_234_clk),
    .D(booth_b24_m23),
    .Q(pp_row47_12));
 sky130_fd_sc_hd__dfxtp_1 _1750_ (.CLK(clknet_leaf_123_clk),
    .D(booth_b60_m46),
    .Q(pp_row106_10));
 sky130_fd_sc_hd__dfxtp_1 _1751_ (.CLK(clknet_leaf_233_clk),
    .D(booth_b26_m21),
    .Q(pp_row47_13));
 sky130_fd_sc_hd__dfxtp_1 _1752_ (.CLK(clknet_leaf_234_clk),
    .D(booth_b28_m19),
    .Q(pp_row47_14));
 sky130_fd_sc_hd__dfxtp_1 _1753_ (.CLK(clknet_leaf_223_clk),
    .D(booth_b30_m17),
    .Q(pp_row47_15));
 sky130_fd_sc_hd__dfxtp_1 _1754_ (.CLK(clknet_leaf_238_clk),
    .D(booth_b32_m15),
    .Q(pp_row47_16));
 sky130_fd_sc_hd__dfxtp_1 _1755_ (.CLK(clknet_leaf_238_clk),
    .D(booth_b34_m13),
    .Q(pp_row47_17));
 sky130_fd_sc_hd__dfxtp_1 _1756_ (.CLK(clknet_leaf_239_clk),
    .D(booth_b36_m11),
    .Q(pp_row47_18));
 sky130_fd_sc_hd__dfxtp_1 _1757_ (.CLK(clknet_leaf_239_clk),
    .D(booth_b38_m9),
    .Q(pp_row47_19));
 sky130_fd_sc_hd__dfxtp_1 _1758_ (.CLK(clknet_leaf_219_clk),
    .D(booth_b40_m7),
    .Q(pp_row47_20));
 sky130_fd_sc_hd__dfxtp_1 _1759_ (.CLK(clknet_leaf_23_clk),
    .D(booth_b42_m5),
    .Q(pp_row47_21));
 sky130_fd_sc_hd__dfxtp_1 _1760_ (.CLK(clknet_leaf_23_clk),
    .D(booth_b44_m3),
    .Q(pp_row47_22));
 sky130_fd_sc_hd__dfxtp_1 _1761_ (.CLK(clknet_leaf_187_clk),
    .D(booth_b62_m44),
    .Q(pp_row106_11));
 sky130_fd_sc_hd__dfxtp_1 _1762_ (.CLK(clknet_leaf_220_clk),
    .D(booth_b46_m1),
    .Q(pp_row47_23));
 sky130_fd_sc_hd__dfxtp_1 _1763_ (.CLK(clknet_leaf_235_clk),
    .D(net198),
    .Q(pp_row47_24));
 sky130_fd_sc_hd__dfxtp_1 _1764_ (.CLK(clknet_leaf_235_clk),
    .D(booth_b0_m48),
    .Q(pp_row48_0));
 sky130_fd_sc_hd__dfxtp_1 _1765_ (.CLK(clknet_leaf_234_clk),
    .D(booth_b2_m46),
    .Q(pp_row48_1));
 sky130_fd_sc_hd__dfxtp_1 _1766_ (.CLK(clknet_leaf_236_clk),
    .D(booth_b4_m44),
    .Q(pp_row48_2));
 sky130_fd_sc_hd__dfxtp_1 _1767_ (.CLK(clknet_leaf_237_clk),
    .D(booth_b6_m42),
    .Q(pp_row48_3));
 sky130_fd_sc_hd__dfxtp_1 _1768_ (.CLK(clknet_leaf_238_clk),
    .D(booth_b8_m40),
    .Q(pp_row48_4));
 sky130_fd_sc_hd__dfxtp_1 _1769_ (.CLK(clknet_leaf_237_clk),
    .D(booth_b10_m38),
    .Q(pp_row48_5));
 sky130_fd_sc_hd__dfxtp_1 _1770_ (.CLK(clknet_leaf_238_clk),
    .D(booth_b12_m36),
    .Q(pp_row48_6));
 sky130_fd_sc_hd__dfxtp_1 _1771_ (.CLK(clknet_leaf_238_clk),
    .D(booth_b14_m34),
    .Q(pp_row48_7));
 sky130_fd_sc_hd__dfxtp_1 _1772_ (.CLK(clknet_leaf_187_clk),
    .D(booth_b64_m42),
    .Q(pp_row106_12));
 sky130_fd_sc_hd__dfxtp_1 _1773_ (.CLK(clknet_leaf_238_clk),
    .D(booth_b16_m32),
    .Q(pp_row48_8));
 sky130_fd_sc_hd__dfxtp_1 _1774_ (.CLK(clknet_leaf_238_clk),
    .D(booth_b18_m30),
    .Q(pp_row48_9));
 sky130_fd_sc_hd__dfxtp_1 _1775_ (.CLK(clknet_leaf_239_clk),
    .D(booth_b20_m28),
    .Q(pp_row48_10));
 sky130_fd_sc_hd__dfxtp_1 _1776_ (.CLK(clknet_leaf_238_clk),
    .D(booth_b22_m26),
    .Q(pp_row48_11));
 sky130_fd_sc_hd__dfxtp_1 _1777_ (.CLK(clknet_leaf_221_clk),
    .D(booth_b24_m24),
    .Q(pp_row48_12));
 sky130_fd_sc_hd__dfxtp_1 _1778_ (.CLK(clknet_leaf_220_clk),
    .D(booth_b26_m22),
    .Q(pp_row48_13));
 sky130_fd_sc_hd__dfxtp_1 _1779_ (.CLK(clknet_leaf_220_clk),
    .D(booth_b28_m20),
    .Q(pp_row48_14));
 sky130_fd_sc_hd__dfxtp_1 _1780_ (.CLK(clknet_leaf_222_clk),
    .D(booth_b30_m18),
    .Q(pp_row48_15));
 sky130_fd_sc_hd__dfxtp_1 _1781_ (.CLK(clknet_leaf_222_clk),
    .D(booth_b32_m16),
    .Q(pp_row48_16));
 sky130_fd_sc_hd__dfxtp_1 _1782_ (.CLK(clknet_leaf_222_clk),
    .D(booth_b34_m14),
    .Q(pp_row48_17));
 sky130_fd_sc_hd__dfxtp_1 _1783_ (.CLK(clknet_leaf_184_clk),
    .D(net136),
    .Q(pp_row106_13));
 sky130_fd_sc_hd__dfxtp_1 _1784_ (.CLK(clknet_leaf_222_clk),
    .D(booth_b36_m12),
    .Q(pp_row48_18));
 sky130_fd_sc_hd__dfxtp_1 _1785_ (.CLK(clknet_leaf_222_clk),
    .D(booth_b38_m10),
    .Q(pp_row48_19));
 sky130_fd_sc_hd__dfxtp_1 _1786_ (.CLK(clknet_leaf_222_clk),
    .D(booth_b40_m8),
    .Q(pp_row48_20));
 sky130_fd_sc_hd__dfxtp_1 _1787_ (.CLK(clknet_leaf_220_clk),
    .D(booth_b42_m6),
    .Q(pp_row48_21));
 sky130_fd_sc_hd__dfxtp_1 _1788_ (.CLK(clknet_leaf_220_clk),
    .D(booth_b44_m4),
    .Q(pp_row48_22));
 sky130_fd_sc_hd__dfxtp_1 _1789_ (.CLK(clknet_leaf_221_clk),
    .D(booth_b46_m2),
    .Q(pp_row48_23));
 sky130_fd_sc_hd__dfxtp_1 _1790_ (.CLK(clknet_leaf_221_clk),
    .D(booth_b48_m0),
    .Q(pp_row48_24));
 sky130_fd_sc_hd__dfxtp_1 _1791_ (.CLK(clknet_leaf_222_clk),
    .D(net1338),
    .Q(pp_row48_25));
 sky130_fd_sc_hd__dfxtp_1 _1792_ (.CLK(clknet_leaf_232_clk),
    .D(net199),
    .Q(pp_row48_26));
 sky130_fd_sc_hd__dfxtp_1 _1793_ (.CLK(clknet_leaf_35_clk),
    .D(booth_b0_m49),
    .Q(pp_row49_0));
 sky130_fd_sc_hd__dfxtp_1 _1794_ (.CLK(clknet_leaf_142_clk),
    .D(\notsign$5944 ),
    .Q(pp_row107_0));
 sky130_fd_sc_hd__dfxtp_1 _1795_ (.CLK(clknet_leaf_32_clk),
    .D(booth_b2_m47),
    .Q(pp_row49_1));
 sky130_fd_sc_hd__dfxtp_1 _1796_ (.CLK(clknet_leaf_37_clk),
    .D(booth_b4_m45),
    .Q(pp_row49_2));
 sky130_fd_sc_hd__dfxtp_1 _1797_ (.CLK(clknet_leaf_218_clk),
    .D(booth_b6_m43),
    .Q(pp_row49_3));
 sky130_fd_sc_hd__dfxtp_1 _1798_ (.CLK(clknet_leaf_219_clk),
    .D(booth_b8_m41),
    .Q(pp_row49_4));
 sky130_fd_sc_hd__dfxtp_1 _1799_ (.CLK(clknet_leaf_220_clk),
    .D(booth_b10_m39),
    .Q(pp_row49_5));
 sky130_fd_sc_hd__dfxtp_1 _1800_ (.CLK(clknet_leaf_220_clk),
    .D(booth_b12_m37),
    .Q(pp_row49_6));
 sky130_fd_sc_hd__dfxtp_1 _1801_ (.CLK(clknet_leaf_219_clk),
    .D(booth_b14_m35),
    .Q(pp_row49_7));
 sky130_fd_sc_hd__dfxtp_1 _1802_ (.CLK(clknet_leaf_219_clk),
    .D(booth_b16_m33),
    .Q(pp_row49_8));
 sky130_fd_sc_hd__dfxtp_1 _1803_ (.CLK(clknet_leaf_220_clk),
    .D(booth_b18_m31),
    .Q(pp_row49_9));
 sky130_fd_sc_hd__dfxtp_1 _1804_ (.CLK(clknet_leaf_220_clk),
    .D(booth_b20_m29),
    .Q(pp_row49_10));
 sky130_fd_sc_hd__dfxtp_1 _1805_ (.CLK(clknet_leaf_141_clk),
    .D(booth_b44_m63),
    .Q(pp_row107_1));
 sky130_fd_sc_hd__dfxtp_1 _1806_ (.CLK(clknet_leaf_220_clk),
    .D(booth_b22_m27),
    .Q(pp_row49_11));
 sky130_fd_sc_hd__dfxtp_1 _1807_ (.CLK(clknet_leaf_24_clk),
    .D(booth_b24_m25),
    .Q(pp_row49_12));
 sky130_fd_sc_hd__dfxtp_1 _1808_ (.CLK(clknet_leaf_24_clk),
    .D(booth_b26_m23),
    .Q(pp_row49_13));
 sky130_fd_sc_hd__dfxtp_1 _1809_ (.CLK(clknet_leaf_24_clk),
    .D(booth_b28_m21),
    .Q(pp_row49_14));
 sky130_fd_sc_hd__dfxtp_1 _1810_ (.CLK(clknet_leaf_26_clk),
    .D(booth_b30_m19),
    .Q(pp_row49_15));
 sky130_fd_sc_hd__dfxtp_1 _1811_ (.CLK(clknet_leaf_26_clk),
    .D(booth_b32_m17),
    .Q(pp_row49_16));
 sky130_fd_sc_hd__dfxtp_1 _1812_ (.CLK(clknet_leaf_26_clk),
    .D(booth_b34_m15),
    .Q(pp_row49_17));
 sky130_fd_sc_hd__dfxtp_1 _1813_ (.CLK(clknet_leaf_25_clk),
    .D(booth_b36_m13),
    .Q(pp_row49_18));
 sky130_fd_sc_hd__dfxtp_1 _1814_ (.CLK(clknet_leaf_26_clk),
    .D(booth_b38_m11),
    .Q(pp_row49_19));
 sky130_fd_sc_hd__dfxtp_1 _1815_ (.CLK(clknet_leaf_25_clk),
    .D(booth_b40_m9),
    .Q(pp_row49_20));
 sky130_fd_sc_hd__dfxtp_1 _1816_ (.CLK(clknet_leaf_141_clk),
    .D(booth_b46_m61),
    .Q(pp_row107_2));
 sky130_fd_sc_hd__dfxtp_1 _1817_ (.CLK(clknet_leaf_224_clk),
    .D(booth_b42_m7),
    .Q(pp_row49_21));
 sky130_fd_sc_hd__dfxtp_1 _1818_ (.CLK(clknet_leaf_222_clk),
    .D(booth_b44_m5),
    .Q(pp_row49_22));
 sky130_fd_sc_hd__dfxtp_1 _1819_ (.CLK(clknet_leaf_220_clk),
    .D(booth_b46_m3),
    .Q(pp_row49_23));
 sky130_fd_sc_hd__dfxtp_1 _1820_ (.CLK(clknet_leaf_220_clk),
    .D(booth_b48_m1),
    .Q(pp_row49_24));
 sky130_fd_sc_hd__dfxtp_1 _1821_ (.CLK(clknet_leaf_235_clk),
    .D(net200),
    .Q(pp_row49_25));
 sky130_fd_sc_hd__dfxtp_1 _1822_ (.CLK(clknet_leaf_232_clk),
    .D(booth_b0_m50),
    .Q(pp_row50_0));
 sky130_fd_sc_hd__dfxtp_1 _1823_ (.CLK(clknet_leaf_234_clk),
    .D(booth_b2_m48),
    .Q(pp_row50_1));
 sky130_fd_sc_hd__dfxtp_1 _1824_ (.CLK(clknet_leaf_234_clk),
    .D(booth_b4_m46),
    .Q(pp_row50_2));
 sky130_fd_sc_hd__dfxtp_1 _1825_ (.CLK(clknet_leaf_234_clk),
    .D(booth_b6_m44),
    .Q(pp_row50_3));
 sky130_fd_sc_hd__dfxtp_1 _1826_ (.CLK(clknet_leaf_234_clk),
    .D(booth_b8_m42),
    .Q(pp_row50_4));
 sky130_fd_sc_hd__dfxtp_1 _1827_ (.CLK(clknet_leaf_135_clk),
    .D(booth_b48_m59),
    .Q(pp_row107_3));
 sky130_fd_sc_hd__dfxtp_1 _1828_ (.CLK(clknet_leaf_234_clk),
    .D(booth_b10_m40),
    .Q(pp_row50_5));
 sky130_fd_sc_hd__dfxtp_1 _1829_ (.CLK(clknet_leaf_34_clk),
    .D(booth_b12_m38),
    .Q(pp_row50_6));
 sky130_fd_sc_hd__dfxtp_1 _1830_ (.CLK(clknet_leaf_34_clk),
    .D(booth_b14_m36),
    .Q(pp_row50_7));
 sky130_fd_sc_hd__dfxtp_1 _1831_ (.CLK(clknet_leaf_25_clk),
    .D(booth_b16_m34),
    .Q(pp_row50_8));
 sky130_fd_sc_hd__dfxtp_1 _1832_ (.CLK(clknet_leaf_18_clk),
    .D(booth_b18_m32),
    .Q(pp_row50_9));
 sky130_fd_sc_hd__dfxtp_1 _1833_ (.CLK(clknet_leaf_18_clk),
    .D(booth_b20_m30),
    .Q(pp_row50_10));
 sky130_fd_sc_hd__dfxtp_1 _1834_ (.CLK(clknet_leaf_18_clk),
    .D(booth_b22_m28),
    .Q(pp_row50_11));
 sky130_fd_sc_hd__dfxtp_1 _1835_ (.CLK(clknet_leaf_25_clk),
    .D(booth_b24_m26),
    .Q(pp_row50_12));
 sky130_fd_sc_hd__dfxtp_1 _1836_ (.CLK(clknet_leaf_25_clk),
    .D(booth_b26_m24),
    .Q(pp_row50_13));
 sky130_fd_sc_hd__dfxtp_1 _1837_ (.CLK(clknet_leaf_25_clk),
    .D(booth_b28_m22),
    .Q(pp_row50_14));
 sky130_fd_sc_hd__dfxtp_1 _1838_ (.CLK(clknet_leaf_135_clk),
    .D(booth_b50_m57),
    .Q(pp_row107_4));
 sky130_fd_sc_hd__dfxtp_2 _1839_ (.CLK(clknet_leaf_181_clk),
    .D(net155),
    .Q(pp_row123_4));
 sky130_fd_sc_hd__dfxtp_1 _1840_ (.CLK(clknet_leaf_62_clk),
    .D(booth_b30_m20),
    .Q(pp_row50_15));
 sky130_fd_sc_hd__dfxtp_1 _1841_ (.CLK(clknet_leaf_62_clk),
    .D(booth_b32_m18),
    .Q(pp_row50_16));
 sky130_fd_sc_hd__dfxtp_1 _1842_ (.CLK(clknet_leaf_62_clk),
    .D(booth_b34_m16),
    .Q(pp_row50_17));
 sky130_fd_sc_hd__dfxtp_1 _1843_ (.CLK(clknet_leaf_71_clk),
    .D(booth_b36_m14),
    .Q(pp_row50_18));
 sky130_fd_sc_hd__dfxtp_1 _1844_ (.CLK(clknet_leaf_71_clk),
    .D(booth_b38_m12),
    .Q(pp_row50_19));
 sky130_fd_sc_hd__dfxtp_1 _1845_ (.CLK(clknet_leaf_71_clk),
    .D(booth_b40_m10),
    .Q(pp_row50_20));
 sky130_fd_sc_hd__dfxtp_1 _1846_ (.CLK(clknet_leaf_71_clk),
    .D(booth_b42_m8),
    .Q(pp_row50_21));
 sky130_fd_sc_hd__dfxtp_1 _1847_ (.CLK(clknet_leaf_70_clk),
    .D(booth_b44_m6),
    .Q(pp_row50_22));
 sky130_fd_sc_hd__dfxtp_1 _1848_ (.CLK(clknet_leaf_73_clk),
    .D(booth_b46_m4),
    .Q(pp_row50_23));
 sky130_fd_sc_hd__dfxtp_1 _1849_ (.CLK(clknet_leaf_25_clk),
    .D(booth_b48_m2),
    .Q(pp_row50_24));
 sky130_fd_sc_hd__dfxtp_1 _1850_ (.CLK(clknet_leaf_135_clk),
    .D(booth_b52_m55),
    .Q(pp_row107_5));
 sky130_fd_sc_hd__dfxtp_1 _1851_ (.CLK(clknet_leaf_25_clk),
    .D(booth_b50_m0),
    .Q(pp_row50_25));
 sky130_fd_sc_hd__dfxtp_1 _1852_ (.CLK(clknet_leaf_25_clk),
    .D(net1332),
    .Q(pp_row50_26));
 sky130_fd_sc_hd__dfxtp_2 _1853_ (.CLK(clknet_leaf_232_clk),
    .D(net202),
    .Q(pp_row50_27));
 sky130_fd_sc_hd__dfxtp_1 _1854_ (.CLK(clknet_leaf_67_clk),
    .D(booth_b0_m51),
    .Q(pp_row51_0));
 sky130_fd_sc_hd__dfxtp_1 _1855_ (.CLK(clknet_leaf_68_clk),
    .D(booth_b2_m49),
    .Q(pp_row51_1));
 sky130_fd_sc_hd__dfxtp_1 _1856_ (.CLK(clknet_leaf_67_clk),
    .D(booth_b4_m47),
    .Q(pp_row51_2));
 sky130_fd_sc_hd__dfxtp_1 _1857_ (.CLK(clknet_leaf_79_clk),
    .D(booth_b6_m45),
    .Q(pp_row51_3));
 sky130_fd_sc_hd__dfxtp_1 _1858_ (.CLK(clknet_leaf_78_clk),
    .D(booth_b8_m43),
    .Q(pp_row51_4));
 sky130_fd_sc_hd__dfxtp_1 _1859_ (.CLK(clknet_leaf_79_clk),
    .D(booth_b10_m41),
    .Q(pp_row51_5));
 sky130_fd_sc_hd__dfxtp_1 _1860_ (.CLK(clknet_leaf_80_clk),
    .D(booth_b12_m39),
    .Q(pp_row51_6));
 sky130_fd_sc_hd__dfxtp_1 _1861_ (.CLK(clknet_leaf_133_clk),
    .D(booth_b54_m53),
    .Q(pp_row107_6));
 sky130_fd_sc_hd__dfxtp_1 _1862_ (.CLK(clknet_leaf_66_clk),
    .D(booth_b14_m37),
    .Q(pp_row51_7));
 sky130_fd_sc_hd__dfxtp_1 _1863_ (.CLK(clknet_leaf_66_clk),
    .D(booth_b16_m35),
    .Q(pp_row51_8));
 sky130_fd_sc_hd__dfxtp_1 _1864_ (.CLK(clknet_leaf_67_clk),
    .D(booth_b18_m33),
    .Q(pp_row51_9));
 sky130_fd_sc_hd__dfxtp_1 _1865_ (.CLK(clknet_leaf_66_clk),
    .D(booth_b20_m31),
    .Q(pp_row51_10));
 sky130_fd_sc_hd__dfxtp_1 _1866_ (.CLK(clknet_leaf_67_clk),
    .D(booth_b22_m29),
    .Q(pp_row51_11));
 sky130_fd_sc_hd__dfxtp_1 _1867_ (.CLK(clknet_leaf_66_clk),
    .D(booth_b24_m27),
    .Q(pp_row51_12));
 sky130_fd_sc_hd__dfxtp_1 _1868_ (.CLK(clknet_leaf_66_clk),
    .D(booth_b26_m25),
    .Q(pp_row51_13));
 sky130_fd_sc_hd__dfxtp_1 _1869_ (.CLK(clknet_leaf_66_clk),
    .D(booth_b28_m23),
    .Q(pp_row51_14));
 sky130_fd_sc_hd__dfxtp_1 _1870_ (.CLK(clknet_leaf_68_clk),
    .D(booth_b30_m21),
    .Q(pp_row51_15));
 sky130_fd_sc_hd__dfxtp_1 _1871_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b32_m19),
    .Q(pp_row51_16));
 sky130_fd_sc_hd__dfxtp_1 _1872_ (.CLK(clknet_leaf_134_clk),
    .D(booth_b56_m51),
    .Q(pp_row107_7));
 sky130_fd_sc_hd__dfxtp_1 _1873_ (.CLK(clknet_leaf_71_clk),
    .D(booth_b34_m17),
    .Q(pp_row51_17));
 sky130_fd_sc_hd__dfxtp_1 _1874_ (.CLK(clknet_leaf_69_clk),
    .D(booth_b36_m15),
    .Q(pp_row51_18));
 sky130_fd_sc_hd__dfxtp_1 _1875_ (.CLK(clknet_leaf_69_clk),
    .D(booth_b38_m13),
    .Q(pp_row51_19));
 sky130_fd_sc_hd__dfxtp_1 _1876_ (.CLK(clknet_leaf_69_clk),
    .D(booth_b40_m11),
    .Q(pp_row51_20));
 sky130_fd_sc_hd__dfxtp_1 _1877_ (.CLK(clknet_leaf_70_clk),
    .D(booth_b42_m9),
    .Q(pp_row51_21));
 sky130_fd_sc_hd__dfxtp_1 _1878_ (.CLK(clknet_leaf_70_clk),
    .D(booth_b44_m7),
    .Q(pp_row51_22));
 sky130_fd_sc_hd__dfxtp_1 _1879_ (.CLK(clknet_leaf_70_clk),
    .D(booth_b46_m5),
    .Q(pp_row51_23));
 sky130_fd_sc_hd__dfxtp_1 _1880_ (.CLK(clknet_leaf_27_clk),
    .D(booth_b48_m3),
    .Q(pp_row51_24));
 sky130_fd_sc_hd__dfxtp_1 _1881_ (.CLK(clknet_leaf_25_clk),
    .D(booth_b50_m1),
    .Q(pp_row51_25));
 sky130_fd_sc_hd__dfxtp_1 _1882_ (.CLK(clknet_leaf_232_clk),
    .D(net203),
    .Q(pp_row51_26));
 sky130_fd_sc_hd__dfxtp_1 _1883_ (.CLK(clknet_leaf_134_clk),
    .D(booth_b58_m49),
    .Q(pp_row107_8));
 sky130_fd_sc_hd__dfxtp_1 _1884_ (.CLK(clknet_leaf_78_clk),
    .D(booth_b0_m52),
    .Q(pp_row52_0));
 sky130_fd_sc_hd__dfxtp_1 _1885_ (.CLK(clknet_leaf_78_clk),
    .D(booth_b2_m50),
    .Q(pp_row52_1));
 sky130_fd_sc_hd__dfxtp_1 _1886_ (.CLK(clknet_leaf_80_clk),
    .D(booth_b4_m48),
    .Q(pp_row52_2));
 sky130_fd_sc_hd__dfxtp_1 _1887_ (.CLK(clknet_leaf_80_clk),
    .D(booth_b6_m46),
    .Q(pp_row52_3));
 sky130_fd_sc_hd__dfxtp_1 _1888_ (.CLK(clknet_leaf_39_clk),
    .D(booth_b8_m44),
    .Q(pp_row52_4));
 sky130_fd_sc_hd__dfxtp_1 _1889_ (.CLK(clknet_leaf_39_clk),
    .D(booth_b10_m42),
    .Q(pp_row52_5));
 sky130_fd_sc_hd__dfxtp_1 _1890_ (.CLK(clknet_leaf_39_clk),
    .D(booth_b12_m40),
    .Q(pp_row52_6));
 sky130_fd_sc_hd__dfxtp_1 _1891_ (.CLK(clknet_leaf_39_clk),
    .D(booth_b14_m38),
    .Q(pp_row52_7));
 sky130_fd_sc_hd__dfxtp_1 _1892_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b16_m36),
    .Q(pp_row52_8));
 sky130_fd_sc_hd__dfxtp_1 _1893_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b18_m34),
    .Q(pp_row52_9));
 sky130_fd_sc_hd__dfxtp_1 _1894_ (.CLK(clknet_leaf_137_clk),
    .D(booth_b60_m47),
    .Q(pp_row107_9));
 sky130_fd_sc_hd__dfxtp_1 _1895_ (.CLK(clknet_leaf_65_clk),
    .D(booth_b20_m32),
    .Q(pp_row52_10));
 sky130_fd_sc_hd__dfxtp_1 _1896_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b22_m30),
    .Q(pp_row52_11));
 sky130_fd_sc_hd__dfxtp_1 _1897_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b24_m28),
    .Q(pp_row52_12));
 sky130_fd_sc_hd__dfxtp_1 _1898_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b26_m26),
    .Q(pp_row52_13));
 sky130_fd_sc_hd__dfxtp_1 _1899_ (.CLK(clknet_leaf_63_clk),
    .D(booth_b28_m24),
    .Q(pp_row52_14));
 sky130_fd_sc_hd__dfxtp_1 _1900_ (.CLK(clknet_leaf_63_clk),
    .D(booth_b30_m22),
    .Q(pp_row52_15));
 sky130_fd_sc_hd__dfxtp_1 _1901_ (.CLK(clknet_leaf_63_clk),
    .D(booth_b32_m20),
    .Q(pp_row52_16));
 sky130_fd_sc_hd__dfxtp_1 _1902_ (.CLK(clknet_leaf_71_clk),
    .D(booth_b34_m18),
    .Q(pp_row52_17));
 sky130_fd_sc_hd__dfxtp_1 _1903_ (.CLK(clknet_leaf_71_clk),
    .D(booth_b36_m16),
    .Q(pp_row52_18));
 sky130_fd_sc_hd__dfxtp_1 _1904_ (.CLK(clknet_leaf_71_clk),
    .D(booth_b38_m14),
    .Q(pp_row52_19));
 sky130_fd_sc_hd__dfxtp_1 _1905_ (.CLK(clknet_leaf_138_clk),
    .D(booth_b62_m45),
    .Q(pp_row107_10));
 sky130_fd_sc_hd__dfxtp_1 _1906_ (.CLK(clknet_leaf_70_clk),
    .D(booth_b40_m12),
    .Q(pp_row52_20));
 sky130_fd_sc_hd__dfxtp_1 _1907_ (.CLK(clknet_leaf_70_clk),
    .D(booth_b42_m10),
    .Q(pp_row52_21));
 sky130_fd_sc_hd__dfxtp_1 _1908_ (.CLK(clknet_leaf_70_clk),
    .D(booth_b44_m8),
    .Q(pp_row52_22));
 sky130_fd_sc_hd__dfxtp_1 _1909_ (.CLK(clknet_leaf_70_clk),
    .D(booth_b46_m6),
    .Q(pp_row52_23));
 sky130_fd_sc_hd__dfxtp_1 _1910_ (.CLK(clknet_leaf_70_clk),
    .D(booth_b48_m4),
    .Q(pp_row52_24));
 sky130_fd_sc_hd__dfxtp_1 _1911_ (.CLK(clknet_leaf_70_clk),
    .D(booth_b50_m2),
    .Q(pp_row52_25));
 sky130_fd_sc_hd__dfxtp_1 _1912_ (.CLK(clknet_leaf_31_clk),
    .D(booth_b52_m0),
    .Q(pp_row52_26));
 sky130_fd_sc_hd__dfxtp_1 _1913_ (.CLK(clknet_leaf_31_clk),
    .D(net1320),
    .Q(pp_row52_27));
 sky130_fd_sc_hd__dfxtp_2 _1914_ (.CLK(clknet_leaf_232_clk),
    .D(net204),
    .Q(pp_row52_28));
 sky130_fd_sc_hd__dfxtp_1 _1915_ (.CLK(clknet_leaf_67_clk),
    .D(booth_b0_m53),
    .Q(pp_row53_0));
 sky130_fd_sc_hd__dfxtp_1 _1916_ (.CLK(clknet_leaf_138_clk),
    .D(booth_b64_m43),
    .Q(pp_row107_11));
 sky130_fd_sc_hd__dfxtp_1 _1917_ (.CLK(clknet_leaf_68_clk),
    .D(booth_b2_m51),
    .Q(pp_row53_1));
 sky130_fd_sc_hd__dfxtp_1 _1918_ (.CLK(clknet_leaf_81_clk),
    .D(booth_b4_m49),
    .Q(pp_row53_2));
 sky130_fd_sc_hd__dfxtp_1 _1919_ (.CLK(clknet_leaf_80_clk),
    .D(booth_b6_m47),
    .Q(pp_row53_3));
 sky130_fd_sc_hd__dfxtp_1 _1920_ (.CLK(clknet_leaf_81_clk),
    .D(booth_b8_m45),
    .Q(pp_row53_4));
 sky130_fd_sc_hd__dfxtp_1 _1921_ (.CLK(clknet_leaf_80_clk),
    .D(booth_b10_m43),
    .Q(pp_row53_5));
 sky130_fd_sc_hd__dfxtp_1 _1922_ (.CLK(clknet_leaf_80_clk),
    .D(booth_b12_m41),
    .Q(pp_row53_6));
 sky130_fd_sc_hd__dfxtp_1 _1923_ (.CLK(clknet_leaf_80_clk),
    .D(booth_b14_m39),
    .Q(pp_row53_7));
 sky130_fd_sc_hd__dfxtp_1 _1924_ (.CLK(clknet_leaf_65_clk),
    .D(booth_b16_m37),
    .Q(pp_row53_8));
 sky130_fd_sc_hd__dfxtp_1 _1925_ (.CLK(clknet_leaf_65_clk),
    .D(booth_b18_m35),
    .Q(pp_row53_9));
 sky130_fd_sc_hd__dfxtp_1 _1926_ (.CLK(clknet_leaf_65_clk),
    .D(booth_b20_m33),
    .Q(pp_row53_10));
 sky130_fd_sc_hd__dfxtp_2 _1927_ (.CLK(clknet_leaf_184_clk),
    .D(net137),
    .Q(pp_row107_12));
 sky130_fd_sc_hd__dfxtp_1 _1928_ (.CLK(clknet_leaf_69_clk),
    .D(booth_b22_m31),
    .Q(pp_row53_11));
 sky130_fd_sc_hd__dfxtp_1 _1929_ (.CLK(clknet_leaf_67_clk),
    .D(booth_b24_m29),
    .Q(pp_row53_12));
 sky130_fd_sc_hd__dfxtp_1 _1930_ (.CLK(clknet_leaf_62_clk),
    .D(booth_b26_m27),
    .Q(pp_row53_13));
 sky130_fd_sc_hd__dfxtp_1 _1931_ (.CLK(clknet_leaf_62_clk),
    .D(booth_b28_m25),
    .Q(pp_row53_14));
 sky130_fd_sc_hd__dfxtp_1 _1932_ (.CLK(clknet_leaf_62_clk),
    .D(booth_b30_m23),
    .Q(pp_row53_15));
 sky130_fd_sc_hd__dfxtp_1 _1933_ (.CLK(clknet_leaf_62_clk),
    .D(booth_b32_m21),
    .Q(pp_row53_16));
 sky130_fd_sc_hd__dfxtp_1 _1934_ (.CLK(clknet_leaf_69_clk),
    .D(booth_b34_m19),
    .Q(pp_row53_17));
 sky130_fd_sc_hd__dfxtp_1 _1935_ (.CLK(clknet_leaf_70_clk),
    .D(booth_b36_m17),
    .Q(pp_row53_18));
 sky130_fd_sc_hd__dfxtp_1 _1936_ (.CLK(clknet_leaf_70_clk),
    .D(booth_b38_m15),
    .Q(pp_row53_19));
 sky130_fd_sc_hd__dfxtp_1 _1937_ (.CLK(clknet_leaf_70_clk),
    .D(booth_b40_m13),
    .Q(pp_row53_20));
 sky130_fd_sc_hd__dfxtp_1 _1938_ (.CLK(clknet_leaf_136_clk),
    .D(booth_b44_m64),
    .Q(pp_row108_1));
 sky130_fd_sc_hd__dfxtp_1 _1939_ (.CLK(clknet_leaf_70_clk),
    .D(booth_b42_m11),
    .Q(pp_row53_21));
 sky130_fd_sc_hd__dfxtp_1 _1940_ (.CLK(clknet_leaf_70_clk),
    .D(booth_b44_m9),
    .Q(pp_row53_22));
 sky130_fd_sc_hd__dfxtp_1 _1941_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b46_m7),
    .Q(pp_row53_23));
 sky130_fd_sc_hd__dfxtp_1 _1942_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b48_m5),
    .Q(pp_row53_24));
 sky130_fd_sc_hd__dfxtp_1 _1943_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b50_m3),
    .Q(pp_row53_25));
 sky130_fd_sc_hd__dfxtp_1 _1944_ (.CLK(clknet_leaf_78_clk),
    .D(booth_b52_m1),
    .Q(pp_row53_26));
 sky130_fd_sc_hd__dfxtp_4 _1945_ (.CLK(clknet_leaf_231_clk),
    .D(net205),
    .Q(pp_row53_27));
 sky130_fd_sc_hd__dfxtp_1 _1946_ (.CLK(clknet_leaf_78_clk),
    .D(booth_b0_m54),
    .Q(pp_row54_0));
 sky130_fd_sc_hd__dfxtp_1 _1947_ (.CLK(clknet_leaf_78_clk),
    .D(booth_b2_m52),
    .Q(pp_row54_1));
 sky130_fd_sc_hd__dfxtp_1 _1948_ (.CLK(clknet_leaf_78_clk),
    .D(booth_b4_m50),
    .Q(pp_row54_2));
 sky130_fd_sc_hd__dfxtp_1 _1949_ (.CLK(clknet_leaf_137_clk),
    .D(booth_b46_m62),
    .Q(pp_row108_2));
 sky130_fd_sc_hd__dfxtp_1 _1950_ (.CLK(clknet_leaf_164_clk),
    .D(booth_b60_m64),
    .Q(pp_row124_1));
 sky130_fd_sc_hd__dfxtp_1 _1951_ (.CLK(clknet_leaf_66_clk),
    .D(booth_b6_m48),
    .Q(pp_row54_3));
 sky130_fd_sc_hd__dfxtp_1 _1952_ (.CLK(clknet_leaf_66_clk),
    .D(booth_b8_m46),
    .Q(pp_row54_4));
 sky130_fd_sc_hd__dfxtp_1 _1953_ (.CLK(clknet_leaf_66_clk),
    .D(booth_b10_m44),
    .Q(pp_row54_5));
 sky130_fd_sc_hd__dfxtp_1 _1954_ (.CLK(clknet_leaf_66_clk),
    .D(booth_b12_m42),
    .Q(pp_row54_6));
 sky130_fd_sc_hd__dfxtp_1 _1955_ (.CLK(clknet_leaf_66_clk),
    .D(booth_b14_m40),
    .Q(pp_row54_7));
 sky130_fd_sc_hd__dfxtp_1 _1956_ (.CLK(clknet_leaf_66_clk),
    .D(booth_b16_m38),
    .Q(pp_row54_8));
 sky130_fd_sc_hd__dfxtp_1 _1957_ (.CLK(clknet_leaf_66_clk),
    .D(booth_b18_m36),
    .Q(pp_row54_9));
 sky130_fd_sc_hd__dfxtp_1 _1958_ (.CLK(clknet_leaf_66_clk),
    .D(booth_b20_m34),
    .Q(pp_row54_10));
 sky130_fd_sc_hd__dfxtp_1 _1959_ (.CLK(clknet_leaf_63_clk),
    .D(booth_b22_m32),
    .Q(pp_row54_11));
 sky130_fd_sc_hd__dfxtp_1 _1960_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b24_m30),
    .Q(pp_row54_12));
 sky130_fd_sc_hd__dfxtp_1 _1961_ (.CLK(clknet_leaf_138_clk),
    .D(booth_b48_m60),
    .Q(pp_row108_3));
 sky130_fd_sc_hd__dfxtp_1 _1962_ (.CLK(clknet_leaf_64_clk),
    .D(booth_b26_m28),
    .Q(pp_row54_13));
 sky130_fd_sc_hd__dfxtp_1 _1963_ (.CLK(clknet_leaf_63_clk),
    .D(booth_b28_m26),
    .Q(pp_row54_14));
 sky130_fd_sc_hd__dfxtp_1 _1964_ (.CLK(clknet_leaf_63_clk),
    .D(booth_b30_m24),
    .Q(pp_row54_15));
 sky130_fd_sc_hd__dfxtp_1 _1965_ (.CLK(clknet_leaf_62_clk),
    .D(booth_b32_m22),
    .Q(pp_row54_16));
 sky130_fd_sc_hd__dfxtp_1 _1966_ (.CLK(clknet_leaf_63_clk),
    .D(booth_b34_m20),
    .Q(pp_row54_17));
 sky130_fd_sc_hd__dfxtp_1 _1967_ (.CLK(clknet_leaf_63_clk),
    .D(booth_b36_m18),
    .Q(pp_row54_18));
 sky130_fd_sc_hd__dfxtp_1 _1968_ (.CLK(clknet_leaf_62_clk),
    .D(booth_b38_m16),
    .Q(pp_row54_19));
 sky130_fd_sc_hd__dfxtp_1 _1969_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b40_m14),
    .Q(pp_row54_20));
 sky130_fd_sc_hd__dfxtp_1 _1970_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b42_m12),
    .Q(pp_row54_21));
 sky130_fd_sc_hd__dfxtp_1 _1971_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b44_m10),
    .Q(pp_row54_22));
 sky130_fd_sc_hd__dfxtp_1 _1972_ (.CLK(clknet_leaf_138_clk),
    .D(booth_b50_m58),
    .Q(pp_row108_4));
 sky130_fd_sc_hd__dfxtp_1 _1973_ (.CLK(clknet_leaf_71_clk),
    .D(booth_b46_m8),
    .Q(pp_row54_23));
 sky130_fd_sc_hd__dfxtp_1 _1974_ (.CLK(clknet_leaf_71_clk),
    .D(booth_b48_m6),
    .Q(pp_row54_24));
 sky130_fd_sc_hd__dfxtp_1 _1975_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b50_m4),
    .Q(pp_row54_25));
 sky130_fd_sc_hd__dfxtp_1 _1976_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b52_m2),
    .Q(pp_row54_26));
 sky130_fd_sc_hd__dfxtp_1 _1977_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b54_m0),
    .Q(pp_row54_27));
 sky130_fd_sc_hd__dfxtp_1 _1978_ (.CLK(clknet_leaf_72_clk),
    .D(net1304),
    .Q(pp_row54_28));
 sky130_fd_sc_hd__dfxtp_4 _1979_ (.CLK(clknet_leaf_235_clk),
    .D(net206),
    .Q(pp_row54_29));
 sky130_fd_sc_hd__dfxtp_1 _1980_ (.CLK(clknet_leaf_78_clk),
    .D(booth_b0_m55),
    .Q(pp_row55_0));
 sky130_fd_sc_hd__dfxtp_1 _1981_ (.CLK(clknet_leaf_78_clk),
    .D(booth_b2_m53),
    .Q(pp_row55_1));
 sky130_fd_sc_hd__dfxtp_1 _1982_ (.CLK(clknet_leaf_78_clk),
    .D(booth_b4_m51),
    .Q(pp_row55_2));
 sky130_fd_sc_hd__dfxtp_1 _1983_ (.CLK(clknet_leaf_136_clk),
    .D(booth_b52_m56),
    .Q(pp_row108_5));
 sky130_fd_sc_hd__dfxtp_1 _1984_ (.CLK(clknet_leaf_79_clk),
    .D(booth_b6_m49),
    .Q(pp_row55_3));
 sky130_fd_sc_hd__dfxtp_1 _1985_ (.CLK(clknet_leaf_79_clk),
    .D(booth_b8_m47),
    .Q(pp_row55_4));
 sky130_fd_sc_hd__dfxtp_1 _1986_ (.CLK(clknet_leaf_81_clk),
    .D(booth_b10_m45),
    .Q(pp_row55_5));
 sky130_fd_sc_hd__dfxtp_1 _1987_ (.CLK(clknet_leaf_81_clk),
    .D(booth_b12_m43),
    .Q(pp_row55_6));
 sky130_fd_sc_hd__dfxtp_1 _1988_ (.CLK(clknet_leaf_38_clk),
    .D(booth_b14_m41),
    .Q(pp_row55_7));
 sky130_fd_sc_hd__dfxtp_1 _1989_ (.CLK(clknet_leaf_81_clk),
    .D(booth_b16_m39),
    .Q(pp_row55_8));
 sky130_fd_sc_hd__dfxtp_1 _1990_ (.CLK(clknet_leaf_81_clk),
    .D(booth_b18_m37),
    .Q(pp_row55_9));
 sky130_fd_sc_hd__dfxtp_1 _1991_ (.CLK(clknet_leaf_81_clk),
    .D(booth_b20_m35),
    .Q(pp_row55_10));
 sky130_fd_sc_hd__dfxtp_1 _1992_ (.CLK(clknet_leaf_69_clk),
    .D(booth_b22_m33),
    .Q(pp_row55_11));
 sky130_fd_sc_hd__dfxtp_1 _1993_ (.CLK(clknet_leaf_67_clk),
    .D(booth_b24_m31),
    .Q(pp_row55_12));
 sky130_fd_sc_hd__dfxtp_1 _1994_ (.CLK(clknet_leaf_143_clk),
    .D(booth_b54_m54),
    .Q(pp_row108_6));
 sky130_fd_sc_hd__dfxtp_1 _1995_ (.CLK(clknet_leaf_67_clk),
    .D(booth_b26_m29),
    .Q(pp_row55_13));
 sky130_fd_sc_hd__dfxtp_1 _1996_ (.CLK(clknet_leaf_69_clk),
    .D(booth_b28_m27),
    .Q(pp_row55_14));
 sky130_fd_sc_hd__dfxtp_1 _1997_ (.CLK(clknet_leaf_69_clk),
    .D(booth_b30_m25),
    .Q(pp_row55_15));
 sky130_fd_sc_hd__dfxtp_1 _1998_ (.CLK(clknet_leaf_69_clk),
    .D(booth_b32_m23),
    .Q(pp_row55_16));
 sky130_fd_sc_hd__dfxtp_1 _1999_ (.CLK(clknet_leaf_62_clk),
    .D(booth_b34_m21),
    .Q(pp_row55_17));
 sky130_fd_sc_hd__dfxtp_1 _2000_ (.CLK(clknet_leaf_69_clk),
    .D(booth_b36_m19),
    .Q(pp_row55_18));
 sky130_fd_sc_hd__dfxtp_1 _2001_ (.CLK(clknet_leaf_62_clk),
    .D(booth_b38_m17),
    .Q(pp_row55_19));
 sky130_fd_sc_hd__dfxtp_1 _2002_ (.CLK(clknet_leaf_73_clk),
    .D(booth_b40_m15),
    .Q(pp_row55_20));
 sky130_fd_sc_hd__dfxtp_1 _2003_ (.CLK(clknet_leaf_73_clk),
    .D(booth_b42_m13),
    .Q(pp_row55_21));
 sky130_fd_sc_hd__dfxtp_1 _2004_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b44_m11),
    .Q(pp_row55_22));
 sky130_fd_sc_hd__dfxtp_1 _2005_ (.CLK(clknet_leaf_142_clk),
    .D(booth_b56_m52),
    .Q(pp_row108_7));
 sky130_fd_sc_hd__dfxtp_1 _2006_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b46_m9),
    .Q(pp_row55_23));
 sky130_fd_sc_hd__dfxtp_1 _2007_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b48_m7),
    .Q(pp_row55_24));
 sky130_fd_sc_hd__dfxtp_1 _2008_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b50_m5),
    .Q(pp_row55_25));
 sky130_fd_sc_hd__dfxtp_1 _2009_ (.CLK(clknet_leaf_76_clk),
    .D(booth_b52_m3),
    .Q(pp_row55_26));
 sky130_fd_sc_hd__dfxtp_1 _2010_ (.CLK(clknet_leaf_75_clk),
    .D(booth_b54_m1),
    .Q(pp_row55_27));
 sky130_fd_sc_hd__dfxtp_4 _2011_ (.CLK(clknet_leaf_231_clk),
    .D(net207),
    .Q(pp_row55_28));
 sky130_fd_sc_hd__dfxtp_1 _2012_ (.CLK(clknet_leaf_83_clk),
    .D(booth_b0_m56),
    .Q(pp_row56_0));
 sky130_fd_sc_hd__dfxtp_1 _2013_ (.CLK(clknet_leaf_83_clk),
    .D(booth_b2_m54),
    .Q(pp_row56_1));
 sky130_fd_sc_hd__dfxtp_1 _2014_ (.CLK(clknet_leaf_81_clk),
    .D(booth_b4_m52),
    .Q(pp_row56_2));
 sky130_fd_sc_hd__dfxtp_1 _2015_ (.CLK(clknet_leaf_81_clk),
    .D(booth_b6_m50),
    .Q(pp_row56_3));
 sky130_fd_sc_hd__dfxtp_1 _2016_ (.CLK(clknet_leaf_135_clk),
    .D(booth_b58_m50),
    .Q(pp_row108_8));
 sky130_fd_sc_hd__dfxtp_1 _2017_ (.CLK(clknet_leaf_81_clk),
    .D(booth_b8_m48),
    .Q(pp_row56_4));
 sky130_fd_sc_hd__dfxtp_1 _2018_ (.CLK(clknet_leaf_81_clk),
    .D(booth_b10_m46),
    .Q(pp_row56_5));
 sky130_fd_sc_hd__dfxtp_1 _2019_ (.CLK(clknet_leaf_81_clk),
    .D(booth_b12_m44),
    .Q(pp_row56_6));
 sky130_fd_sc_hd__dfxtp_1 _2020_ (.CLK(clknet_leaf_38_clk),
    .D(booth_b14_m42),
    .Q(pp_row56_7));
 sky130_fd_sc_hd__dfxtp_1 _2021_ (.CLK(clknet_leaf_33_clk),
    .D(booth_b16_m40),
    .Q(pp_row56_8));
 sky130_fd_sc_hd__dfxtp_1 _2022_ (.CLK(clknet_leaf_34_clk),
    .D(booth_b18_m38),
    .Q(pp_row56_9));
 sky130_fd_sc_hd__dfxtp_1 _2023_ (.CLK(clknet_leaf_34_clk),
    .D(booth_b20_m36),
    .Q(pp_row56_10));
 sky130_fd_sc_hd__dfxtp_1 _2024_ (.CLK(clknet_leaf_35_clk),
    .D(booth_b22_m34),
    .Q(pp_row56_11));
 sky130_fd_sc_hd__dfxtp_1 _2025_ (.CLK(clknet_leaf_36_clk),
    .D(booth_b24_m32),
    .Q(pp_row56_12));
 sky130_fd_sc_hd__dfxtp_1 _2026_ (.CLK(clknet_leaf_35_clk),
    .D(booth_b26_m30),
    .Q(pp_row56_13));
 sky130_fd_sc_hd__dfxtp_1 _2027_ (.CLK(clknet_leaf_135_clk),
    .D(booth_b60_m48),
    .Q(pp_row108_9));
 sky130_fd_sc_hd__dfxtp_1 _2028_ (.CLK(clknet_leaf_76_clk),
    .D(booth_b28_m28),
    .Q(pp_row56_14));
 sky130_fd_sc_hd__dfxtp_1 _2029_ (.CLK(clknet_leaf_76_clk),
    .D(booth_b30_m26),
    .Q(pp_row56_15));
 sky130_fd_sc_hd__dfxtp_1 _2030_ (.CLK(clknet_leaf_76_clk),
    .D(booth_b32_m24),
    .Q(pp_row56_16));
 sky130_fd_sc_hd__dfxtp_1 _2031_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b34_m22),
    .Q(pp_row56_17));
 sky130_fd_sc_hd__dfxtp_1 _2032_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b36_m20),
    .Q(pp_row56_18));
 sky130_fd_sc_hd__dfxtp_1 _2033_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b38_m18),
    .Q(pp_row56_19));
 sky130_fd_sc_hd__dfxtp_1 _2034_ (.CLK(clknet_leaf_73_clk),
    .D(booth_b40_m16),
    .Q(pp_row56_20));
 sky130_fd_sc_hd__dfxtp_1 _2035_ (.CLK(clknet_leaf_73_clk),
    .D(booth_b42_m14),
    .Q(pp_row56_21));
 sky130_fd_sc_hd__dfxtp_1 _2036_ (.CLK(clknet_leaf_72_clk),
    .D(booth_b44_m12),
    .Q(pp_row56_22));
 sky130_fd_sc_hd__dfxtp_1 _2037_ (.CLK(clknet_leaf_83_clk),
    .D(booth_b46_m10),
    .Q(pp_row56_23));
 sky130_fd_sc_hd__dfxtp_1 _2038_ (.CLK(clknet_leaf_135_clk),
    .D(booth_b62_m46),
    .Q(pp_row108_10));
 sky130_fd_sc_hd__dfxtp_1 _2039_ (.CLK(clknet_leaf_81_clk),
    .D(booth_b48_m8),
    .Q(pp_row56_24));
 sky130_fd_sc_hd__dfxtp_1 _2040_ (.CLK(clknet_leaf_83_clk),
    .D(booth_b50_m6),
    .Q(pp_row56_25));
 sky130_fd_sc_hd__dfxtp_1 _2041_ (.CLK(clknet_leaf_82_clk),
    .D(booth_b52_m4),
    .Q(pp_row56_26));
 sky130_fd_sc_hd__dfxtp_1 _2042_ (.CLK(clknet_leaf_82_clk),
    .D(booth_b54_m2),
    .Q(pp_row56_27));
 sky130_fd_sc_hd__dfxtp_1 _2043_ (.CLK(clknet_leaf_85_clk),
    .D(booth_b56_m0),
    .Q(pp_row56_28));
 sky130_fd_sc_hd__dfxtp_1 _2044_ (.CLK(clknet_leaf_83_clk),
    .D(net1296),
    .Q(pp_row56_29));
 sky130_fd_sc_hd__dfxtp_2 _2045_ (.CLK(clknet_leaf_231_clk),
    .D(net208),
    .Q(pp_row56_30));
 sky130_fd_sc_hd__dfxtp_1 _2046_ (.CLK(clknet_leaf_82_clk),
    .D(booth_b0_m57),
    .Q(pp_row57_0));
 sky130_fd_sc_hd__dfxtp_1 _2047_ (.CLK(clknet_leaf_82_clk),
    .D(booth_b2_m55),
    .Q(pp_row57_1));
 sky130_fd_sc_hd__dfxtp_1 _2048_ (.CLK(clknet_leaf_38_clk),
    .D(booth_b4_m53),
    .Q(pp_row57_2));
 sky130_fd_sc_hd__dfxtp_1 _2049_ (.CLK(clknet_leaf_136_clk),
    .D(booth_b64_m44),
    .Q(pp_row108_11));
 sky130_fd_sc_hd__dfxtp_1 _2050_ (.CLK(clknet_leaf_38_clk),
    .D(booth_b6_m51),
    .Q(pp_row57_3));
 sky130_fd_sc_hd__dfxtp_1 _2051_ (.CLK(clknet_leaf_38_clk),
    .D(booth_b8_m49),
    .Q(pp_row57_4));
 sky130_fd_sc_hd__dfxtp_1 _2052_ (.CLK(clknet_leaf_38_clk),
    .D(booth_b10_m47),
    .Q(pp_row57_5));
 sky130_fd_sc_hd__dfxtp_1 _2053_ (.CLK(clknet_leaf_38_clk),
    .D(booth_b12_m45),
    .Q(pp_row57_6));
 sky130_fd_sc_hd__dfxtp_1 _2054_ (.CLK(clknet_leaf_38_clk),
    .D(booth_b14_m43),
    .Q(pp_row57_7));
 sky130_fd_sc_hd__dfxtp_1 _2055_ (.CLK(clknet_leaf_38_clk),
    .D(booth_b16_m41),
    .Q(pp_row57_8));
 sky130_fd_sc_hd__dfxtp_1 _2056_ (.CLK(clknet_leaf_38_clk),
    .D(booth_b18_m39),
    .Q(pp_row57_9));
 sky130_fd_sc_hd__dfxtp_1 _2057_ (.CLK(clknet_leaf_36_clk),
    .D(booth_b20_m37),
    .Q(pp_row57_10));
 sky130_fd_sc_hd__dfxtp_1 _2058_ (.CLK(clknet_leaf_42_clk),
    .D(booth_b22_m35),
    .Q(pp_row57_11));
 sky130_fd_sc_hd__dfxtp_1 _2059_ (.CLK(clknet_leaf_39_clk),
    .D(booth_b24_m33),
    .Q(pp_row57_12));
 sky130_fd_sc_hd__dfxtp_2 _2060_ (.CLK(clknet_leaf_184_clk),
    .D(net138),
    .Q(pp_row108_12));
 sky130_fd_sc_hd__dfxtp_1 _2061_ (.CLK(clknet_leaf_164_clk),
    .D(booth_b62_m62),
    .Q(pp_row124_2));
 sky130_fd_sc_hd__dfxtp_1 _2062_ (.CLK(clknet_leaf_36_clk),
    .D(booth_b26_m31),
    .Q(pp_row57_13));
 sky130_fd_sc_hd__dfxtp_1 _2063_ (.CLK(clknet_leaf_43_clk),
    .D(booth_b28_m29),
    .Q(pp_row57_14));
 sky130_fd_sc_hd__dfxtp_1 _2064_ (.CLK(clknet_leaf_35_clk),
    .D(booth_b30_m27),
    .Q(pp_row57_15));
 sky130_fd_sc_hd__dfxtp_1 _2065_ (.CLK(clknet_leaf_34_clk),
    .D(booth_b32_m25),
    .Q(pp_row57_16));
 sky130_fd_sc_hd__dfxtp_1 _2066_ (.CLK(clknet_leaf_43_clk),
    .D(booth_b34_m23),
    .Q(pp_row57_17));
 sky130_fd_sc_hd__dfxtp_1 _2067_ (.CLK(clknet_leaf_35_clk),
    .D(booth_b36_m21),
    .Q(pp_row57_18));
 sky130_fd_sc_hd__dfxtp_1 _2068_ (.CLK(clknet_leaf_43_clk),
    .D(booth_b38_m19),
    .Q(pp_row57_19));
 sky130_fd_sc_hd__dfxtp_1 _2069_ (.CLK(clknet_leaf_35_clk),
    .D(booth_b40_m17),
    .Q(pp_row57_20));
 sky130_fd_sc_hd__dfxtp_1 _2070_ (.CLK(clknet_leaf_36_clk),
    .D(booth_b42_m15),
    .Q(pp_row57_21));
 sky130_fd_sc_hd__dfxtp_1 _2071_ (.CLK(clknet_leaf_35_clk),
    .D(booth_b44_m13),
    .Q(pp_row57_22));
 sky130_fd_sc_hd__dfxtp_1 _2072_ (.CLK(clknet_leaf_143_clk),
    .D(\notsign$6014 ),
    .Q(pp_row109_0));
 sky130_fd_sc_hd__dfxtp_1 _2073_ (.CLK(clknet_leaf_32_clk),
    .D(booth_b46_m11),
    .Q(pp_row57_23));
 sky130_fd_sc_hd__dfxtp_1 _2074_ (.CLK(clknet_leaf_32_clk),
    .D(booth_b48_m9),
    .Q(pp_row57_24));
 sky130_fd_sc_hd__dfxtp_1 _2075_ (.CLK(clknet_leaf_32_clk),
    .D(booth_b50_m7),
    .Q(pp_row57_25));
 sky130_fd_sc_hd__dfxtp_1 _2076_ (.CLK(clknet_leaf_85_clk),
    .D(booth_b52_m5),
    .Q(pp_row57_26));
 sky130_fd_sc_hd__dfxtp_1 _2077_ (.CLK(clknet_leaf_82_clk),
    .D(booth_b54_m3),
    .Q(pp_row57_27));
 sky130_fd_sc_hd__dfxtp_1 _2078_ (.CLK(clknet_leaf_85_clk),
    .D(booth_b56_m1),
    .Q(pp_row57_28));
 sky130_fd_sc_hd__dfxtp_2 _2079_ (.CLK(clknet_leaf_231_clk),
    .D(net209),
    .Q(pp_row57_29));
 sky130_fd_sc_hd__dfxtp_1 _2080_ (.CLK(clknet_leaf_86_clk),
    .D(booth_b0_m58),
    .Q(pp_row58_0));
 sky130_fd_sc_hd__dfxtp_1 _2081_ (.CLK(clknet_leaf_86_clk),
    .D(booth_b2_m56),
    .Q(pp_row58_1));
 sky130_fd_sc_hd__dfxtp_1 _2082_ (.CLK(clknet_leaf_86_clk),
    .D(booth_b4_m54),
    .Q(pp_row58_2));
 sky130_fd_sc_hd__dfxtp_1 _2083_ (.CLK(clknet_leaf_143_clk),
    .D(booth_b46_m63),
    .Q(pp_row109_1));
 sky130_fd_sc_hd__dfxtp_1 _2084_ (.CLK(clknet_leaf_31_clk),
    .D(booth_b6_m52),
    .Q(pp_row58_3));
 sky130_fd_sc_hd__dfxtp_1 _2085_ (.CLK(clknet_leaf_32_clk),
    .D(booth_b8_m50),
    .Q(pp_row58_4));
 sky130_fd_sc_hd__dfxtp_1 _2086_ (.CLK(clknet_leaf_32_clk),
    .D(booth_b10_m48),
    .Q(pp_row58_5));
 sky130_fd_sc_hd__dfxtp_1 _2087_ (.CLK(clknet_leaf_37_clk),
    .D(booth_b12_m46),
    .Q(pp_row58_6));
 sky130_fd_sc_hd__dfxtp_1 _2088_ (.CLK(clknet_leaf_37_clk),
    .D(booth_b14_m44),
    .Q(pp_row58_7));
 sky130_fd_sc_hd__dfxtp_1 _2089_ (.CLK(clknet_leaf_37_clk),
    .D(booth_b16_m42),
    .Q(pp_row58_8));
 sky130_fd_sc_hd__dfxtp_1 _2090_ (.CLK(clknet_leaf_37_clk),
    .D(booth_b18_m40),
    .Q(pp_row58_9));
 sky130_fd_sc_hd__dfxtp_1 _2091_ (.CLK(clknet_leaf_37_clk),
    .D(booth_b20_m38),
    .Q(pp_row58_10));
 sky130_fd_sc_hd__dfxtp_1 _2092_ (.CLK(clknet_leaf_149_clk),
    .D(booth_b22_m36),
    .Q(pp_row58_11));
 sky130_fd_sc_hd__dfxtp_1 _2093_ (.CLK(clknet_leaf_149_clk),
    .D(booth_b24_m34),
    .Q(pp_row58_12));
 sky130_fd_sc_hd__dfxtp_1 _2094_ (.CLK(clknet_leaf_143_clk),
    .D(booth_b48_m61),
    .Q(pp_row109_2));
 sky130_fd_sc_hd__dfxtp_1 _2095_ (.CLK(clknet_leaf_88_clk),
    .D(booth_b26_m32),
    .Q(pp_row58_13));
 sky130_fd_sc_hd__dfxtp_1 _2096_ (.CLK(clknet_leaf_86_clk),
    .D(booth_b28_m30),
    .Q(pp_row58_14));
 sky130_fd_sc_hd__dfxtp_1 _2097_ (.CLK(clknet_leaf_86_clk),
    .D(booth_b30_m28),
    .Q(pp_row58_15));
 sky130_fd_sc_hd__dfxtp_1 _2098_ (.CLK(clknet_leaf_86_clk),
    .D(booth_b32_m26),
    .Q(pp_row58_16));
 sky130_fd_sc_hd__dfxtp_1 _2099_ (.CLK(clknet_leaf_32_clk),
    .D(booth_b34_m24),
    .Q(pp_row58_17));
 sky130_fd_sc_hd__dfxtp_1 _2100_ (.CLK(clknet_leaf_32_clk),
    .D(booth_b36_m22),
    .Q(pp_row58_18));
 sky130_fd_sc_hd__dfxtp_1 _2101_ (.CLK(clknet_leaf_32_clk),
    .D(booth_b38_m20),
    .Q(pp_row58_19));
 sky130_fd_sc_hd__dfxtp_1 _2102_ (.CLK(clknet_leaf_29_clk),
    .D(booth_b40_m18),
    .Q(pp_row58_20));
 sky130_fd_sc_hd__dfxtp_1 _2103_ (.CLK(clknet_leaf_30_clk),
    .D(booth_b42_m16),
    .Q(pp_row58_21));
 sky130_fd_sc_hd__dfxtp_1 _2104_ (.CLK(clknet_leaf_30_clk),
    .D(booth_b44_m14),
    .Q(pp_row58_22));
 sky130_fd_sc_hd__dfxtp_1 _2105_ (.CLK(clknet_leaf_137_clk),
    .D(booth_b50_m59),
    .Q(pp_row109_3));
 sky130_fd_sc_hd__dfxtp_1 _2106_ (.CLK(clknet_leaf_33_clk),
    .D(booth_b46_m12),
    .Q(pp_row58_23));
 sky130_fd_sc_hd__dfxtp_1 _2107_ (.CLK(clknet_leaf_33_clk),
    .D(booth_b48_m10),
    .Q(pp_row58_24));
 sky130_fd_sc_hd__dfxtp_1 _2108_ (.CLK(clknet_leaf_33_clk),
    .D(booth_b50_m8),
    .Q(pp_row58_25));
 sky130_fd_sc_hd__dfxtp_1 _2109_ (.CLK(clknet_leaf_85_clk),
    .D(booth_b52_m6),
    .Q(pp_row58_26));
 sky130_fd_sc_hd__dfxtp_1 _2110_ (.CLK(clknet_leaf_86_clk),
    .D(booth_b54_m4),
    .Q(pp_row58_27));
 sky130_fd_sc_hd__dfxtp_1 _2111_ (.CLK(clknet_leaf_85_clk),
    .D(booth_b56_m2),
    .Q(pp_row58_28));
 sky130_fd_sc_hd__dfxtp_1 _2112_ (.CLK(clknet_leaf_86_clk),
    .D(booth_b58_m0),
    .Q(pp_row58_29));
 sky130_fd_sc_hd__dfxtp_1 _2113_ (.CLK(clknet_leaf_85_clk),
    .D(net1287),
    .Q(pp_row58_30));
 sky130_fd_sc_hd__dfxtp_2 _2114_ (.CLK(clknet_leaf_231_clk),
    .D(net210),
    .Q(pp_row58_31));
 sky130_fd_sc_hd__dfxtp_1 _2115_ (.CLK(clknet_leaf_218_clk),
    .D(booth_b0_m59),
    .Q(pp_row59_0));
 sky130_fd_sc_hd__dfxtp_1 _2116_ (.CLK(clknet_leaf_137_clk),
    .D(booth_b52_m57),
    .Q(pp_row109_4));
 sky130_fd_sc_hd__dfxtp_1 _2117_ (.CLK(clknet_leaf_224_clk),
    .D(booth_b2_m57),
    .Q(pp_row59_1));
 sky130_fd_sc_hd__dfxtp_1 _2118_ (.CLK(clknet_leaf_218_clk),
    .D(booth_b4_m55),
    .Q(pp_row59_2));
 sky130_fd_sc_hd__dfxtp_1 _2119_ (.CLK(clknet_leaf_218_clk),
    .D(booth_b6_m53),
    .Q(pp_row59_3));
 sky130_fd_sc_hd__dfxtp_1 _2120_ (.CLK(clknet_leaf_218_clk),
    .D(booth_b8_m51),
    .Q(pp_row59_4));
 sky130_fd_sc_hd__dfxtp_1 _2121_ (.CLK(clknet_leaf_218_clk),
    .D(booth_b10_m49),
    .Q(pp_row59_5));
 sky130_fd_sc_hd__dfxtp_1 _2122_ (.CLK(clknet_leaf_218_clk),
    .D(booth_b12_m47),
    .Q(pp_row59_6));
 sky130_fd_sc_hd__dfxtp_1 _2123_ (.CLK(clknet_leaf_219_clk),
    .D(booth_b14_m45),
    .Q(pp_row59_7));
 sky130_fd_sc_hd__dfxtp_1 _2124_ (.CLK(clknet_leaf_218_clk),
    .D(booth_b16_m43),
    .Q(pp_row59_8));
 sky130_fd_sc_hd__dfxtp_1 _2125_ (.CLK(clknet_leaf_217_clk),
    .D(booth_b18_m41),
    .Q(pp_row59_9));
 sky130_fd_sc_hd__dfxtp_1 _2126_ (.CLK(clknet_leaf_217_clk),
    .D(booth_b20_m39),
    .Q(pp_row59_10));
 sky130_fd_sc_hd__dfxtp_1 _2127_ (.CLK(clknet_leaf_129_clk),
    .D(booth_b54_m55),
    .Q(pp_row109_5));
 sky130_fd_sc_hd__dfxtp_1 _2128_ (.CLK(clknet_leaf_26_clk),
    .D(booth_b22_m37),
    .Q(pp_row59_11));
 sky130_fd_sc_hd__dfxtp_1 _2129_ (.CLK(clknet_leaf_29_clk),
    .D(booth_b24_m35),
    .Q(pp_row59_12));
 sky130_fd_sc_hd__dfxtp_1 _2130_ (.CLK(clknet_leaf_29_clk),
    .D(booth_b26_m33),
    .Q(pp_row59_13));
 sky130_fd_sc_hd__dfxtp_1 _2131_ (.CLK(clknet_leaf_32_clk),
    .D(booth_b28_m31),
    .Q(pp_row59_14));
 sky130_fd_sc_hd__dfxtp_1 _2132_ (.CLK(clknet_leaf_32_clk),
    .D(booth_b30_m29),
    .Q(pp_row59_15));
 sky130_fd_sc_hd__dfxtp_1 _2133_ (.CLK(clknet_leaf_32_clk),
    .D(booth_b32_m27),
    .Q(pp_row59_16));
 sky130_fd_sc_hd__dfxtp_1 _2134_ (.CLK(clknet_leaf_27_clk),
    .D(booth_b34_m25),
    .Q(pp_row59_17));
 sky130_fd_sc_hd__dfxtp_1 _2135_ (.CLK(clknet_leaf_27_clk),
    .D(booth_b36_m23),
    .Q(pp_row59_18));
 sky130_fd_sc_hd__dfxtp_1 _2136_ (.CLK(clknet_leaf_27_clk),
    .D(booth_b38_m21),
    .Q(pp_row59_19));
 sky130_fd_sc_hd__dfxtp_1 _2137_ (.CLK(clknet_leaf_26_clk),
    .D(booth_b40_m19),
    .Q(pp_row59_20));
 sky130_fd_sc_hd__dfxtp_1 _2138_ (.CLK(clknet_leaf_143_clk),
    .D(booth_b56_m53),
    .Q(pp_row109_6));
 sky130_fd_sc_hd__dfxtp_1 _2139_ (.CLK(clknet_leaf_26_clk),
    .D(booth_b42_m17),
    .Q(pp_row59_21));
 sky130_fd_sc_hd__dfxtp_1 _2140_ (.CLK(clknet_leaf_33_clk),
    .D(booth_b44_m15),
    .Q(pp_row59_22));
 sky130_fd_sc_hd__dfxtp_1 _2141_ (.CLK(clknet_leaf_219_clk),
    .D(booth_b46_m13),
    .Q(pp_row59_23));
 sky130_fd_sc_hd__dfxtp_1 _2142_ (.CLK(clknet_leaf_219_clk),
    .D(booth_b48_m11),
    .Q(pp_row59_24));
 sky130_fd_sc_hd__dfxtp_1 _2143_ (.CLK(clknet_leaf_219_clk),
    .D(booth_b50_m9),
    .Q(pp_row59_25));
 sky130_fd_sc_hd__dfxtp_1 _2144_ (.CLK(clknet_leaf_31_clk),
    .D(booth_b52_m7),
    .Q(pp_row59_26));
 sky130_fd_sc_hd__dfxtp_1 _2145_ (.CLK(clknet_leaf_31_clk),
    .D(booth_b54_m5),
    .Q(pp_row59_27));
 sky130_fd_sc_hd__dfxtp_1 _2146_ (.CLK(clknet_leaf_31_clk),
    .D(booth_b56_m3),
    .Q(pp_row59_28));
 sky130_fd_sc_hd__dfxtp_1 _2147_ (.CLK(clknet_leaf_87_clk),
    .D(booth_b58_m1),
    .Q(pp_row59_29));
 sky130_fd_sc_hd__dfxtp_2 _2148_ (.CLK(clknet_leaf_231_clk),
    .D(net211),
    .Q(pp_row59_30));
 sky130_fd_sc_hd__dfxtp_1 _2149_ (.CLK(clknet_leaf_144_clk),
    .D(booth_b58_m51),
    .Q(pp_row109_7));
 sky130_fd_sc_hd__dfxtp_1 _2150_ (.CLK(clknet_leaf_215_clk),
    .D(booth_b0_m60),
    .Q(pp_row60_0));
 sky130_fd_sc_hd__dfxtp_1 _2151_ (.CLK(clknet_leaf_215_clk),
    .D(booth_b2_m58),
    .Q(pp_row60_1));
 sky130_fd_sc_hd__dfxtp_1 _2152_ (.CLK(clknet_leaf_215_clk),
    .D(booth_b4_m56),
    .Q(pp_row60_2));
 sky130_fd_sc_hd__dfxtp_1 _2153_ (.CLK(clknet_leaf_214_clk),
    .D(booth_b6_m54),
    .Q(pp_row60_3));
 sky130_fd_sc_hd__dfxtp_1 _2154_ (.CLK(clknet_leaf_214_clk),
    .D(booth_b8_m52),
    .Q(pp_row60_4));
 sky130_fd_sc_hd__dfxtp_1 _2155_ (.CLK(clknet_leaf_214_clk),
    .D(booth_b10_m50),
    .Q(pp_row60_5));
 sky130_fd_sc_hd__dfxtp_1 _2156_ (.CLK(clknet_leaf_215_clk),
    .D(booth_b12_m48),
    .Q(pp_row60_6));
 sky130_fd_sc_hd__dfxtp_1 _2157_ (.CLK(clknet_leaf_215_clk),
    .D(booth_b14_m46),
    .Q(pp_row60_7));
 sky130_fd_sc_hd__dfxtp_1 _2158_ (.CLK(clknet_leaf_215_clk),
    .D(booth_b16_m44),
    .Q(pp_row60_8));
 sky130_fd_sc_hd__dfxtp_1 _2159_ (.CLK(clknet_leaf_214_clk),
    .D(booth_b18_m42),
    .Q(pp_row60_9));
 sky130_fd_sc_hd__dfxtp_1 _2160_ (.CLK(clknet_leaf_136_clk),
    .D(booth_b60_m49),
    .Q(pp_row109_8));
 sky130_fd_sc_hd__dfxtp_1 _2161_ (.CLK(clknet_leaf_214_clk),
    .D(booth_b20_m40),
    .Q(pp_row60_10));
 sky130_fd_sc_hd__dfxtp_1 _2162_ (.CLK(clknet_leaf_214_clk),
    .D(booth_b22_m38),
    .Q(pp_row60_11));
 sky130_fd_sc_hd__dfxtp_1 _2163_ (.CLK(clknet_leaf_30_clk),
    .D(booth_b24_m36),
    .Q(pp_row60_12));
 sky130_fd_sc_hd__dfxtp_1 _2164_ (.CLK(clknet_leaf_29_clk),
    .D(booth_b26_m34),
    .Q(pp_row60_13));
 sky130_fd_sc_hd__dfxtp_1 _2165_ (.CLK(clknet_leaf_28_clk),
    .D(booth_b28_m32),
    .Q(pp_row60_14));
 sky130_fd_sc_hd__dfxtp_1 _2166_ (.CLK(clknet_leaf_28_clk),
    .D(booth_b30_m30),
    .Q(pp_row60_15));
 sky130_fd_sc_hd__dfxtp_1 _2167_ (.CLK(clknet_leaf_27_clk),
    .D(booth_b32_m28),
    .Q(pp_row60_16));
 sky130_fd_sc_hd__dfxtp_1 _2168_ (.CLK(clknet_leaf_28_clk),
    .D(booth_b34_m26),
    .Q(pp_row60_17));
 sky130_fd_sc_hd__dfxtp_1 _2169_ (.CLK(clknet_leaf_215_clk),
    .D(booth_b36_m24),
    .Q(pp_row60_18));
 sky130_fd_sc_hd__dfxtp_1 _2170_ (.CLK(clknet_leaf_28_clk),
    .D(booth_b38_m22),
    .Q(pp_row60_19));
 sky130_fd_sc_hd__dfxtp_1 _2171_ (.CLK(clknet_leaf_136_clk),
    .D(booth_b62_m47),
    .Q(pp_row109_9));
 sky130_fd_sc_hd__dfxtp_1 _2172_ (.CLK(clknet_leaf_163_clk),
    .D(booth_b64_m60),
    .Q(pp_row124_3));
 sky130_fd_sc_hd__dfxtp_1 _2173_ (.CLK(clknet_leaf_224_clk),
    .D(booth_b40_m20),
    .Q(pp_row60_20));
 sky130_fd_sc_hd__dfxtp_1 _2174_ (.CLK(clknet_leaf_224_clk),
    .D(booth_b42_m18),
    .Q(pp_row60_21));
 sky130_fd_sc_hd__dfxtp_1 _2175_ (.CLK(clknet_leaf_224_clk),
    .D(booth_b44_m16),
    .Q(pp_row60_22));
 sky130_fd_sc_hd__dfxtp_1 _2176_ (.CLK(clknet_leaf_223_clk),
    .D(booth_b46_m14),
    .Q(pp_row60_23));
 sky130_fd_sc_hd__dfxtp_1 _2177_ (.CLK(clknet_leaf_224_clk),
    .D(booth_b48_m12),
    .Q(pp_row60_24));
 sky130_fd_sc_hd__dfxtp_1 _2178_ (.CLK(clknet_leaf_224_clk),
    .D(booth_b50_m10),
    .Q(pp_row60_25));
 sky130_fd_sc_hd__dfxtp_1 _2179_ (.CLK(clknet_leaf_218_clk),
    .D(booth_b52_m8),
    .Q(pp_row60_26));
 sky130_fd_sc_hd__dfxtp_1 _2180_ (.CLK(clknet_leaf_218_clk),
    .D(booth_b54_m6),
    .Q(pp_row60_27));
 sky130_fd_sc_hd__dfxtp_1 _2181_ (.CLK(clknet_leaf_218_clk),
    .D(booth_b56_m4),
    .Q(pp_row60_28));
 sky130_fd_sc_hd__dfxtp_1 _2182_ (.CLK(clknet_leaf_216_clk),
    .D(booth_b58_m2),
    .Q(pp_row60_29));
 sky130_fd_sc_hd__dfxtp_1 _2183_ (.CLK(clknet_leaf_136_clk),
    .D(booth_b64_m45),
    .Q(pp_row109_10));
 sky130_fd_sc_hd__dfxtp_1 _2184_ (.CLK(clknet_leaf_216_clk),
    .D(booth_b60_m0),
    .Q(pp_row60_30));
 sky130_fd_sc_hd__dfxtp_1 _2185_ (.CLK(clknet_leaf_216_clk),
    .D(net1263),
    .Q(pp_row60_31));
 sky130_fd_sc_hd__dfxtp_1 _2186_ (.CLK(clknet_leaf_231_clk),
    .D(net213),
    .Q(pp_row60_32));
 sky130_fd_sc_hd__dfxtp_1 _2187_ (.CLK(clknet_leaf_227_clk),
    .D(booth_b0_m61),
    .Q(pp_row61_0));
 sky130_fd_sc_hd__dfxtp_1 _2188_ (.CLK(clknet_leaf_227_clk),
    .D(booth_b2_m59),
    .Q(pp_row61_1));
 sky130_fd_sc_hd__dfxtp_1 _2189_ (.CLK(clknet_leaf_227_clk),
    .D(booth_b4_m57),
    .Q(pp_row61_2));
 sky130_fd_sc_hd__dfxtp_1 _2190_ (.CLK(clknet_leaf_223_clk),
    .D(booth_b6_m55),
    .Q(pp_row61_3));
 sky130_fd_sc_hd__dfxtp_1 _2191_ (.CLK(clknet_leaf_223_clk),
    .D(booth_b8_m53),
    .Q(pp_row61_4));
 sky130_fd_sc_hd__dfxtp_1 _2192_ (.CLK(clknet_leaf_223_clk),
    .D(booth_b10_m51),
    .Q(pp_row61_5));
 sky130_fd_sc_hd__dfxtp_1 _2193_ (.CLK(clknet_leaf_227_clk),
    .D(booth_b12_m49),
    .Q(pp_row61_6));
 sky130_fd_sc_hd__dfxtp_2 _2194_ (.CLK(clknet_leaf_184_clk),
    .D(net139),
    .Q(pp_row109_11));
 sky130_fd_sc_hd__dfxtp_1 _2195_ (.CLK(clknet_leaf_223_clk),
    .D(booth_b14_m47),
    .Q(pp_row61_7));
 sky130_fd_sc_hd__dfxtp_1 _2196_ (.CLK(clknet_leaf_223_clk),
    .D(booth_b16_m45),
    .Q(pp_row61_8));
 sky130_fd_sc_hd__dfxtp_1 _2197_ (.CLK(clknet_leaf_228_clk),
    .D(booth_b18_m43),
    .Q(pp_row61_9));
 sky130_fd_sc_hd__dfxtp_1 _2198_ (.CLK(clknet_leaf_228_clk),
    .D(booth_b20_m41),
    .Q(pp_row61_10));
 sky130_fd_sc_hd__dfxtp_1 _2199_ (.CLK(clknet_leaf_228_clk),
    .D(booth_b22_m39),
    .Q(pp_row61_11));
 sky130_fd_sc_hd__dfxtp_1 _2200_ (.CLK(clknet_leaf_228_clk),
    .D(booth_b24_m37),
    .Q(pp_row61_12));
 sky130_fd_sc_hd__dfxtp_1 _2201_ (.CLK(clknet_leaf_223_clk),
    .D(booth_b26_m35),
    .Q(pp_row61_13));
 sky130_fd_sc_hd__dfxtp_1 _2202_ (.CLK(clknet_leaf_88_clk),
    .D(booth_b28_m33),
    .Q(pp_row61_14));
 sky130_fd_sc_hd__dfxtp_1 _2203_ (.CLK(clknet_leaf_88_clk),
    .D(booth_b30_m31),
    .Q(pp_row61_15));
 sky130_fd_sc_hd__dfxtp_1 _2204_ (.CLK(clknet_leaf_88_clk),
    .D(booth_b32_m29),
    .Q(pp_row61_16));
 sky130_fd_sc_hd__dfxtp_1 _2205_ (.CLK(clknet_leaf_133_clk),
    .D(booth_b46_m64),
    .Q(pp_row110_1));
 sky130_fd_sc_hd__dfxtp_1 _2206_ (.CLK(clknet_leaf_29_clk),
    .D(booth_b34_m27),
    .Q(pp_row61_17));
 sky130_fd_sc_hd__dfxtp_1 _2207_ (.CLK(clknet_leaf_29_clk),
    .D(booth_b36_m25),
    .Q(pp_row61_18));
 sky130_fd_sc_hd__dfxtp_1 _2208_ (.CLK(clknet_leaf_29_clk),
    .D(booth_b38_m23),
    .Q(pp_row61_19));
 sky130_fd_sc_hd__dfxtp_1 _2209_ (.CLK(clknet_leaf_212_clk),
    .D(booth_b40_m21),
    .Q(pp_row61_20));
 sky130_fd_sc_hd__dfxtp_1 _2210_ (.CLK(clknet_leaf_212_clk),
    .D(booth_b42_m19),
    .Q(pp_row61_21));
 sky130_fd_sc_hd__dfxtp_1 _2211_ (.CLK(clknet_leaf_212_clk),
    .D(booth_b44_m17),
    .Q(pp_row61_22));
 sky130_fd_sc_hd__dfxtp_1 _2212_ (.CLK(clknet_leaf_217_clk),
    .D(booth_b46_m15),
    .Q(pp_row61_23));
 sky130_fd_sc_hd__dfxtp_1 _2213_ (.CLK(clknet_leaf_217_clk),
    .D(booth_b48_m13),
    .Q(pp_row61_24));
 sky130_fd_sc_hd__dfxtp_1 _2214_ (.CLK(clknet_leaf_217_clk),
    .D(booth_b50_m11),
    .Q(pp_row61_25));
 sky130_fd_sc_hd__dfxtp_1 _2215_ (.CLK(clknet_leaf_29_clk),
    .D(booth_b52_m9),
    .Q(pp_row61_26));
 sky130_fd_sc_hd__dfxtp_1 _2216_ (.CLK(clknet_leaf_133_clk),
    .D(booth_b48_m62),
    .Q(pp_row110_2));
 sky130_fd_sc_hd__dfxtp_1 _2217_ (.CLK(clknet_leaf_29_clk),
    .D(booth_b54_m7),
    .Q(pp_row61_27));
 sky130_fd_sc_hd__dfxtp_1 _2218_ (.CLK(clknet_leaf_29_clk),
    .D(booth_b56_m5),
    .Q(pp_row61_28));
 sky130_fd_sc_hd__dfxtp_1 _2219_ (.CLK(clknet_leaf_216_clk),
    .D(booth_b58_m3),
    .Q(pp_row61_29));
 sky130_fd_sc_hd__dfxtp_1 _2220_ (.CLK(clknet_leaf_215_clk),
    .D(booth_b60_m1),
    .Q(pp_row61_30));
 sky130_fd_sc_hd__dfxtp_1 _2221_ (.CLK(clknet_leaf_231_clk),
    .D(net214),
    .Q(pp_row61_31));
 sky130_fd_sc_hd__dfxtp_1 _2222_ (.CLK(clknet_leaf_229_clk),
    .D(booth_b0_m62),
    .Q(pp_row62_0));
 sky130_fd_sc_hd__dfxtp_1 _2223_ (.CLK(clknet_leaf_227_clk),
    .D(booth_b2_m60),
    .Q(pp_row62_1));
 sky130_fd_sc_hd__dfxtp_1 _2224_ (.CLK(clknet_leaf_227_clk),
    .D(booth_b4_m58),
    .Q(pp_row62_2));
 sky130_fd_sc_hd__dfxtp_1 _2225_ (.CLK(clknet_leaf_227_clk),
    .D(booth_b6_m56),
    .Q(pp_row62_3));
 sky130_fd_sc_hd__dfxtp_1 _2226_ (.CLK(clknet_leaf_227_clk),
    .D(booth_b8_m54),
    .Q(pp_row62_4));
 sky130_fd_sc_hd__dfxtp_1 _2227_ (.CLK(clknet_leaf_136_clk),
    .D(booth_b50_m60),
    .Q(pp_row110_3));
 sky130_fd_sc_hd__dfxtp_1 _2228_ (.CLK(clknet_leaf_227_clk),
    .D(booth_b10_m52),
    .Q(pp_row62_5));
 sky130_fd_sc_hd__dfxtp_1 _2229_ (.CLK(clknet_leaf_229_clk),
    .D(booth_b12_m50),
    .Q(pp_row62_6));
 sky130_fd_sc_hd__dfxtp_1 _2230_ (.CLK(clknet_leaf_233_clk),
    .D(booth_b14_m48),
    .Q(pp_row62_7));
 sky130_fd_sc_hd__dfxtp_1 _2231_ (.CLK(clknet_leaf_233_clk),
    .D(booth_b16_m46),
    .Q(pp_row62_8));
 sky130_fd_sc_hd__dfxtp_1 _2232_ (.CLK(clknet_leaf_233_clk),
    .D(booth_b18_m44),
    .Q(pp_row62_9));
 sky130_fd_sc_hd__dfxtp_1 _2233_ (.CLK(clknet_leaf_233_clk),
    .D(booth_b20_m42),
    .Q(pp_row62_10));
 sky130_fd_sc_hd__dfxtp_1 _2234_ (.CLK(clknet_leaf_232_clk),
    .D(booth_b22_m40),
    .Q(pp_row62_11));
 sky130_fd_sc_hd__dfxtp_1 _2235_ (.CLK(clknet_leaf_228_clk),
    .D(booth_b24_m38),
    .Q(pp_row62_12));
 sky130_fd_sc_hd__dfxtp_1 _2236_ (.CLK(clknet_leaf_228_clk),
    .D(booth_b26_m36),
    .Q(pp_row62_13));
 sky130_fd_sc_hd__dfxtp_1 _2237_ (.CLK(clknet_leaf_228_clk),
    .D(booth_b28_m34),
    .Q(pp_row62_14));
 sky130_fd_sc_hd__dfxtp_1 _2238_ (.CLK(clknet_leaf_136_clk),
    .D(booth_b52_m58),
    .Q(pp_row110_4));
 sky130_fd_sc_hd__dfxtp_1 _2239_ (.CLK(clknet_leaf_230_clk),
    .D(booth_b30_m32),
    .Q(pp_row62_15));
 sky130_fd_sc_hd__dfxtp_1 _2240_ (.CLK(clknet_leaf_227_clk),
    .D(booth_b32_m30),
    .Q(pp_row62_16));
 sky130_fd_sc_hd__dfxtp_1 _2241_ (.CLK(clknet_leaf_148_clk),
    .D(booth_b34_m28),
    .Q(pp_row62_17));
 sky130_fd_sc_hd__dfxtp_1 _2242_ (.CLK(clknet_leaf_150_clk),
    .D(booth_b36_m26),
    .Q(pp_row62_18));
 sky130_fd_sc_hd__dfxtp_1 _2243_ (.CLK(clknet_leaf_150_clk),
    .D(booth_b38_m24),
    .Q(pp_row62_19));
 sky130_fd_sc_hd__dfxtp_1 _2244_ (.CLK(clknet_leaf_30_clk),
    .D(booth_b40_m22),
    .Q(pp_row62_20));
 sky130_fd_sc_hd__dfxtp_1 _2245_ (.CLK(clknet_leaf_29_clk),
    .D(booth_b42_m20),
    .Q(pp_row62_21));
 sky130_fd_sc_hd__dfxtp_1 _2246_ (.CLK(clknet_leaf_30_clk),
    .D(booth_b44_m18),
    .Q(pp_row62_22));
 sky130_fd_sc_hd__dfxtp_1 _2247_ (.CLK(clknet_leaf_213_clk),
    .D(booth_b46_m16),
    .Q(pp_row62_23));
 sky130_fd_sc_hd__dfxtp_1 _2248_ (.CLK(clknet_leaf_149_clk),
    .D(booth_b48_m14),
    .Q(pp_row62_24));
 sky130_fd_sc_hd__dfxtp_1 _2249_ (.CLK(clknet_leaf_136_clk),
    .D(booth_b54_m56),
    .Q(pp_row110_5));
 sky130_fd_sc_hd__dfxtp_1 _2250_ (.CLK(clknet_leaf_149_clk),
    .D(booth_b50_m12),
    .Q(pp_row62_25));
 sky130_fd_sc_hd__dfxtp_1 _2251_ (.CLK(clknet_leaf_212_clk),
    .D(booth_b52_m10),
    .Q(pp_row62_26));
 sky130_fd_sc_hd__dfxtp_1 _2252_ (.CLK(clknet_leaf_149_clk),
    .D(booth_b54_m8),
    .Q(pp_row62_27));
 sky130_fd_sc_hd__dfxtp_1 _2253_ (.CLK(clknet_leaf_150_clk),
    .D(booth_b56_m6),
    .Q(pp_row62_28));
 sky130_fd_sc_hd__dfxtp_1 _2254_ (.CLK(clknet_leaf_148_clk),
    .D(booth_b58_m4),
    .Q(pp_row62_29));
 sky130_fd_sc_hd__dfxtp_1 _2255_ (.CLK(clknet_leaf_149_clk),
    .D(booth_b60_m2),
    .Q(pp_row62_30));
 sky130_fd_sc_hd__dfxtp_1 _2256_ (.CLK(clknet_leaf_149_clk),
    .D(booth_b62_m0),
    .Q(pp_row62_31));
 sky130_fd_sc_hd__dfxtp_1 _2257_ (.CLK(clknet_leaf_227_clk),
    .D(net1254),
    .Q(pp_row62_32));
 sky130_fd_sc_hd__dfxtp_1 _2258_ (.CLK(clknet_leaf_231_clk),
    .D(net215),
    .Q(pp_row62_33));
 sky130_fd_sc_hd__dfxtp_1 _2259_ (.CLK(clknet_leaf_230_clk),
    .D(booth_b0_m63),
    .Q(pp_row63_0));
 sky130_fd_sc_hd__dfxtp_1 _2260_ (.CLK(clknet_leaf_137_clk),
    .D(booth_b56_m54),
    .Q(pp_row110_6));
 sky130_fd_sc_hd__dfxtp_1 _2261_ (.CLK(clknet_leaf_199_clk),
    .D(booth_b2_m61),
    .Q(pp_row63_1));
 sky130_fd_sc_hd__dfxtp_1 _2262_ (.CLK(clknet_leaf_230_clk),
    .D(booth_b4_m59),
    .Q(pp_row63_2));
 sky130_fd_sc_hd__dfxtp_1 _2263_ (.CLK(clknet_leaf_230_clk),
    .D(booth_b6_m57),
    .Q(pp_row63_3));
 sky130_fd_sc_hd__dfxtp_1 _2264_ (.CLK(clknet_leaf_230_clk),
    .D(booth_b8_m55),
    .Q(pp_row63_4));
 sky130_fd_sc_hd__dfxtp_1 _2265_ (.CLK(clknet_leaf_230_clk),
    .D(booth_b10_m53),
    .Q(pp_row63_5));
 sky130_fd_sc_hd__dfxtp_1 _2266_ (.CLK(clknet_leaf_214_clk),
    .D(booth_b12_m51),
    .Q(pp_row63_6));
 sky130_fd_sc_hd__dfxtp_1 _2267_ (.CLK(clknet_leaf_214_clk),
    .D(booth_b14_m49),
    .Q(pp_row63_7));
 sky130_fd_sc_hd__dfxtp_1 _2268_ (.CLK(clknet_leaf_214_clk),
    .D(booth_b16_m47),
    .Q(pp_row63_8));
 sky130_fd_sc_hd__dfxtp_1 _2269_ (.CLK(clknet_leaf_210_clk),
    .D(booth_b18_m45),
    .Q(pp_row63_9));
 sky130_fd_sc_hd__dfxtp_1 _2270_ (.CLK(clknet_leaf_210_clk),
    .D(booth_b20_m43),
    .Q(pp_row63_10));
 sky130_fd_sc_hd__dfxtp_1 _2271_ (.CLK(clknet_leaf_129_clk),
    .D(booth_b58_m52),
    .Q(pp_row110_7));
 sky130_fd_sc_hd__dfxtp_1 _2272_ (.CLK(clknet_leaf_210_clk),
    .D(booth_b22_m41),
    .Q(pp_row63_11));
 sky130_fd_sc_hd__dfxtp_1 _2273_ (.CLK(clknet_leaf_216_clk),
    .D(booth_b24_m39),
    .Q(pp_row63_12));
 sky130_fd_sc_hd__dfxtp_1 _2274_ (.CLK(clknet_leaf_209_clk),
    .D(booth_b26_m37),
    .Q(pp_row63_13));
 sky130_fd_sc_hd__dfxtp_1 _2275_ (.CLK(clknet_leaf_217_clk),
    .D(booth_b28_m35),
    .Q(pp_row63_14));
 sky130_fd_sc_hd__dfxtp_1 _2276_ (.CLK(clknet_leaf_213_clk),
    .D(booth_b30_m33),
    .Q(pp_row63_15));
 sky130_fd_sc_hd__dfxtp_1 _2277_ (.CLK(clknet_leaf_212_clk),
    .D(booth_b32_m31),
    .Q(pp_row63_16));
 sky130_fd_sc_hd__dfxtp_1 _2278_ (.CLK(clknet_leaf_212_clk),
    .D(booth_b34_m29),
    .Q(pp_row63_17));
 sky130_fd_sc_hd__dfxtp_1 _2279_ (.CLK(clknet_leaf_212_clk),
    .D(booth_b36_m27),
    .Q(pp_row63_18));
 sky130_fd_sc_hd__dfxtp_1 _2280_ (.CLK(clknet_leaf_212_clk),
    .D(booth_b38_m25),
    .Q(pp_row63_19));
 sky130_fd_sc_hd__dfxtp_1 _2281_ (.CLK(clknet_leaf_153_clk),
    .D(booth_b40_m23),
    .Q(pp_row63_20));
 sky130_fd_sc_hd__dfxtp_1 _2282_ (.CLK(clknet_leaf_129_clk),
    .D(booth_b60_m50),
    .Q(pp_row110_8));
 sky130_fd_sc_hd__dfxtp_1 _2283_ (.CLK(clknet_leaf_181_clk),
    .D(net156),
    .Q(pp_row124_4));
 sky130_fd_sc_hd__dfxtp_1 _2284_ (.CLK(clknet_leaf_152_clk),
    .D(booth_b42_m21),
    .Q(pp_row63_21));
 sky130_fd_sc_hd__dfxtp_1 _2285_ (.CLK(clknet_leaf_152_clk),
    .D(booth_b44_m19),
    .Q(pp_row63_22));
 sky130_fd_sc_hd__dfxtp_1 _2286_ (.CLK(clknet_leaf_216_clk),
    .D(booth_b46_m17),
    .Q(pp_row63_23));
 sky130_fd_sc_hd__dfxtp_1 _2287_ (.CLK(clknet_leaf_210_clk),
    .D(booth_b48_m15),
    .Q(pp_row63_24));
 sky130_fd_sc_hd__dfxtp_1 _2288_ (.CLK(clknet_leaf_210_clk),
    .D(booth_b50_m13),
    .Q(pp_row63_25));
 sky130_fd_sc_hd__dfxtp_1 _2289_ (.CLK(clknet_leaf_214_clk),
    .D(booth_b52_m11),
    .Q(pp_row63_26));
 sky130_fd_sc_hd__dfxtp_1 _2290_ (.CLK(clknet_leaf_216_clk),
    .D(booth_b54_m9),
    .Q(pp_row63_27));
 sky130_fd_sc_hd__dfxtp_1 _2291_ (.CLK(clknet_leaf_214_clk),
    .D(booth_b56_m7),
    .Q(pp_row63_28));
 sky130_fd_sc_hd__dfxtp_1 _2292_ (.CLK(clknet_leaf_212_clk),
    .D(booth_b58_m5),
    .Q(pp_row63_29));
 sky130_fd_sc_hd__dfxtp_1 _2293_ (.CLK(clknet_leaf_212_clk),
    .D(booth_b60_m3),
    .Q(pp_row63_30));
 sky130_fd_sc_hd__dfxtp_1 _2294_ (.CLK(clknet_leaf_130_clk),
    .D(booth_b62_m48),
    .Q(pp_row110_9));
 sky130_fd_sc_hd__dfxtp_1 _2295_ (.CLK(clknet_leaf_209_clk),
    .D(booth_b62_m1),
    .Q(pp_row63_31));
 sky130_fd_sc_hd__dfxtp_1 _2296_ (.CLK(clknet_leaf_231_clk),
    .D(net216),
    .Q(pp_row63_32));
 sky130_fd_sc_hd__dfxtp_1 _2297_ (.CLK(clknet_leaf_199_clk),
    .D(booth_b0_m64),
    .Q(pp_row64_0));
 sky130_fd_sc_hd__dfxtp_1 _2298_ (.CLK(clknet_leaf_199_clk),
    .D(booth_b2_m62),
    .Q(pp_row64_1));
 sky130_fd_sc_hd__dfxtp_1 _2299_ (.CLK(clknet_leaf_199_clk),
    .D(booth_b4_m60),
    .Q(pp_row64_2));
 sky130_fd_sc_hd__dfxtp_1 _2300_ (.CLK(clknet_leaf_198_clk),
    .D(booth_b6_m58),
    .Q(pp_row64_3));
 sky130_fd_sc_hd__dfxtp_1 _2301_ (.CLK(clknet_leaf_198_clk),
    .D(booth_b8_m56),
    .Q(pp_row64_4));
 sky130_fd_sc_hd__dfxtp_1 _2302_ (.CLK(clknet_leaf_198_clk),
    .D(booth_b10_m54),
    .Q(pp_row64_5));
 sky130_fd_sc_hd__dfxtp_1 _2303_ (.CLK(clknet_leaf_91_clk),
    .D(booth_b12_m52),
    .Q(pp_row64_6));
 sky130_fd_sc_hd__dfxtp_1 _2304_ (.CLK(clknet_leaf_91_clk),
    .D(booth_b14_m50),
    .Q(pp_row64_7));
 sky130_fd_sc_hd__dfxtp_1 _2305_ (.CLK(clknet_leaf_133_clk),
    .D(booth_b64_m46),
    .Q(pp_row110_10));
 sky130_fd_sc_hd__dfxtp_1 _2306_ (.CLK(clknet_leaf_84_clk),
    .D(booth_b16_m48),
    .Q(pp_row64_8));
 sky130_fd_sc_hd__dfxtp_1 _2307_ (.CLK(clknet_leaf_91_clk),
    .D(booth_b18_m46),
    .Q(pp_row64_9));
 sky130_fd_sc_hd__dfxtp_1 _2308_ (.CLK(clknet_leaf_90_clk),
    .D(booth_b20_m44),
    .Q(pp_row64_10));
 sky130_fd_sc_hd__dfxtp_1 _2309_ (.CLK(clknet_leaf_91_clk),
    .D(booth_b22_m42),
    .Q(pp_row64_11));
 sky130_fd_sc_hd__dfxtp_1 _2310_ (.CLK(clknet_leaf_84_clk),
    .D(booth_b24_m40),
    .Q(pp_row64_12));
 sky130_fd_sc_hd__dfxtp_1 _2311_ (.CLK(clknet_leaf_85_clk),
    .D(booth_b26_m38),
    .Q(pp_row64_13));
 sky130_fd_sc_hd__dfxtp_1 _2312_ (.CLK(clknet_leaf_87_clk),
    .D(booth_b28_m36),
    .Q(pp_row64_14));
 sky130_fd_sc_hd__dfxtp_1 _2313_ (.CLK(clknet_leaf_30_clk),
    .D(booth_b30_m34),
    .Q(pp_row64_15));
 sky130_fd_sc_hd__dfxtp_1 _2314_ (.CLK(clknet_leaf_30_clk),
    .D(booth_b32_m32),
    .Q(pp_row64_16));
 sky130_fd_sc_hd__dfxtp_1 _2315_ (.CLK(clknet_leaf_30_clk),
    .D(booth_b34_m30),
    .Q(pp_row64_17));
 sky130_fd_sc_hd__dfxtp_2 _2316_ (.CLK(clknet_leaf_184_clk),
    .D(net141),
    .Q(pp_row110_11));
 sky130_fd_sc_hd__dfxtp_1 _2317_ (.CLK(clknet_leaf_96_clk),
    .D(booth_b36_m28),
    .Q(pp_row64_18));
 sky130_fd_sc_hd__dfxtp_1 _2318_ (.CLK(clknet_leaf_77_clk),
    .D(booth_b38_m26),
    .Q(pp_row64_19));
 sky130_fd_sc_hd__dfxtp_1 _2319_ (.CLK(clknet_leaf_77_clk),
    .D(booth_b40_m24),
    .Q(pp_row64_20));
 sky130_fd_sc_hd__dfxtp_1 _2320_ (.CLK(clknet_leaf_77_clk),
    .D(booth_b42_m22),
    .Q(pp_row64_21));
 sky130_fd_sc_hd__dfxtp_1 _2321_ (.CLK(clknet_leaf_77_clk),
    .D(booth_b44_m20),
    .Q(pp_row64_22));
 sky130_fd_sc_hd__dfxtp_1 _2322_ (.CLK(clknet_leaf_77_clk),
    .D(booth_b46_m18),
    .Q(pp_row64_23));
 sky130_fd_sc_hd__dfxtp_1 _2323_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b48_m16),
    .Q(pp_row64_24));
 sky130_fd_sc_hd__dfxtp_1 _2324_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b50_m14),
    .Q(pp_row64_25));
 sky130_fd_sc_hd__dfxtp_1 _2325_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b52_m12),
    .Q(pp_row64_26));
 sky130_fd_sc_hd__dfxtp_1 _2326_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b54_m10),
    .Q(pp_row64_27));
 sky130_fd_sc_hd__dfxtp_1 _2327_ (.CLK(clknet_leaf_127_clk),
    .D(\notsign$6084 ),
    .Q(pp_row111_0));
 sky130_fd_sc_hd__dfxtp_1 _2328_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b56_m8),
    .Q(pp_row64_28));
 sky130_fd_sc_hd__dfxtp_1 _2329_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b58_m6),
    .Q(pp_row64_29));
 sky130_fd_sc_hd__dfxtp_1 _2330_ (.CLK(clknet_leaf_99_clk),
    .D(booth_b60_m4),
    .Q(pp_row64_30));
 sky130_fd_sc_hd__dfxtp_1 _2331_ (.CLK(clknet_leaf_99_clk),
    .D(booth_b62_m2),
    .Q(pp_row64_31));
 sky130_fd_sc_hd__dfxtp_1 _2332_ (.CLK(clknet_leaf_100_clk),
    .D(booth_b64_m0),
    .Q(pp_row64_32));
 sky130_fd_sc_hd__dfxtp_1 _2333_ (.CLK(clknet_leaf_198_clk),
    .D(net217),
    .Q(pp_row64_33));
 sky130_fd_sc_hd__dfxtp_1 _2334_ (.CLK(clknet_leaf_86_clk),
    .D(booth_b2_m63),
    .Q(pp_row65_1));
 sky130_fd_sc_hd__dfxtp_1 _2335_ (.CLK(clknet_leaf_86_clk),
    .D(booth_b4_m61),
    .Q(pp_row65_2));
 sky130_fd_sc_hd__dfxtp_1 _2336_ (.CLK(clknet_leaf_89_clk),
    .D(booth_b6_m59),
    .Q(pp_row65_3));
 sky130_fd_sc_hd__dfxtp_1 _2337_ (.CLK(clknet_leaf_127_clk),
    .D(booth_b48_m63),
    .Q(pp_row111_1));
 sky130_fd_sc_hd__dfxtp_1 _2338_ (.CLK(clknet_leaf_91_clk),
    .D(booth_b8_m57),
    .Q(pp_row65_4));
 sky130_fd_sc_hd__dfxtp_1 _2339_ (.CLK(clknet_leaf_89_clk),
    .D(booth_b10_m55),
    .Q(pp_row65_5));
 sky130_fd_sc_hd__dfxtp_1 _2340_ (.CLK(clknet_leaf_89_clk),
    .D(booth_b12_m53),
    .Q(pp_row65_6));
 sky130_fd_sc_hd__dfxtp_1 _2341_ (.CLK(clknet_leaf_89_clk),
    .D(booth_b14_m51),
    .Q(pp_row65_7));
 sky130_fd_sc_hd__dfxtp_1 _2342_ (.CLK(clknet_leaf_89_clk),
    .D(booth_b16_m49),
    .Q(pp_row65_8));
 sky130_fd_sc_hd__dfxtp_1 _2343_ (.CLK(clknet_leaf_87_clk),
    .D(booth_b18_m47),
    .Q(pp_row65_9));
 sky130_fd_sc_hd__dfxtp_1 _2344_ (.CLK(clknet_leaf_87_clk),
    .D(booth_b20_m45),
    .Q(pp_row65_10));
 sky130_fd_sc_hd__dfxtp_1 _2345_ (.CLK(clknet_leaf_87_clk),
    .D(booth_b22_m43),
    .Q(pp_row65_11));
 sky130_fd_sc_hd__dfxtp_1 _2346_ (.CLK(clknet_leaf_88_clk),
    .D(booth_b24_m41),
    .Q(pp_row65_12));
 sky130_fd_sc_hd__dfxtp_1 _2347_ (.CLK(clknet_leaf_88_clk),
    .D(booth_b26_m39),
    .Q(pp_row65_13));
 sky130_fd_sc_hd__dfxtp_1 _2348_ (.CLK(clknet_leaf_127_clk),
    .D(booth_b50_m61),
    .Q(pp_row111_2));
 sky130_fd_sc_hd__dfxtp_1 _2349_ (.CLK(clknet_leaf_88_clk),
    .D(booth_b28_m37),
    .Q(pp_row65_14));
 sky130_fd_sc_hd__dfxtp_1 _2350_ (.CLK(clknet_leaf_77_clk),
    .D(booth_b30_m35),
    .Q(pp_row65_15));
 sky130_fd_sc_hd__dfxtp_1 _2351_ (.CLK(clknet_leaf_77_clk),
    .D(booth_b32_m33),
    .Q(pp_row65_16));
 sky130_fd_sc_hd__dfxtp_1 _2352_ (.CLK(clknet_leaf_77_clk),
    .D(booth_b34_m31),
    .Q(pp_row65_17));
 sky130_fd_sc_hd__dfxtp_1 _2353_ (.CLK(clknet_leaf_77_clk),
    .D(booth_b36_m29),
    .Q(pp_row65_18));
 sky130_fd_sc_hd__dfxtp_1 _2354_ (.CLK(clknet_leaf_75_clk),
    .D(booth_b38_m27),
    .Q(pp_row65_19));
 sky130_fd_sc_hd__dfxtp_1 _2355_ (.CLK(clknet_leaf_75_clk),
    .D(booth_b40_m25),
    .Q(pp_row65_20));
 sky130_fd_sc_hd__dfxtp_1 _2356_ (.CLK(clknet_leaf_98_clk),
    .D(booth_b42_m23),
    .Q(pp_row65_21));
 sky130_fd_sc_hd__dfxtp_1 _2357_ (.CLK(clknet_leaf_75_clk),
    .D(booth_b44_m21),
    .Q(pp_row65_22));
 sky130_fd_sc_hd__dfxtp_1 _2358_ (.CLK(clknet_leaf_77_clk),
    .D(booth_b46_m19),
    .Q(pp_row65_23));
 sky130_fd_sc_hd__dfxtp_1 _2359_ (.CLK(clknet_leaf_127_clk),
    .D(booth_b52_m59),
    .Q(pp_row111_3));
 sky130_fd_sc_hd__dfxtp_1 _2360_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b48_m17),
    .Q(pp_row65_24));
 sky130_fd_sc_hd__dfxtp_1 _2361_ (.CLK(clknet_leaf_75_clk),
    .D(booth_b50_m15),
    .Q(pp_row65_25));
 sky130_fd_sc_hd__dfxtp_1 _2362_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b52_m13),
    .Q(pp_row65_26));
 sky130_fd_sc_hd__dfxtp_1 _2363_ (.CLK(clknet_leaf_98_clk),
    .D(booth_b54_m11),
    .Q(pp_row65_27));
 sky130_fd_sc_hd__dfxtp_1 _2364_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b56_m9),
    .Q(pp_row65_28));
 sky130_fd_sc_hd__dfxtp_1 _2365_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b58_m7),
    .Q(pp_row65_29));
 sky130_fd_sc_hd__dfxtp_1 _2366_ (.CLK(clknet_leaf_98_clk),
    .D(booth_b60_m5),
    .Q(pp_row65_30));
 sky130_fd_sc_hd__dfxtp_1 _2367_ (.CLK(clknet_leaf_98_clk),
    .D(booth_b62_m3),
    .Q(pp_row65_31));
 sky130_fd_sc_hd__dfxtp_1 _2368_ (.CLK(clknet_leaf_98_clk),
    .D(booth_b64_m1),
    .Q(pp_row65_32));
 sky130_fd_sc_hd__dfxtp_1 _2369_ (.CLK(clknet_leaf_198_clk),
    .D(net218),
    .Q(pp_row65_33));
 sky130_fd_sc_hd__dfxtp_1 _2370_ (.CLK(clknet_leaf_127_clk),
    .D(booth_b54_m57),
    .Q(pp_row111_4));
 sky130_fd_sc_hd__dfxtp_1 _2371_ (.CLK(clknet_leaf_85_clk),
    .D(booth_b2_m64),
    .Q(pp_row66_1));
 sky130_fd_sc_hd__dfxtp_1 _2372_ (.CLK(clknet_leaf_85_clk),
    .D(booth_b4_m62),
    .Q(pp_row66_2));
 sky130_fd_sc_hd__dfxtp_1 _2373_ (.CLK(clknet_leaf_84_clk),
    .D(booth_b6_m60),
    .Q(pp_row66_3));
 sky130_fd_sc_hd__dfxtp_1 _2374_ (.CLK(clknet_leaf_84_clk),
    .D(booth_b8_m58),
    .Q(pp_row66_4));
 sky130_fd_sc_hd__dfxtp_1 _2375_ (.CLK(clknet_leaf_85_clk),
    .D(booth_b10_m56),
    .Q(pp_row66_5));
 sky130_fd_sc_hd__dfxtp_1 _2376_ (.CLK(clknet_leaf_85_clk),
    .D(booth_b12_m54),
    .Q(pp_row66_6));
 sky130_fd_sc_hd__dfxtp_1 _2377_ (.CLK(clknet_leaf_83_clk),
    .D(booth_b14_m52),
    .Q(pp_row66_7));
 sky130_fd_sc_hd__dfxtp_1 _2378_ (.CLK(clknet_leaf_83_clk),
    .D(booth_b16_m50),
    .Q(pp_row66_8));
 sky130_fd_sc_hd__dfxtp_1 _2379_ (.CLK(clknet_leaf_83_clk),
    .D(booth_b18_m48),
    .Q(pp_row66_9));
 sky130_fd_sc_hd__dfxtp_1 _2380_ (.CLK(clknet_leaf_127_clk),
    .D(booth_b56_m55),
    .Q(pp_row111_5));
 sky130_fd_sc_hd__dfxtp_1 _2381_ (.CLK(clknet_leaf_83_clk),
    .D(booth_b20_m46),
    .Q(pp_row66_10));
 sky130_fd_sc_hd__dfxtp_1 _2382_ (.CLK(clknet_leaf_83_clk),
    .D(booth_b22_m44),
    .Q(pp_row66_11));
 sky130_fd_sc_hd__dfxtp_1 _2383_ (.CLK(clknet_leaf_83_clk),
    .D(booth_b24_m42),
    .Q(pp_row66_12));
 sky130_fd_sc_hd__dfxtp_1 _2384_ (.CLK(clknet_leaf_83_clk),
    .D(booth_b26_m40),
    .Q(pp_row66_13));
 sky130_fd_sc_hd__dfxtp_1 _2385_ (.CLK(clknet_leaf_83_clk),
    .D(booth_b28_m38),
    .Q(pp_row66_14));
 sky130_fd_sc_hd__dfxtp_1 _2386_ (.CLK(clknet_leaf_77_clk),
    .D(booth_b30_m36),
    .Q(pp_row66_15));
 sky130_fd_sc_hd__dfxtp_1 _2387_ (.CLK(clknet_leaf_77_clk),
    .D(booth_b32_m34),
    .Q(pp_row66_16));
 sky130_fd_sc_hd__dfxtp_1 _2388_ (.CLK(clknet_leaf_77_clk),
    .D(booth_b34_m32),
    .Q(pp_row66_17));
 sky130_fd_sc_hd__dfxtp_1 _2389_ (.CLK(clknet_leaf_96_clk),
    .D(booth_b36_m30),
    .Q(pp_row66_18));
 sky130_fd_sc_hd__dfxtp_1 _2390_ (.CLK(clknet_leaf_96_clk),
    .D(booth_b38_m28),
    .Q(pp_row66_19));
 sky130_fd_sc_hd__dfxtp_1 _2391_ (.CLK(clknet_leaf_128_clk),
    .D(booth_b58_m53),
    .Q(pp_row111_6));
 sky130_fd_sc_hd__dfxtp_1 _2392_ (.CLK(clknet_leaf_179_clk),
    .D(\notsign$6574 ),
    .Q(pp_row125_0));
 sky130_fd_sc_hd__dfxtp_1 _2393_ (.CLK(clknet_leaf_96_clk),
    .D(booth_b40_m26),
    .Q(pp_row66_20));
 sky130_fd_sc_hd__dfxtp_1 _2394_ (.CLK(clknet_leaf_96_clk),
    .D(booth_b42_m24),
    .Q(pp_row66_21));
 sky130_fd_sc_hd__dfxtp_1 _2395_ (.CLK(clknet_leaf_96_clk),
    .D(booth_b44_m22),
    .Q(pp_row66_22));
 sky130_fd_sc_hd__dfxtp_1 _2396_ (.CLK(clknet_leaf_96_clk),
    .D(booth_b46_m20),
    .Q(pp_row66_23));
 sky130_fd_sc_hd__dfxtp_1 _2397_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b48_m18),
    .Q(pp_row66_24));
 sky130_fd_sc_hd__dfxtp_1 _2398_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b50_m16),
    .Q(pp_row66_25));
 sky130_fd_sc_hd__dfxtp_1 _2399_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b52_m14),
    .Q(pp_row66_26));
 sky130_fd_sc_hd__dfxtp_1 _2400_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b54_m12),
    .Q(pp_row66_27));
 sky130_fd_sc_hd__dfxtp_1 _2401_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b56_m10),
    .Q(pp_row66_28));
 sky130_fd_sc_hd__dfxtp_1 _2402_ (.CLK(clknet_leaf_99_clk),
    .D(booth_b58_m8),
    .Q(pp_row66_29));
 sky130_fd_sc_hd__dfxtp_1 _2403_ (.CLK(clknet_leaf_127_clk),
    .D(booth_b60_m51),
    .Q(pp_row111_7));
 sky130_fd_sc_hd__dfxtp_1 _2404_ (.CLK(clknet_leaf_99_clk),
    .D(booth_b60_m6),
    .Q(pp_row66_30));
 sky130_fd_sc_hd__dfxtp_1 _2405_ (.CLK(clknet_leaf_99_clk),
    .D(booth_b62_m4),
    .Q(pp_row66_31));
 sky130_fd_sc_hd__dfxtp_1 _2406_ (.CLK(clknet_leaf_99_clk),
    .D(booth_b64_m2),
    .Q(pp_row66_32));
 sky130_fd_sc_hd__dfxtp_2 _2407_ (.CLK(clknet_leaf_198_clk),
    .D(net219),
    .Q(pp_row66_33));
 sky130_fd_sc_hd__dfxtp_1 _2408_ (.CLK(clknet_leaf_84_clk),
    .D(notsign),
    .Q(pp_row67_0));
 sky130_fd_sc_hd__dfxtp_1 _2409_ (.CLK(clknet_leaf_84_clk),
    .D(\notsign$4544 ),
    .Q(pp_row67_1));
 sky130_fd_sc_hd__dfxtp_1 _2410_ (.CLK(clknet_leaf_84_clk),
    .D(booth_b4_m63),
    .Q(pp_row67_2));
 sky130_fd_sc_hd__dfxtp_1 _2411_ (.CLK(clknet_leaf_77_clk),
    .D(booth_b6_m61),
    .Q(pp_row67_3));
 sky130_fd_sc_hd__dfxtp_1 _2412_ (.CLK(clknet_leaf_84_clk),
    .D(booth_b8_m59),
    .Q(pp_row67_4));
 sky130_fd_sc_hd__dfxtp_1 _2413_ (.CLK(clknet_leaf_84_clk),
    .D(booth_b10_m57),
    .Q(pp_row67_5));
 sky130_fd_sc_hd__dfxtp_1 _2414_ (.CLK(clknet_leaf_127_clk),
    .D(booth_b62_m49),
    .Q(pp_row111_8));
 sky130_fd_sc_hd__dfxtp_1 _2415_ (.CLK(clknet_leaf_92_clk),
    .D(booth_b12_m55),
    .Q(pp_row67_6));
 sky130_fd_sc_hd__dfxtp_1 _2416_ (.CLK(clknet_leaf_92_clk),
    .D(booth_b14_m53),
    .Q(pp_row67_7));
 sky130_fd_sc_hd__dfxtp_1 _2417_ (.CLK(clknet_leaf_92_clk),
    .D(booth_b16_m51),
    .Q(pp_row67_8));
 sky130_fd_sc_hd__dfxtp_1 _2418_ (.CLK(clknet_leaf_145_clk),
    .D(booth_b18_m49),
    .Q(pp_row67_9));
 sky130_fd_sc_hd__dfxtp_1 _2419_ (.CLK(clknet_leaf_145_clk),
    .D(booth_b20_m47),
    .Q(pp_row67_10));
 sky130_fd_sc_hd__dfxtp_1 _2420_ (.CLK(clknet_leaf_145_clk),
    .D(booth_b22_m45),
    .Q(pp_row67_11));
 sky130_fd_sc_hd__dfxtp_1 _2421_ (.CLK(clknet_leaf_142_clk),
    .D(booth_b24_m43),
    .Q(pp_row67_12));
 sky130_fd_sc_hd__dfxtp_1 _2422_ (.CLK(clknet_leaf_142_clk),
    .D(booth_b26_m41),
    .Q(pp_row67_13));
 sky130_fd_sc_hd__dfxtp_1 _2423_ (.CLK(clknet_leaf_142_clk),
    .D(booth_b28_m39),
    .Q(pp_row67_14));
 sky130_fd_sc_hd__dfxtp_1 _2424_ (.CLK(clknet_leaf_98_clk),
    .D(booth_b30_m37),
    .Q(pp_row67_15));
 sky130_fd_sc_hd__dfxtp_1 _2425_ (.CLK(clknet_leaf_124_clk),
    .D(booth_b64_m47),
    .Q(pp_row111_9));
 sky130_fd_sc_hd__dfxtp_1 _2426_ (.CLK(clknet_leaf_98_clk),
    .D(booth_b32_m35),
    .Q(pp_row67_16));
 sky130_fd_sc_hd__dfxtp_1 _2427_ (.CLK(clknet_leaf_98_clk),
    .D(booth_b34_m33),
    .Q(pp_row67_17));
 sky130_fd_sc_hd__dfxtp_1 _2428_ (.CLK(clknet_leaf_96_clk),
    .D(booth_b36_m31),
    .Q(pp_row67_18));
 sky130_fd_sc_hd__dfxtp_1 _2429_ (.CLK(clknet_leaf_96_clk),
    .D(booth_b38_m29),
    .Q(pp_row67_19));
 sky130_fd_sc_hd__dfxtp_1 _2430_ (.CLK(clknet_leaf_96_clk),
    .D(booth_b40_m27),
    .Q(pp_row67_20));
 sky130_fd_sc_hd__dfxtp_1 _2431_ (.CLK(clknet_leaf_96_clk),
    .D(booth_b42_m25),
    .Q(pp_row67_21));
 sky130_fd_sc_hd__dfxtp_1 _2432_ (.CLK(clknet_leaf_96_clk),
    .D(booth_b44_m23),
    .Q(pp_row67_22));
 sky130_fd_sc_hd__dfxtp_1 _2433_ (.CLK(clknet_leaf_96_clk),
    .D(booth_b46_m21),
    .Q(pp_row67_23));
 sky130_fd_sc_hd__dfxtp_1 _2434_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b48_m19),
    .Q(pp_row67_24));
 sky130_fd_sc_hd__dfxtp_1 _2435_ (.CLK(clknet_leaf_75_clk),
    .D(booth_b50_m17),
    .Q(pp_row67_25));
 sky130_fd_sc_hd__dfxtp_2 _2436_ (.CLK(clknet_leaf_184_clk),
    .D(net142),
    .Q(pp_row111_10));
 sky130_fd_sc_hd__dfxtp_1 _2437_ (.CLK(clknet_leaf_74_clk),
    .D(booth_b52_m15),
    .Q(pp_row67_26));
 sky130_fd_sc_hd__dfxtp_1 _2438_ (.CLK(clknet_leaf_75_clk),
    .D(booth_b54_m13),
    .Q(pp_row67_27));
 sky130_fd_sc_hd__dfxtp_1 _2439_ (.CLK(clknet_leaf_75_clk),
    .D(booth_b56_m11),
    .Q(pp_row67_28));
 sky130_fd_sc_hd__dfxtp_1 _2440_ (.CLK(clknet_leaf_75_clk),
    .D(booth_b58_m9),
    .Q(pp_row67_29));
 sky130_fd_sc_hd__dfxtp_1 _2441_ (.CLK(clknet_leaf_98_clk),
    .D(booth_b60_m7),
    .Q(pp_row67_30));
 sky130_fd_sc_hd__dfxtp_1 _2442_ (.CLK(clknet_leaf_98_clk),
    .D(booth_b62_m5),
    .Q(pp_row67_31));
 sky130_fd_sc_hd__dfxtp_1 _2443_ (.CLK(clknet_leaf_97_clk),
    .D(booth_b64_m3),
    .Q(pp_row67_32));
 sky130_fd_sc_hd__dfxtp_2 _2444_ (.CLK(clknet_leaf_198_clk),
    .D(net220),
    .Q(pp_row67_33));
 sky130_fd_sc_hd__dfxtp_1 _2445_ (.CLK(clknet_leaf_89_clk),
    .D(booth_b4_m64),
    .Q(pp_row68_1));
 sky130_fd_sc_hd__dfxtp_1 _2446_ (.CLK(clknet_leaf_90_clk),
    .D(booth_b6_m62),
    .Q(pp_row68_2));
 sky130_fd_sc_hd__dfxtp_1 _2447_ (.CLK(clknet_leaf_128_clk),
    .D(booth_b48_m64),
    .Q(pp_row112_1));
 sky130_fd_sc_hd__dfxtp_1 _2448_ (.CLK(clknet_leaf_91_clk),
    .D(booth_b8_m60),
    .Q(pp_row68_3));
 sky130_fd_sc_hd__dfxtp_1 _2449_ (.CLK(clknet_leaf_91_clk),
    .D(booth_b10_m58),
    .Q(pp_row68_4));
 sky130_fd_sc_hd__dfxtp_1 _2450_ (.CLK(clknet_leaf_91_clk),
    .D(booth_b12_m56),
    .Q(pp_row68_5));
 sky130_fd_sc_hd__dfxtp_1 _2451_ (.CLK(clknet_leaf_92_clk),
    .D(booth_b14_m54),
    .Q(pp_row68_6));
 sky130_fd_sc_hd__dfxtp_1 _2452_ (.CLK(clknet_leaf_92_clk),
    .D(booth_b16_m52),
    .Q(pp_row68_7));
 sky130_fd_sc_hd__dfxtp_1 _2453_ (.CLK(clknet_leaf_92_clk),
    .D(booth_b18_m50),
    .Q(pp_row68_8));
 sky130_fd_sc_hd__dfxtp_1 _2454_ (.CLK(clknet_leaf_141_clk),
    .D(booth_b20_m48),
    .Q(pp_row68_9));
 sky130_fd_sc_hd__dfxtp_1 _2455_ (.CLK(clknet_leaf_92_clk),
    .D(booth_b22_m46),
    .Q(pp_row68_10));
 sky130_fd_sc_hd__dfxtp_1 _2456_ (.CLK(clknet_leaf_92_clk),
    .D(booth_b24_m44),
    .Q(pp_row68_11));
 sky130_fd_sc_hd__dfxtp_1 _2457_ (.CLK(clknet_leaf_145_clk),
    .D(booth_b26_m42),
    .Q(pp_row68_12));
 sky130_fd_sc_hd__dfxtp_1 _2458_ (.CLK(clknet_leaf_128_clk),
    .D(booth_b50_m62),
    .Q(pp_row112_2));
 sky130_fd_sc_hd__dfxtp_1 _2459_ (.CLK(clknet_leaf_148_clk),
    .D(booth_b28_m40),
    .Q(pp_row68_13));
 sky130_fd_sc_hd__dfxtp_1 _2460_ (.CLK(clknet_leaf_148_clk),
    .D(booth_b30_m38),
    .Q(pp_row68_14));
 sky130_fd_sc_hd__dfxtp_1 _2461_ (.CLK(clknet_leaf_95_clk),
    .D(booth_b32_m36),
    .Q(pp_row68_15));
 sky130_fd_sc_hd__dfxtp_1 _2462_ (.CLK(clknet_leaf_95_clk),
    .D(booth_b34_m34),
    .Q(pp_row68_16));
 sky130_fd_sc_hd__dfxtp_1 _2463_ (.CLK(clknet_leaf_94_clk),
    .D(booth_b36_m32),
    .Q(pp_row68_17));
 sky130_fd_sc_hd__dfxtp_1 _2464_ (.CLK(clknet_leaf_94_clk),
    .D(booth_b38_m30),
    .Q(pp_row68_18));
 sky130_fd_sc_hd__dfxtp_1 _2465_ (.CLK(clknet_leaf_95_clk),
    .D(booth_b40_m28),
    .Q(pp_row68_19));
 sky130_fd_sc_hd__dfxtp_1 _2466_ (.CLK(clknet_leaf_95_clk),
    .D(booth_b42_m26),
    .Q(pp_row68_20));
 sky130_fd_sc_hd__dfxtp_1 _2467_ (.CLK(clknet_leaf_95_clk),
    .D(booth_b44_m24),
    .Q(pp_row68_21));
 sky130_fd_sc_hd__dfxtp_1 _2468_ (.CLK(clknet_leaf_102_clk),
    .D(booth_b46_m22),
    .Q(pp_row68_22));
 sky130_fd_sc_hd__dfxtp_1 _2469_ (.CLK(clknet_leaf_124_clk),
    .D(booth_b52_m60),
    .Q(pp_row112_3));
 sky130_fd_sc_hd__dfxtp_1 _2470_ (.CLK(clknet_leaf_98_clk),
    .D(booth_b48_m20),
    .Q(pp_row68_23));
 sky130_fd_sc_hd__dfxtp_1 _2471_ (.CLK(clknet_leaf_98_clk),
    .D(booth_b50_m18),
    .Q(pp_row68_24));
 sky130_fd_sc_hd__dfxtp_1 _2472_ (.CLK(clknet_leaf_98_clk),
    .D(booth_b52_m16),
    .Q(pp_row68_25));
 sky130_fd_sc_hd__dfxtp_1 _2473_ (.CLK(clknet_leaf_98_clk),
    .D(booth_b54_m14),
    .Q(pp_row68_26));
 sky130_fd_sc_hd__dfxtp_1 _2474_ (.CLK(clknet_leaf_99_clk),
    .D(booth_b56_m12),
    .Q(pp_row68_27));
 sky130_fd_sc_hd__dfxtp_1 _2475_ (.CLK(clknet_leaf_99_clk),
    .D(booth_b58_m10),
    .Q(pp_row68_28));
 sky130_fd_sc_hd__dfxtp_1 _2476_ (.CLK(clknet_leaf_99_clk),
    .D(booth_b60_m8),
    .Q(pp_row68_29));
 sky130_fd_sc_hd__dfxtp_1 _2477_ (.CLK(clknet_leaf_99_clk),
    .D(booth_b62_m6),
    .Q(pp_row68_30));
 sky130_fd_sc_hd__dfxtp_1 _2478_ (.CLK(clknet_leaf_99_clk),
    .D(booth_b64_m4),
    .Q(pp_row68_31));
 sky130_fd_sc_hd__dfxtp_2 _2479_ (.CLK(clknet_leaf_198_clk),
    .D(net221),
    .Q(pp_row68_32));
 sky130_fd_sc_hd__dfxtp_1 _2480_ (.CLK(clknet_leaf_125_clk),
    .D(booth_b54_m58),
    .Q(pp_row112_4));
 sky130_fd_sc_hd__dfxtp_1 _2481_ (.CLK(clknet_leaf_147_clk),
    .D(\notsign$4614 ),
    .Q(pp_row69_0));
 sky130_fd_sc_hd__dfxtp_1 _2482_ (.CLK(clknet_leaf_142_clk),
    .D(booth_b6_m63),
    .Q(pp_row69_1));
 sky130_fd_sc_hd__dfxtp_1 _2483_ (.CLK(clknet_leaf_147_clk),
    .D(booth_b8_m61),
    .Q(pp_row69_2));
 sky130_fd_sc_hd__dfxtp_1 _2484_ (.CLK(clknet_leaf_146_clk),
    .D(booth_b10_m59),
    .Q(pp_row69_3));
 sky130_fd_sc_hd__dfxtp_1 _2485_ (.CLK(clknet_leaf_146_clk),
    .D(booth_b12_m57),
    .Q(pp_row69_4));
 sky130_fd_sc_hd__dfxtp_1 _2486_ (.CLK(clknet_leaf_146_clk),
    .D(booth_b14_m55),
    .Q(pp_row69_5));
 sky130_fd_sc_hd__dfxtp_1 _2487_ (.CLK(clknet_leaf_90_clk),
    .D(booth_b16_m53),
    .Q(pp_row69_6));
 sky130_fd_sc_hd__dfxtp_1 _2488_ (.CLK(clknet_leaf_90_clk),
    .D(booth_b18_m51),
    .Q(pp_row69_7));
 sky130_fd_sc_hd__dfxtp_1 _2489_ (.CLK(clknet_leaf_90_clk),
    .D(booth_b20_m49),
    .Q(pp_row69_8));
 sky130_fd_sc_hd__dfxtp_1 _2490_ (.CLK(clknet_leaf_90_clk),
    .D(booth_b22_m47),
    .Q(pp_row69_9));
 sky130_fd_sc_hd__dfxtp_1 _2491_ (.CLK(clknet_leaf_125_clk),
    .D(booth_b56_m56),
    .Q(pp_row112_5));
 sky130_fd_sc_hd__dfxtp_1 _2492_ (.CLK(clknet_leaf_90_clk),
    .D(booth_b24_m45),
    .Q(pp_row69_10));
 sky130_fd_sc_hd__dfxtp_1 _2493_ (.CLK(clknet_leaf_90_clk),
    .D(booth_b26_m43),
    .Q(pp_row69_11));
 sky130_fd_sc_hd__dfxtp_1 _2494_ (.CLK(clknet_leaf_142_clk),
    .D(booth_b28_m41),
    .Q(pp_row69_12));
 sky130_fd_sc_hd__dfxtp_1 _2495_ (.CLK(clknet_leaf_142_clk),
    .D(booth_b30_m39),
    .Q(pp_row69_13));
 sky130_fd_sc_hd__dfxtp_1 _2496_ (.CLK(clknet_leaf_141_clk),
    .D(booth_b32_m37),
    .Q(pp_row69_14));
 sky130_fd_sc_hd__dfxtp_1 _2497_ (.CLK(clknet_leaf_97_clk),
    .D(booth_b34_m35),
    .Q(pp_row69_15));
 sky130_fd_sc_hd__dfxtp_1 _2498_ (.CLK(clknet_leaf_97_clk),
    .D(booth_b36_m33),
    .Q(pp_row69_16));
 sky130_fd_sc_hd__dfxtp_1 _2499_ (.CLK(clknet_leaf_97_clk),
    .D(booth_b38_m31),
    .Q(pp_row69_17));
 sky130_fd_sc_hd__dfxtp_1 _2500_ (.CLK(clknet_leaf_147_clk),
    .D(booth_b40_m29),
    .Q(pp_row69_18));
 sky130_fd_sc_hd__dfxtp_1 _2501_ (.CLK(clknet_leaf_147_clk),
    .D(booth_b42_m27),
    .Q(pp_row69_19));
 sky130_fd_sc_hd__dfxtp_1 _2502_ (.CLK(clknet_leaf_125_clk),
    .D(booth_b58_m54),
    .Q(pp_row112_6));
 sky130_fd_sc_hd__dfxtp_1 _2503_ (.CLK(clknet_leaf_179_clk),
    .D(booth_b62_m63),
    .Q(pp_row125_1));
 sky130_fd_sc_hd__conb_1 dadda_fa_0_70_0_1892 (.HI(net1892));
 sky130_fd_sc_hd__conb_1 dadda_fa_0_72_0_1893 (.HI(net1893));
 sky130_fd_sc_hd__conb_1 dadda_fa_0_74_0_1894 (.HI(net1894));
 sky130_fd_sc_hd__conb_1 dadda_fa_0_76_0_1895 (.HI(net1895));
 sky130_fd_sc_hd__conb_1 dadda_fa_1_80_0_1896 (.HI(net1896));
 sky130_fd_sc_hd__conb_1 dadda_fa_1_82_0_1897 (.HI(net1897));
 sky130_fd_sc_hd__conb_1 dadda_fa_1_84_0_1898 (.HI(net1898));
 sky130_fd_sc_hd__conb_1 dadda_fa_1_86_0_1899 (.HI(net1899));
 sky130_fd_sc_hd__conb_1 dadda_fa_1_88_0_1900 (.HI(net1900));
 sky130_fd_sc_hd__conb_1 dadda_fa_1_90_0_1901 (.HI(net1901));
 sky130_fd_sc_hd__conb_1 dadda_fa_1_92_0_1902 (.HI(net1902));
 sky130_fd_sc_hd__conb_1 dadda_fa_1_94_0_1903 (.HI(net1903));
 sky130_fd_sc_hd__conb_1 dadda_fa_2_100_0_1904 (.HI(net1904));
 sky130_fd_sc_hd__conb_1 dadda_fa_2_102_0_1905 (.HI(net1905));
 sky130_fd_sc_hd__conb_1 dadda_fa_2_104_0_1906 (.HI(net1906));
 sky130_fd_sc_hd__conb_1 dadda_fa_2_106_0_1907 (.HI(net1907));
 sky130_fd_sc_hd__conb_1 dadda_fa_2_98_0_1908 (.HI(net1908));
 sky130_fd_sc_hd__conb_1 dadda_fa_3_110_0_1909 (.HI(net1909));
 sky130_fd_sc_hd__conb_1 dadda_fa_3_112_0_1910 (.HI(net1910));
 sky130_fd_sc_hd__conb_1 dadda_fa_3_114_0_1911 (.HI(net1911));
 sky130_fd_sc_hd__conb_1 dadda_fa_4_118_0_1912 (.HI(net1912));
 sky130_fd_sc_hd__conb_1 dadda_fa_4_120_0_1913 (.HI(net1913));
 sky130_fd_sc_hd__conb_1 dadda_fa_5_124_0_1914 (.HI(net1914));
 sky130_fd_sc_hd__conb_1 dadda_ha_0_78_0_1915 (.HI(net1915));
 sky130_fd_sc_hd__conb_1 dadda_ha_1_96_0_1916 (.HI(net1916));
 sky130_fd_sc_hd__conb_1 dadda_ha_2_108_0_1917 (.HI(net1917));
 sky130_fd_sc_hd__conb_1 dadda_ha_3_116_0_1918 (.HI(net1918));
 sky130_fd_sc_hd__conb_1 dadda_ha_4_122_0_1919 (.HI(net1919));
 sky130_fd_sc_hd__conb_1 dadda_ha_5_126_0_1920 (.HI(net1920));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__conb_1 \U$$1093_1754  (.LO(net1754));
 sky130_fd_sc_hd__conb_1 \U$$1102_1755  (.LO(net1755));
 sky130_fd_sc_hd__conb_1 \U$$1230_1756  (.LO(net1756));
 sky130_fd_sc_hd__conb_1 \U$$1239_1757  (.LO(net1757));
 sky130_fd_sc_hd__conb_1 \U$$134_1758  (.LO(net1758));
 sky130_fd_sc_hd__conb_1 \U$$1367_1759  (.LO(net1759));
 sky130_fd_sc_hd__conb_1 \U$$1376_1760  (.LO(net1760));
 sky130_fd_sc_hd__conb_1 \U$$143_1761  (.LO(net1761));
 sky130_fd_sc_hd__conb_1 \U$$1504_1762  (.LO(net1762));
 sky130_fd_sc_hd__conb_1 \U$$1513_1763  (.LO(net1763));
 sky130_fd_sc_hd__conb_1 \U$$1641_1764  (.LO(net1764));
 sky130_fd_sc_hd__conb_1 \U$$1650_1765  (.LO(net1765));
 sky130_fd_sc_hd__conb_1 \U$$1778_1766  (.LO(net1766));
 sky130_fd_sc_hd__conb_1 \U$$1787_1767  (.LO(net1767));
 sky130_fd_sc_hd__conb_1 \U$$1915_1768  (.LO(net1768));
 sky130_fd_sc_hd__conb_1 \U$$1924_1769  (.LO(net1769));
 sky130_fd_sc_hd__conb_1 \U$$2052_1770  (.LO(net1770));
 sky130_fd_sc_hd__conb_1 \U$$2061_1771  (.LO(net1771));
 sky130_fd_sc_hd__conb_1 \U$$2189_1772  (.LO(net1772));
 sky130_fd_sc_hd__conb_1 \U$$2198_1773  (.LO(net1773));
 sky130_fd_sc_hd__conb_1 \U$$2326_1774  (.LO(net1774));
 sky130_fd_sc_hd__conb_1 \U$$2335_1775  (.LO(net1775));
 sky130_fd_sc_hd__conb_1 \U$$2463_1776  (.LO(net1776));
 sky130_fd_sc_hd__conb_1 \U$$2472_1777  (.LO(net1777));
 sky130_fd_sc_hd__conb_1 \U$$2600_1778  (.LO(net1778));
 sky130_fd_sc_hd__conb_1 \U$$2609_1779  (.LO(net1779));
 sky130_fd_sc_hd__conb_1 \U$$271_1780  (.LO(net1780));
 sky130_fd_sc_hd__conb_1 \U$$2737_1781  (.LO(net1781));
 sky130_fd_sc_hd__conb_1 \U$$2746_1782  (.LO(net1782));
 sky130_fd_sc_hd__conb_1 \U$$280_1783  (.LO(net1783));
 sky130_fd_sc_hd__conb_1 \U$$2874_1784  (.LO(net1784));
 sky130_fd_sc_hd__conb_1 \U$$2883_1785  (.LO(net1785));
 sky130_fd_sc_hd__conb_1 \U$$3011_1786  (.LO(net1786));
 sky130_fd_sc_hd__conb_1 \U$$3020_1787  (.LO(net1787));
 sky130_fd_sc_hd__conb_1 \U$$3148_1788  (.LO(net1788));
 sky130_fd_sc_hd__conb_1 \U$$3157_1789  (.LO(net1789));
 sky130_fd_sc_hd__conb_1 \U$$3285_1790  (.LO(net1790));
 sky130_fd_sc_hd__conb_1 \U$$3294_1791  (.LO(net1791));
 sky130_fd_sc_hd__conb_1 \U$$3422_1792  (.LO(net1792));
 sky130_fd_sc_hd__conb_1 \U$$3431_1793  (.LO(net1793));
 sky130_fd_sc_hd__conb_1 \U$$3559_1794  (.LO(net1794));
 sky130_fd_sc_hd__conb_1 \U$$3568_1795  (.LO(net1795));
 sky130_fd_sc_hd__conb_1 \U$$3696_1796  (.LO(net1796));
 sky130_fd_sc_hd__conb_1 \U$$3705_1797  (.LO(net1797));
 sky130_fd_sc_hd__conb_1 \U$$3833_1798  (.LO(net1798));
 sky130_fd_sc_hd__conb_1 \U$$3842_1799  (.LO(net1799));
 sky130_fd_sc_hd__conb_1 \U$$3970_1800  (.LO(net1800));
 sky130_fd_sc_hd__conb_1 \U$$3979_1801  (.LO(net1801));
 sky130_fd_sc_hd__conb_1 \U$$4_1802  (.LO(net1802));
 sky130_fd_sc_hd__conb_1 \U$$408_1803  (.LO(net1803));
 sky130_fd_sc_hd__conb_1 \U$$4107_1804  (.LO(net1804));
 sky130_fd_sc_hd__conb_1 \U$$4116_1805  (.LO(net1805));
 sky130_fd_sc_hd__conb_1 \U$$417_1806  (.LO(net1806));
 sky130_fd_sc_hd__conb_1 \U$$4244_1807  (.LO(net1807));
 sky130_fd_sc_hd__conb_1 \U$$4253_1808  (.LO(net1808));
 sky130_fd_sc_hd__conb_1 \U$$4381_1809  (.LO(net1809));
 sky130_fd_sc_hd__conb_1 \U$$4385_1810  (.LO(net1810));
 sky130_fd_sc_hd__conb_1 \U$$4386_1811  (.LO(net1811));
 sky130_fd_sc_hd__conb_1 \U$$4387_1812  (.LO(net1812));
 sky130_fd_sc_hd__conb_1 \U$$4388_1813  (.LO(net1813));
 sky130_fd_sc_hd__conb_1 \U$$4389_1814  (.LO(net1814));
 sky130_fd_sc_hd__conb_1 \U$$4390_1815  (.LO(net1815));
 sky130_fd_sc_hd__conb_1 \U$$4391_1816  (.LO(net1816));
 sky130_fd_sc_hd__conb_1 \U$$4393_1817  (.LO(net1817));
 sky130_fd_sc_hd__conb_1 \U$$4395_1818  (.LO(net1818));
 sky130_fd_sc_hd__conb_1 \U$$4397_1819  (.LO(net1819));
 sky130_fd_sc_hd__conb_1 \U$$4399_1820  (.LO(net1820));
 sky130_fd_sc_hd__conb_1 \U$$4401_1821  (.LO(net1821));
 sky130_fd_sc_hd__conb_1 \U$$4403_1822  (.LO(net1822));
 sky130_fd_sc_hd__conb_1 \U$$4405_1823  (.LO(net1823));
 sky130_fd_sc_hd__conb_1 \U$$4407_1824  (.LO(net1824));
 sky130_fd_sc_hd__conb_1 \U$$4409_1825  (.LO(net1825));
 sky130_fd_sc_hd__conb_1 \U$$4411_1826  (.LO(net1826));
 sky130_fd_sc_hd__conb_1 \U$$4413_1827  (.LO(net1827));
 sky130_fd_sc_hd__conb_1 \U$$4415_1828  (.LO(net1828));
 sky130_fd_sc_hd__conb_1 \U$$4417_1829  (.LO(net1829));
 sky130_fd_sc_hd__conb_1 \U$$4419_1830  (.LO(net1830));
 sky130_fd_sc_hd__conb_1 \U$$4421_1831  (.LO(net1831));
 sky130_fd_sc_hd__conb_1 \U$$4423_1832  (.LO(net1832));
 sky130_fd_sc_hd__conb_1 \U$$4425_1833  (.LO(net1833));
 sky130_fd_sc_hd__conb_1 \U$$4427_1834  (.LO(net1834));
 sky130_fd_sc_hd__conb_1 \U$$4429_1835  (.LO(net1835));
 sky130_fd_sc_hd__conb_1 \U$$4431_1836  (.LO(net1836));
 sky130_fd_sc_hd__conb_1 \U$$4433_1837  (.LO(net1837));
 sky130_fd_sc_hd__conb_1 \U$$4435_1838  (.LO(net1838));
 sky130_fd_sc_hd__conb_1 \U$$4437_1839  (.LO(net1839));
 sky130_fd_sc_hd__conb_1 \U$$4439_1840  (.LO(net1840));
 sky130_fd_sc_hd__conb_1 \U$$4441_1841  (.LO(net1841));
 sky130_fd_sc_hd__conb_1 \U$$4443_1842  (.LO(net1842));
 sky130_fd_sc_hd__conb_1 \U$$4445_1843  (.LO(net1843));
 sky130_fd_sc_hd__conb_1 \U$$4447_1844  (.LO(net1844));
 sky130_fd_sc_hd__conb_1 \U$$4449_1845  (.LO(net1845));
 sky130_fd_sc_hd__conb_1 \U$$4451_1846  (.LO(net1846));
 sky130_fd_sc_hd__conb_1 \U$$4453_1847  (.LO(net1847));
 sky130_fd_sc_hd__conb_1 \U$$4455_1848  (.LO(net1848));
 sky130_fd_sc_hd__conb_1 \U$$4457_1849  (.LO(net1849));
 sky130_fd_sc_hd__conb_1 \U$$4459_1850  (.LO(net1850));
 sky130_fd_sc_hd__conb_1 \U$$4461_1851  (.LO(net1851));
 sky130_fd_sc_hd__conb_1 \U$$4463_1852  (.LO(net1852));
 sky130_fd_sc_hd__conb_1 \U$$4465_1853  (.LO(net1853));
 sky130_fd_sc_hd__conb_1 \U$$4467_1854  (.LO(net1854));
 sky130_fd_sc_hd__conb_1 \U$$4469_1855  (.LO(net1855));
 sky130_fd_sc_hd__conb_1 \U$$4471_1856  (.LO(net1856));
 sky130_fd_sc_hd__conb_1 \U$$4473_1857  (.LO(net1857));
 sky130_fd_sc_hd__conb_1 \U$$4475_1858  (.LO(net1858));
 sky130_fd_sc_hd__conb_1 \U$$4477_1859  (.LO(net1859));
 sky130_fd_sc_hd__conb_1 \U$$4479_1860  (.LO(net1860));
 sky130_fd_sc_hd__conb_1 \U$$4481_1861  (.LO(net1861));
 sky130_fd_sc_hd__conb_1 \U$$4483_1862  (.LO(net1862));
 sky130_fd_sc_hd__conb_1 \U$$4485_1863  (.LO(net1863));
 sky130_fd_sc_hd__conb_1 \U$$4487_1864  (.LO(net1864));
 sky130_fd_sc_hd__conb_1 \U$$4489_1865  (.LO(net1865));
 sky130_fd_sc_hd__conb_1 \U$$4491_1866  (.LO(net1866));
 sky130_fd_sc_hd__conb_1 \U$$4493_1867  (.LO(net1867));
 sky130_fd_sc_hd__conb_1 \U$$4495_1868  (.LO(net1868));
 sky130_fd_sc_hd__conb_1 \U$$4497_1869  (.LO(net1869));
 sky130_fd_sc_hd__conb_1 \U$$4499_1870  (.LO(net1870));
 sky130_fd_sc_hd__conb_1 \U$$4501_1871  (.LO(net1871));
 sky130_fd_sc_hd__conb_1 \U$$4503_1872  (.LO(net1872));
 sky130_fd_sc_hd__conb_1 \U$$4505_1873  (.LO(net1873));
 sky130_fd_sc_hd__conb_1 \U$$4507_1874  (.LO(net1874));
 sky130_fd_sc_hd__conb_1 \U$$4509_1875  (.LO(net1875));
 sky130_fd_sc_hd__conb_1 \U$$4511_1876  (.LO(net1876));
 sky130_fd_sc_hd__conb_1 \U$$4513_1877  (.LO(net1877));
 sky130_fd_sc_hd__conb_1 \U$$4515_1878  (.LO(net1878));
 sky130_fd_sc_hd__conb_1 \U$$4517_1879  (.LO(net1879));
 sky130_fd_sc_hd__conb_1 \U$$5_1880  (.LO(net1880));
 sky130_fd_sc_hd__conb_1 \U$$545_1881  (.LO(net1881));
 sky130_fd_sc_hd__conb_1 \U$$554_1882  (.LO(net1882));
 sky130_fd_sc_hd__conb_1 \U$$6_1883  (.LO(net1883));
 sky130_fd_sc_hd__conb_1 \U$$682_1884  (.LO(net1884));
 sky130_fd_sc_hd__conb_1 \U$$691_1885  (.LO(net1885));
 sky130_fd_sc_hd__conb_1 \U$$819_1886  (.LO(net1886));
 sky130_fd_sc_hd__conb_1 \U$$828_1887  (.LO(net1887));
 sky130_fd_sc_hd__conb_1 \U$$956_1888  (.LO(net1888));
 sky130_fd_sc_hd__conb_1 \U$$965_1889  (.LO(net1889));
 sky130_fd_sc_hd__conb_1 \final_adder.U$$961_1890  (.LO(net1890));
 sky130_fd_sc_hd__conb_1 dadda_fa_0_68_0_1891 (.HI(net1891));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_54_0 (.A(pp_row54_0),
    .B(pp_row54_1),
    .CIN(pp_row54_2),
    .COUT(\c$4 ),
    .SUM(\s$5 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_55_0 (.A(pp_row55_0),
    .B(pp_row55_1),
    .CIN(pp_row55_2),
    .COUT(\c$8 ),
    .SUM(\s$9 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_56_0 (.A(pp_row56_0),
    .B(pp_row56_1),
    .CIN(pp_row56_2),
    .COUT(\c$12 ),
    .SUM(\s$13 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_56_1 (.A(pp_row56_3),
    .B(pp_row56_4),
    .CIN(pp_row56_5),
    .COUT(\c$14 ),
    .SUM(\s$15 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_57_0 (.A(pp_row57_0),
    .B(pp_row57_1),
    .CIN(pp_row57_2),
    .COUT(\c$18 ),
    .SUM(\s$19 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_57_1 (.A(pp_row57_3),
    .B(pp_row57_4),
    .CIN(pp_row57_5),
    .COUT(\c$20 ),
    .SUM(\s$21 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_58_0 (.A(pp_row58_0),
    .B(pp_row58_1),
    .CIN(pp_row58_2),
    .COUT(\c$24 ),
    .SUM(\s$25 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_58_1 (.A(pp_row58_3),
    .B(pp_row58_4),
    .CIN(pp_row58_5),
    .COUT(\c$26 ),
    .SUM(\s$27 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_58_2 (.A(pp_row58_6),
    .B(pp_row58_7),
    .CIN(pp_row58_8),
    .COUT(\c$28 ),
    .SUM(\s$29 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_59_0 (.A(pp_row59_0),
    .B(pp_row59_1),
    .CIN(pp_row59_2),
    .COUT(\c$32 ),
    .SUM(\s$33 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_59_1 (.A(pp_row59_3),
    .B(pp_row59_4),
    .CIN(pp_row59_5),
    .COUT(\c$34 ),
    .SUM(\s$35 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_59_2 (.A(pp_row59_6),
    .B(pp_row59_7),
    .CIN(pp_row59_8),
    .COUT(\c$36 ),
    .SUM(\s$37 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_60_0 (.A(pp_row60_0),
    .B(pp_row60_1),
    .CIN(pp_row60_2),
    .COUT(\c$40 ),
    .SUM(\s$41 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_60_1 (.A(pp_row60_3),
    .B(pp_row60_4),
    .CIN(pp_row60_5),
    .COUT(\c$42 ),
    .SUM(\s$43 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_60_2 (.A(pp_row60_6),
    .B(pp_row60_7),
    .CIN(pp_row60_8),
    .COUT(\c$44 ),
    .SUM(\s$45 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_60_3 (.A(pp_row60_9),
    .B(pp_row60_10),
    .CIN(pp_row60_11),
    .COUT(\c$46 ),
    .SUM(\s$47 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_0_61_0 (.A(pp_row61_0),
    .B(pp_row61_1),
    .CIN(pp_row61_2),
    .COUT(\c$50 ),
    .SUM(\s$51 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_61_1 (.A(pp_row61_3),
    .B(pp_row61_4),
    .CIN(pp_row61_5),
    .COUT(\c$52 ),
    .SUM(\s$53 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_61_2 (.A(pp_row61_6),
    .B(pp_row61_7),
    .CIN(pp_row61_8),
    .COUT(\c$54 ),
    .SUM(\s$55 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_61_3 (.A(pp_row61_9),
    .B(pp_row61_10),
    .CIN(pp_row61_11),
    .COUT(\c$56 ),
    .SUM(\s$57 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_62_0 (.A(pp_row62_0),
    .B(pp_row62_1),
    .CIN(pp_row62_2),
    .COUT(\c$60 ),
    .SUM(\s$61 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_62_1 (.A(pp_row62_3),
    .B(pp_row62_4),
    .CIN(pp_row62_5),
    .COUT(\c$62 ),
    .SUM(\s$63 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_62_2 (.A(pp_row62_6),
    .B(pp_row62_7),
    .CIN(pp_row62_8),
    .COUT(\c$64 ),
    .SUM(\s$65 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_62_3 (.A(pp_row62_9),
    .B(pp_row62_10),
    .CIN(pp_row62_11),
    .COUT(\c$66 ),
    .SUM(\s$67 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_62_4 (.A(pp_row62_12),
    .B(pp_row62_13),
    .CIN(pp_row62_14),
    .COUT(\c$68 ),
    .SUM(\s$69 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_63_0 (.A(pp_row63_0),
    .B(pp_row63_1),
    .CIN(pp_row63_2),
    .COUT(\c$72 ),
    .SUM(\s$73 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_63_1 (.A(pp_row63_3),
    .B(pp_row63_4),
    .CIN(pp_row63_5),
    .COUT(\c$74 ),
    .SUM(\s$75 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_63_2 (.A(pp_row63_6),
    .B(pp_row63_7),
    .CIN(pp_row63_8),
    .COUT(\c$76 ),
    .SUM(\s$77 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_63_3 (.A(pp_row63_9),
    .B(pp_row63_10),
    .CIN(pp_row63_11),
    .COUT(\c$78 ),
    .SUM(\s$79 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_63_4 (.A(pp_row63_12),
    .B(pp_row63_13),
    .CIN(pp_row63_14),
    .COUT(\c$80 ),
    .SUM(\s$81 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_0_64_0 (.A(pp_row64_0),
    .B(pp_row64_1),
    .CIN(pp_row64_2),
    .COUT(\c$84 ),
    .SUM(\s$85 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_0_64_1 (.A(pp_row64_3),
    .B(pp_row64_4),
    .CIN(pp_row64_5),
    .COUT(\c$86 ),
    .SUM(\s$87 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_64_2 (.A(pp_row64_6),
    .B(pp_row64_7),
    .CIN(pp_row64_8),
    .COUT(\c$88 ),
    .SUM(\s$89 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_64_3 (.A(pp_row64_9),
    .B(pp_row64_10),
    .CIN(pp_row64_11),
    .COUT(\c$90 ),
    .SUM(\s$91 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_64_4 (.A(pp_row64_12),
    .B(pp_row64_13),
    .CIN(pp_row64_14),
    .COUT(\c$92 ),
    .SUM(\s$93 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_64_5 (.A(pp_row64_15),
    .B(pp_row64_16),
    .CIN(pp_row64_17),
    .COUT(\c$94 ),
    .SUM(\s$95 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_65_0 (.A(pp_row0_1),
    .B(pp_row65_1),
    .CIN(pp_row65_2),
    .COUT(\c$96 ),
    .SUM(\s$97 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_65_1 (.A(pp_row65_3),
    .B(pp_row65_4),
    .CIN(pp_row65_5),
    .COUT(\c$98 ),
    .SUM(\s$99 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_65_2 (.A(pp_row65_6),
    .B(pp_row65_7),
    .CIN(pp_row65_8),
    .COUT(\c$100 ),
    .SUM(\s$101 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_65_3 (.A(pp_row65_9),
    .B(pp_row65_10),
    .CIN(pp_row65_11),
    .COUT(\c$102 ),
    .SUM(\s$103 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_65_4 (.A(pp_row65_12),
    .B(pp_row65_13),
    .CIN(pp_row65_14),
    .COUT(\c$104 ),
    .SUM(\s$105 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_0_65_5 (.A(pp_row65_15),
    .B(pp_row65_16),
    .CIN(pp_row65_17),
    .COUT(\c$106 ),
    .SUM(\s$107 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_66_0 (.A(pp_row0_1),
    .B(pp_row66_1),
    .CIN(pp_row66_2),
    .COUT(\c$108 ),
    .SUM(\s$109 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_66_1 (.A(pp_row66_3),
    .B(pp_row66_4),
    .CIN(pp_row66_5),
    .COUT(\c$110 ),
    .SUM(\s$111 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_66_2 (.A(pp_row66_6),
    .B(pp_row66_7),
    .CIN(pp_row66_8),
    .COUT(\c$112 ),
    .SUM(\s$113 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_66_3 (.A(pp_row66_9),
    .B(pp_row66_10),
    .CIN(pp_row66_11),
    .COUT(\c$114 ),
    .SUM(\s$115 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_66_4 (.A(pp_row66_12),
    .B(pp_row66_13),
    .CIN(pp_row66_14),
    .COUT(\c$116 ),
    .SUM(\s$117 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_0_66_5 (.A(pp_row66_15),
    .B(pp_row66_16),
    .CIN(pp_row66_17),
    .COUT(\c$118 ),
    .SUM(\s$119 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_67_0 (.A(pp_row67_0),
    .B(pp_row67_1),
    .CIN(pp_row67_2),
    .COUT(\c$120 ),
    .SUM(\s$121 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_67_1 (.A(pp_row67_3),
    .B(pp_row67_4),
    .CIN(pp_row67_5),
    .COUT(\c$122 ),
    .SUM(\s$123 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_67_2 (.A(pp_row67_6),
    .B(pp_row67_7),
    .CIN(pp_row67_8),
    .COUT(\c$124 ),
    .SUM(\s$125 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_0_67_3 (.A(pp_row67_9),
    .B(pp_row67_10),
    .CIN(pp_row67_11),
    .COUT(\c$126 ),
    .SUM(\s$127 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_67_4 (.A(pp_row67_12),
    .B(pp_row67_13),
    .CIN(pp_row67_14),
    .COUT(\c$128 ),
    .SUM(\s$129 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_0_67_5 (.A(pp_row67_15),
    .B(pp_row67_16),
    .CIN(pp_row67_17),
    .COUT(\c$130 ),
    .SUM(\s$131 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_68_0 (.A(net1891),
    .B(pp_row68_1),
    .CIN(pp_row68_2),
    .COUT(\c$132 ),
    .SUM(\s$133 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_68_1 (.A(pp_row68_3),
    .B(pp_row68_4),
    .CIN(pp_row68_5),
    .COUT(\c$134 ),
    .SUM(\s$135 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_68_2 (.A(pp_row68_6),
    .B(pp_row68_7),
    .CIN(pp_row68_8),
    .COUT(\c$136 ),
    .SUM(\s$137 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_68_3 (.A(pp_row68_9),
    .B(pp_row68_10),
    .CIN(pp_row68_11),
    .COUT(\c$138 ),
    .SUM(\s$139 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_68_4 (.A(pp_row68_12),
    .B(pp_row68_13),
    .CIN(pp_row68_14),
    .COUT(\c$140 ),
    .SUM(\s$141 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_69_0 (.A(pp_row69_0),
    .B(pp_row69_1),
    .CIN(pp_row69_2),
    .COUT(\c$144 ),
    .SUM(\s$145 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_69_1 (.A(pp_row69_3),
    .B(pp_row69_4),
    .CIN(pp_row69_5),
    .COUT(\c$146 ),
    .SUM(\s$147 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_69_2 (.A(pp_row69_6),
    .B(pp_row69_7),
    .CIN(pp_row69_8),
    .COUT(\c$148 ),
    .SUM(\s$149 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_69_3 (.A(pp_row69_9),
    .B(pp_row69_10),
    .CIN(pp_row69_11),
    .COUT(\c$150 ),
    .SUM(\s$151 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_69_4 (.A(pp_row69_12),
    .B(pp_row69_13),
    .CIN(pp_row69_14),
    .COUT(\c$152 ),
    .SUM(\s$153 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_70_0 (.A(net1892),
    .B(pp_row70_1),
    .CIN(pp_row70_2),
    .COUT(\c$154 ),
    .SUM(\s$155 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_70_1 (.A(pp_row70_3),
    .B(pp_row70_4),
    .CIN(pp_row70_5),
    .COUT(\c$156 ),
    .SUM(\s$157 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_70_2 (.A(pp_row70_6),
    .B(pp_row70_7),
    .CIN(pp_row70_8),
    .COUT(\c$158 ),
    .SUM(\s$159 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_70_3 (.A(pp_row70_9),
    .B(pp_row70_10),
    .CIN(pp_row70_11),
    .COUT(\c$160 ),
    .SUM(\s$161 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_71_0 (.A(pp_row71_0),
    .B(pp_row71_1),
    .CIN(pp_row71_2),
    .COUT(\c$164 ),
    .SUM(\s$165 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_71_1 (.A(pp_row71_3),
    .B(pp_row71_4),
    .CIN(pp_row71_5),
    .COUT(\c$166 ),
    .SUM(\s$167 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_71_2 (.A(pp_row71_6),
    .B(pp_row71_7),
    .CIN(pp_row71_8),
    .COUT(\c$168 ),
    .SUM(\s$169 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_0_71_3 (.A(pp_row71_9),
    .B(pp_row71_10),
    .CIN(pp_row71_11),
    .COUT(\c$170 ),
    .SUM(\s$171 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_72_0 (.A(net1893),
    .B(pp_row72_1),
    .CIN(pp_row72_2),
    .COUT(\c$172 ),
    .SUM(\s$173 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_72_1 (.A(pp_row72_3),
    .B(pp_row72_4),
    .CIN(pp_row72_5),
    .COUT(\c$174 ),
    .SUM(\s$175 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_72_2 (.A(pp_row72_6),
    .B(pp_row72_7),
    .CIN(pp_row72_8),
    .COUT(\c$176 ),
    .SUM(\s$177 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_73_0 (.A(pp_row73_0),
    .B(pp_row73_1),
    .CIN(pp_row73_2),
    .COUT(\c$180 ),
    .SUM(\s$181 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_73_1 (.A(pp_row73_3),
    .B(pp_row73_4),
    .CIN(pp_row73_5),
    .COUT(\c$182 ),
    .SUM(\s$183 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_73_2 (.A(pp_row73_6),
    .B(pp_row73_7),
    .CIN(pp_row73_8),
    .COUT(\c$184 ),
    .SUM(\s$185 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_74_0 (.A(net1894),
    .B(pp_row74_1),
    .CIN(pp_row74_2),
    .COUT(\c$186 ),
    .SUM(\s$187 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_74_1 (.A(pp_row74_3),
    .B(pp_row74_4),
    .CIN(pp_row74_5),
    .COUT(\c$188 ),
    .SUM(\s$189 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_75_0 (.A(pp_row75_0),
    .B(pp_row75_1),
    .CIN(pp_row75_2),
    .COUT(\c$192 ),
    .SUM(\s$193 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_75_1 (.A(pp_row75_3),
    .B(pp_row75_4),
    .CIN(pp_row75_5),
    .COUT(\c$194 ),
    .SUM(\s$195 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_76_0 (.A(net1895),
    .B(pp_row76_1),
    .CIN(pp_row76_2),
    .COUT(\c$196 ),
    .SUM(\s$197 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_0_77_0 (.A(pp_row77_0),
    .B(pp_row77_1),
    .CIN(pp_row77_2),
    .COUT(\c$200 ),
    .SUM(\s$201 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_36_0 (.A(pp_row36_0),
    .B(pp_row36_1),
    .CIN(pp_row36_2),
    .COUT(\c$208 ),
    .SUM(\s$209 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_37_0 (.A(pp_row37_0),
    .B(pp_row37_1),
    .CIN(pp_row37_2),
    .COUT(\c$212 ),
    .SUM(\s$213 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_38_0 (.A(pp_row38_0),
    .B(pp_row38_1),
    .CIN(pp_row38_2),
    .COUT(\c$216 ),
    .SUM(\s$217 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_38_1 (.A(pp_row38_3),
    .B(pp_row38_4),
    .CIN(pp_row38_5),
    .COUT(\c$218 ),
    .SUM(\s$219 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_39_0 (.A(pp_row39_0),
    .B(pp_row39_1),
    .CIN(pp_row39_2),
    .COUT(\c$222 ),
    .SUM(\s$223 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_39_1 (.A(pp_row39_3),
    .B(pp_row39_4),
    .CIN(pp_row39_5),
    .COUT(\c$224 ),
    .SUM(\s$225 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_40_0 (.A(pp_row40_0),
    .B(pp_row40_1),
    .CIN(pp_row40_2),
    .COUT(\c$228 ),
    .SUM(\s$229 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_40_1 (.A(pp_row40_3),
    .B(pp_row40_4),
    .CIN(pp_row40_5),
    .COUT(\c$230 ),
    .SUM(\s$231 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_40_2 (.A(pp_row40_6),
    .B(pp_row40_7),
    .CIN(pp_row40_8),
    .COUT(\c$232 ),
    .SUM(\s$233 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_41_0 (.A(pp_row41_0),
    .B(pp_row41_1),
    .CIN(pp_row41_2),
    .COUT(\c$236 ),
    .SUM(\s$237 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_41_1 (.A(pp_row41_3),
    .B(pp_row41_4),
    .CIN(pp_row41_5),
    .COUT(\c$238 ),
    .SUM(\s$239 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_41_2 (.A(pp_row41_6),
    .B(pp_row41_7),
    .CIN(pp_row41_8),
    .COUT(\c$240 ),
    .SUM(\s$241 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_42_0 (.A(pp_row42_0),
    .B(pp_row42_1),
    .CIN(pp_row42_2),
    .COUT(\c$244 ),
    .SUM(\s$245 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_42_1 (.A(pp_row42_3),
    .B(pp_row42_4),
    .CIN(pp_row42_5),
    .COUT(\c$246 ),
    .SUM(\s$247 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_42_2 (.A(pp_row42_6),
    .B(pp_row42_7),
    .CIN(pp_row42_8),
    .COUT(\c$248 ),
    .SUM(\s$249 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_42_3 (.A(pp_row42_9),
    .B(pp_row42_10),
    .CIN(pp_row42_11),
    .COUT(\c$250 ),
    .SUM(\s$251 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_43_0 (.A(pp_row43_0),
    .B(pp_row43_1),
    .CIN(pp_row43_2),
    .COUT(\c$254 ),
    .SUM(\s$255 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_43_1 (.A(pp_row43_3),
    .B(pp_row43_4),
    .CIN(pp_row43_5),
    .COUT(\c$256 ),
    .SUM(\s$257 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_43_2 (.A(pp_row43_6),
    .B(pp_row43_7),
    .CIN(pp_row43_8),
    .COUT(\c$258 ),
    .SUM(\s$259 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_43_3 (.A(pp_row43_9),
    .B(pp_row43_10),
    .CIN(pp_row43_11),
    .COUT(\c$260 ),
    .SUM(\s$261 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_44_0 (.A(pp_row44_0),
    .B(pp_row44_1),
    .CIN(pp_row44_2),
    .COUT(\c$264 ),
    .SUM(\s$265 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_44_1 (.A(pp_row44_3),
    .B(pp_row44_4),
    .CIN(pp_row44_5),
    .COUT(\c$266 ),
    .SUM(\s$267 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_44_2 (.A(pp_row44_6),
    .B(pp_row44_7),
    .CIN(pp_row44_8),
    .COUT(\c$268 ),
    .SUM(\s$269 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_44_3 (.A(pp_row44_9),
    .B(pp_row44_10),
    .CIN(pp_row44_11),
    .COUT(\c$270 ),
    .SUM(\s$271 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_44_4 (.A(pp_row44_12),
    .B(pp_row44_13),
    .CIN(pp_row44_14),
    .COUT(\c$272 ),
    .SUM(\s$273 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_45_0 (.A(pp_row45_0),
    .B(pp_row45_1),
    .CIN(pp_row45_2),
    .COUT(\c$276 ),
    .SUM(\s$277 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_45_1 (.A(pp_row45_3),
    .B(pp_row45_4),
    .CIN(pp_row45_5),
    .COUT(\c$278 ),
    .SUM(\s$279 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_45_2 (.A(pp_row45_6),
    .B(pp_row45_7),
    .CIN(pp_row45_8),
    .COUT(\c$280 ),
    .SUM(\s$281 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_45_3 (.A(pp_row45_9),
    .B(pp_row45_10),
    .CIN(pp_row45_11),
    .COUT(\c$282 ),
    .SUM(\s$283 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_45_4 (.A(pp_row45_12),
    .B(pp_row45_13),
    .CIN(pp_row45_14),
    .COUT(\c$284 ),
    .SUM(\s$285 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_46_0 (.A(pp_row46_0),
    .B(pp_row46_1),
    .CIN(pp_row46_2),
    .COUT(\c$288 ),
    .SUM(\s$289 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_46_1 (.A(pp_row46_3),
    .B(pp_row46_4),
    .CIN(pp_row46_5),
    .COUT(\c$290 ),
    .SUM(\s$291 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_46_2 (.A(pp_row46_6),
    .B(pp_row46_7),
    .CIN(pp_row46_8),
    .COUT(\c$292 ),
    .SUM(\s$293 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_46_3 (.A(pp_row46_9),
    .B(pp_row46_10),
    .CIN(pp_row46_11),
    .COUT(\c$294 ),
    .SUM(\s$295 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_46_4 (.A(pp_row46_12),
    .B(pp_row46_13),
    .CIN(pp_row46_14),
    .COUT(\c$296 ),
    .SUM(\s$297 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_46_5 (.A(pp_row46_15),
    .B(pp_row46_16),
    .CIN(pp_row46_17),
    .COUT(\c$298 ),
    .SUM(\s$299 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_47_0 (.A(pp_row47_0),
    .B(pp_row47_1),
    .CIN(pp_row47_2),
    .COUT(\c$302 ),
    .SUM(\s$303 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_47_1 (.A(pp_row47_3),
    .B(pp_row47_4),
    .CIN(pp_row47_5),
    .COUT(\c$304 ),
    .SUM(\s$305 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_47_2 (.A(pp_row47_6),
    .B(pp_row47_7),
    .CIN(pp_row47_8),
    .COUT(\c$306 ),
    .SUM(\s$307 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_47_3 (.A(pp_row47_9),
    .B(pp_row47_10),
    .CIN(pp_row47_11),
    .COUT(\c$308 ),
    .SUM(\s$309 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_47_4 (.A(pp_row47_12),
    .B(pp_row47_13),
    .CIN(pp_row47_14),
    .COUT(\c$310 ),
    .SUM(\s$311 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_47_5 (.A(pp_row47_15),
    .B(pp_row47_16),
    .CIN(pp_row47_17),
    .COUT(\c$312 ),
    .SUM(\s$313 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_48_0 (.A(pp_row48_0),
    .B(pp_row48_1),
    .CIN(pp_row48_2),
    .COUT(\c$316 ),
    .SUM(\s$317 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_48_1 (.A(pp_row48_3),
    .B(pp_row48_4),
    .CIN(pp_row48_5),
    .COUT(\c$318 ),
    .SUM(\s$319 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_48_2 (.A(pp_row48_6),
    .B(pp_row48_7),
    .CIN(pp_row48_8),
    .COUT(\c$320 ),
    .SUM(\s$321 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_48_3 (.A(pp_row48_9),
    .B(pp_row48_10),
    .CIN(pp_row48_11),
    .COUT(\c$322 ),
    .SUM(\s$323 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_48_4 (.A(pp_row48_12),
    .B(pp_row48_13),
    .CIN(pp_row48_14),
    .COUT(\c$324 ),
    .SUM(\s$325 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_48_5 (.A(pp_row48_15),
    .B(pp_row48_16),
    .CIN(pp_row48_17),
    .COUT(\c$326 ),
    .SUM(\s$327 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_48_6 (.A(pp_row48_18),
    .B(pp_row48_19),
    .CIN(pp_row48_20),
    .COUT(\c$328 ),
    .SUM(\s$329 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_49_0 (.A(pp_row49_0),
    .B(pp_row49_1),
    .CIN(pp_row49_2),
    .COUT(\c$332 ),
    .SUM(\s$333 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_49_1 (.A(pp_row49_3),
    .B(pp_row49_4),
    .CIN(pp_row49_5),
    .COUT(\c$334 ),
    .SUM(\s$335 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_49_2 (.A(pp_row49_6),
    .B(pp_row49_7),
    .CIN(pp_row49_8),
    .COUT(\c$336 ),
    .SUM(\s$337 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_49_3 (.A(pp_row49_9),
    .B(pp_row49_10),
    .CIN(pp_row49_11),
    .COUT(\c$338 ),
    .SUM(\s$339 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_49_4 (.A(pp_row49_12),
    .B(pp_row49_13),
    .CIN(pp_row49_14),
    .COUT(\c$340 ),
    .SUM(\s$341 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_49_5 (.A(pp_row49_15),
    .B(pp_row49_16),
    .CIN(pp_row49_17),
    .COUT(\c$342 ),
    .SUM(\s$343 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_49_6 (.A(pp_row49_18),
    .B(pp_row49_19),
    .CIN(pp_row49_20),
    .COUT(\c$344 ),
    .SUM(\s$345 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_50_0 (.A(pp_row50_0),
    .B(pp_row50_1),
    .CIN(pp_row50_2),
    .COUT(\c$348 ),
    .SUM(\s$349 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_50_1 (.A(pp_row50_3),
    .B(pp_row50_4),
    .CIN(pp_row50_5),
    .COUT(\c$350 ),
    .SUM(\s$351 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_50_2 (.A(pp_row50_6),
    .B(pp_row50_7),
    .CIN(pp_row50_8),
    .COUT(\c$352 ),
    .SUM(\s$353 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_50_3 (.A(pp_row50_9),
    .B(pp_row50_10),
    .CIN(pp_row50_11),
    .COUT(\c$354 ),
    .SUM(\s$355 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_50_4 (.A(pp_row50_12),
    .B(pp_row50_13),
    .CIN(pp_row50_14),
    .COUT(\c$356 ),
    .SUM(\s$357 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_50_5 (.A(pp_row50_15),
    .B(pp_row50_16),
    .CIN(pp_row50_17),
    .COUT(\c$358 ),
    .SUM(\s$359 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_50_6 (.A(pp_row50_18),
    .B(pp_row50_19),
    .CIN(pp_row50_20),
    .COUT(\c$360 ),
    .SUM(\s$361 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_50_7 (.A(pp_row50_21),
    .B(pp_row50_22),
    .CIN(pp_row50_23),
    .COUT(\c$362 ),
    .SUM(\s$363 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_51_0 (.A(pp_row51_0),
    .B(pp_row51_1),
    .CIN(pp_row51_2),
    .COUT(\c$366 ),
    .SUM(\s$367 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_51_1 (.A(pp_row51_3),
    .B(pp_row51_4),
    .CIN(pp_row51_5),
    .COUT(\c$368 ),
    .SUM(\s$369 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_51_2 (.A(pp_row51_6),
    .B(pp_row51_7),
    .CIN(pp_row51_8),
    .COUT(\c$370 ),
    .SUM(\s$371 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_51_3 (.A(pp_row51_9),
    .B(pp_row51_10),
    .CIN(pp_row51_11),
    .COUT(\c$372 ),
    .SUM(\s$373 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_51_4 (.A(pp_row51_12),
    .B(pp_row51_13),
    .CIN(pp_row51_14),
    .COUT(\c$374 ),
    .SUM(\s$375 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_51_5 (.A(pp_row51_15),
    .B(pp_row51_16),
    .CIN(pp_row51_17),
    .COUT(\c$376 ),
    .SUM(\s$377 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_51_6 (.A(pp_row51_18),
    .B(pp_row51_19),
    .CIN(pp_row51_20),
    .COUT(\c$378 ),
    .SUM(\s$379 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_51_7 (.A(pp_row51_21),
    .B(pp_row51_22),
    .CIN(pp_row51_23),
    .COUT(\c$380 ),
    .SUM(\s$381 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_52_0 (.A(pp_row52_2),
    .B(pp_row52_3),
    .CIN(pp_row52_4),
    .COUT(\c$384 ),
    .SUM(\s$385 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_52_1 (.A(pp_row52_5),
    .B(pp_row52_6),
    .CIN(pp_row52_7),
    .COUT(\c$386 ),
    .SUM(\s$387 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_52_2 (.A(pp_row52_8),
    .B(pp_row52_9),
    .CIN(pp_row52_10),
    .COUT(\c$388 ),
    .SUM(\s$389 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_52_3 (.A(pp_row52_11),
    .B(pp_row52_12),
    .CIN(pp_row52_13),
    .COUT(\c$390 ),
    .SUM(\s$391 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_52_4 (.A(pp_row52_14),
    .B(pp_row52_15),
    .CIN(pp_row52_16),
    .COUT(\c$392 ),
    .SUM(\s$393 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_52_5 (.A(pp_row52_17),
    .B(pp_row52_18),
    .CIN(pp_row52_19),
    .COUT(\c$394 ),
    .SUM(\s$395 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_52_6 (.A(pp_row52_20),
    .B(pp_row52_21),
    .CIN(pp_row52_22),
    .COUT(\c$396 ),
    .SUM(\s$397 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_52_7 (.A(pp_row52_23),
    .B(pp_row52_24),
    .CIN(pp_row52_25),
    .COUT(\c$398 ),
    .SUM(\s$399 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_52_8 (.A(pp_row52_26),
    .B(pp_row52_27),
    .CIN(pp_row52_28),
    .COUT(\c$400 ),
    .SUM(\s$401 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_53_0 (.A(pp_row53_2),
    .B(pp_row53_3),
    .CIN(pp_row53_4),
    .COUT(\c$402 ),
    .SUM(\s$403 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_53_1 (.A(pp_row53_5),
    .B(pp_row53_6),
    .CIN(pp_row53_7),
    .COUT(\c$404 ),
    .SUM(\s$405 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_53_2 (.A(pp_row53_8),
    .B(pp_row53_9),
    .CIN(pp_row53_10),
    .COUT(\c$406 ),
    .SUM(\s$407 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_53_3 (.A(pp_row53_11),
    .B(pp_row53_12),
    .CIN(pp_row53_13),
    .COUT(\c$408 ),
    .SUM(\s$409 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_53_4 (.A(pp_row53_14),
    .B(pp_row53_15),
    .CIN(pp_row53_16),
    .COUT(\c$410 ),
    .SUM(\s$411 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_53_5 (.A(pp_row53_17),
    .B(pp_row53_18),
    .CIN(pp_row53_19),
    .COUT(\c$412 ),
    .SUM(\s$413 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_53_6 (.A(pp_row53_20),
    .B(pp_row53_21),
    .CIN(pp_row53_22),
    .COUT(\c$414 ),
    .SUM(\s$415 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_53_7 (.A(pp_row53_23),
    .B(pp_row53_24),
    .CIN(pp_row53_25),
    .COUT(\c$416 ),
    .SUM(\s$417 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_53_8 (.A(pp_row53_26),
    .B(pp_row53_27),
    .CIN(\c$1 ),
    .COUT(\c$418 ),
    .SUM(\s$419 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_54_0 (.A(pp_row54_5),
    .B(pp_row54_6),
    .CIN(pp_row54_7),
    .COUT(\c$420 ),
    .SUM(\s$421 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_54_1 (.A(pp_row54_8),
    .B(pp_row54_9),
    .CIN(pp_row54_10),
    .COUT(\c$422 ),
    .SUM(\s$423 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_54_2 (.A(pp_row54_11),
    .B(pp_row54_12),
    .CIN(pp_row54_13),
    .COUT(\c$424 ),
    .SUM(\s$425 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_54_3 (.A(pp_row54_14),
    .B(pp_row54_15),
    .CIN(pp_row54_16),
    .COUT(\c$426 ),
    .SUM(\s$427 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_54_4 (.A(pp_row54_17),
    .B(pp_row54_18),
    .CIN(pp_row54_19),
    .COUT(\c$428 ),
    .SUM(\s$429 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_54_5 (.A(pp_row54_20),
    .B(pp_row54_21),
    .CIN(pp_row54_22),
    .COUT(\c$430 ),
    .SUM(\s$431 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_54_6 (.A(pp_row54_23),
    .B(pp_row54_24),
    .CIN(pp_row54_25),
    .COUT(\c$432 ),
    .SUM(\s$433 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_54_7 (.A(pp_row54_26),
    .B(pp_row54_27),
    .CIN(pp_row54_28),
    .COUT(\c$434 ),
    .SUM(\s$435 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_54_8 (.A(pp_row54_29),
    .B(\c$2 ),
    .CIN(\s$5 ),
    .COUT(\c$436 ),
    .SUM(\s$437 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_55_0 (.A(pp_row55_5),
    .B(pp_row55_6),
    .CIN(pp_row55_7),
    .COUT(\c$438 ),
    .SUM(\s$439 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_55_1 (.A(pp_row55_8),
    .B(pp_row55_9),
    .CIN(pp_row55_10),
    .COUT(\c$440 ),
    .SUM(\s$441 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_55_2 (.A(pp_row55_11),
    .B(pp_row55_12),
    .CIN(pp_row55_13),
    .COUT(\c$442 ),
    .SUM(\s$443 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_55_3 (.A(pp_row55_14),
    .B(pp_row55_15),
    .CIN(pp_row55_16),
    .COUT(\c$444 ),
    .SUM(\s$445 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_55_4 (.A(pp_row55_17),
    .B(pp_row55_18),
    .CIN(pp_row55_19),
    .COUT(\c$446 ),
    .SUM(\s$447 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_55_5 (.A(pp_row55_20),
    .B(pp_row55_21),
    .CIN(pp_row55_22),
    .COUT(\c$448 ),
    .SUM(\s$449 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_55_6 (.A(pp_row55_23),
    .B(pp_row55_24),
    .CIN(pp_row55_25),
    .COUT(\c$450 ),
    .SUM(\s$451 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_55_7 (.A(pp_row55_26),
    .B(pp_row55_27),
    .CIN(pp_row55_28),
    .COUT(\c$452 ),
    .SUM(\s$453 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_55_8 (.A(\c$4 ),
    .B(\c$6 ),
    .CIN(\s$9 ),
    .COUT(\c$454 ),
    .SUM(\s$455 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_56_0 (.A(pp_row56_8),
    .B(pp_row56_9),
    .CIN(pp_row56_10),
    .COUT(\c$456 ),
    .SUM(\s$457 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_56_1 (.A(pp_row56_11),
    .B(pp_row56_12),
    .CIN(pp_row56_13),
    .COUT(\c$458 ),
    .SUM(\s$459 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_56_2 (.A(pp_row56_14),
    .B(pp_row56_15),
    .CIN(pp_row56_16),
    .COUT(\c$460 ),
    .SUM(\s$461 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_56_3 (.A(pp_row56_17),
    .B(pp_row56_18),
    .CIN(pp_row56_19),
    .COUT(\c$462 ),
    .SUM(\s$463 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_56_4 (.A(pp_row56_20),
    .B(pp_row56_21),
    .CIN(pp_row56_22),
    .COUT(\c$464 ),
    .SUM(\s$465 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_56_5 (.A(pp_row56_23),
    .B(pp_row56_24),
    .CIN(pp_row56_25),
    .COUT(\c$466 ),
    .SUM(\s$467 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_56_6 (.A(pp_row56_26),
    .B(pp_row56_27),
    .CIN(pp_row56_28),
    .COUT(\c$468 ),
    .SUM(\s$469 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_56_7 (.A(pp_row56_29),
    .B(pp_row56_30),
    .CIN(\c$8 ),
    .COUT(\c$470 ),
    .SUM(\s$471 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_56_8 (.A(\c$10 ),
    .B(\s$13 ),
    .CIN(\s$15 ),
    .COUT(\c$472 ),
    .SUM(\s$473 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_57_0 (.A(pp_row57_8),
    .B(pp_row57_9),
    .CIN(pp_row57_10),
    .COUT(\c$474 ),
    .SUM(\s$475 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_57_1 (.A(pp_row57_11),
    .B(pp_row57_12),
    .CIN(pp_row57_13),
    .COUT(\c$476 ),
    .SUM(\s$477 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_57_2 (.A(pp_row57_14),
    .B(pp_row57_15),
    .CIN(pp_row57_16),
    .COUT(\c$478 ),
    .SUM(\s$479 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_57_3 (.A(pp_row57_17),
    .B(pp_row57_18),
    .CIN(pp_row57_19),
    .COUT(\c$480 ),
    .SUM(\s$481 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_57_4 (.A(pp_row57_20),
    .B(pp_row57_21),
    .CIN(pp_row57_22),
    .COUT(\c$482 ),
    .SUM(\s$483 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_57_5 (.A(pp_row57_23),
    .B(pp_row57_24),
    .CIN(pp_row57_25),
    .COUT(\c$484 ),
    .SUM(\s$485 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_57_6 (.A(pp_row57_26),
    .B(pp_row57_27),
    .CIN(pp_row57_28),
    .COUT(\c$486 ),
    .SUM(\s$487 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_57_7 (.A(pp_row57_29),
    .B(\c$12 ),
    .CIN(\c$14 ),
    .COUT(\c$488 ),
    .SUM(\s$489 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_57_8 (.A(\c$16 ),
    .B(\s$19 ),
    .CIN(\s$21 ),
    .COUT(\c$490 ),
    .SUM(\s$491 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_58_0 (.A(pp_row58_11),
    .B(pp_row58_12),
    .CIN(pp_row58_13),
    .COUT(\c$492 ),
    .SUM(\s$493 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_58_1 (.A(pp_row58_14),
    .B(pp_row58_15),
    .CIN(pp_row58_16),
    .COUT(\c$494 ),
    .SUM(\s$495 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_58_2 (.A(pp_row58_17),
    .B(pp_row58_18),
    .CIN(pp_row58_19),
    .COUT(\c$496 ),
    .SUM(\s$497 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_58_3 (.A(pp_row58_20),
    .B(pp_row58_21),
    .CIN(pp_row58_22),
    .COUT(\c$498 ),
    .SUM(\s$499 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_58_4 (.A(pp_row58_23),
    .B(pp_row58_24),
    .CIN(pp_row58_25),
    .COUT(\c$500 ),
    .SUM(\s$501 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_58_5 (.A(pp_row58_26),
    .B(pp_row58_27),
    .CIN(pp_row58_28),
    .COUT(\c$502 ),
    .SUM(\s$503 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_58_6 (.A(pp_row58_29),
    .B(pp_row58_30),
    .CIN(pp_row58_31),
    .COUT(\c$504 ),
    .SUM(\s$505 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_58_7 (.A(\c$18 ),
    .B(\c$20 ),
    .CIN(\c$22 ),
    .COUT(\c$506 ),
    .SUM(\s$507 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_58_8 (.A(\s$25 ),
    .B(\s$27 ),
    .CIN(\s$29 ),
    .COUT(\c$508 ),
    .SUM(\s$509 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_59_0 (.A(pp_row59_11),
    .B(pp_row59_12),
    .CIN(pp_row59_13),
    .COUT(\c$510 ),
    .SUM(\s$511 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_59_1 (.A(pp_row59_14),
    .B(pp_row59_15),
    .CIN(pp_row59_16),
    .COUT(\c$512 ),
    .SUM(\s$513 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_59_2 (.A(pp_row59_17),
    .B(pp_row59_18),
    .CIN(pp_row59_19),
    .COUT(\c$514 ),
    .SUM(\s$515 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_59_3 (.A(pp_row59_20),
    .B(pp_row59_21),
    .CIN(pp_row59_22),
    .COUT(\c$516 ),
    .SUM(\s$517 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_59_4 (.A(pp_row59_23),
    .B(pp_row59_24),
    .CIN(pp_row59_25),
    .COUT(\c$518 ),
    .SUM(\s$519 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_59_5 (.A(pp_row59_26),
    .B(pp_row59_27),
    .CIN(pp_row59_28),
    .COUT(\c$520 ),
    .SUM(\s$521 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_59_6 (.A(pp_row59_29),
    .B(pp_row59_30),
    .CIN(\c$24 ),
    .COUT(\c$522 ),
    .SUM(\s$523 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_59_7 (.A(\c$26 ),
    .B(\c$28 ),
    .CIN(\c$30 ),
    .COUT(\c$524 ),
    .SUM(\s$525 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_59_8 (.A(\s$33 ),
    .B(\s$35 ),
    .CIN(\s$37 ),
    .COUT(\c$526 ),
    .SUM(\s$527 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_60_0 (.A(pp_row60_14),
    .B(pp_row60_15),
    .CIN(pp_row60_16),
    .COUT(\c$528 ),
    .SUM(\s$529 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_60_1 (.A(pp_row60_17),
    .B(pp_row60_18),
    .CIN(pp_row60_19),
    .COUT(\c$530 ),
    .SUM(\s$531 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_60_2 (.A(pp_row60_20),
    .B(pp_row60_21),
    .CIN(pp_row60_22),
    .COUT(\c$532 ),
    .SUM(\s$533 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_60_3 (.A(pp_row60_23),
    .B(pp_row60_24),
    .CIN(pp_row60_25),
    .COUT(\c$534 ),
    .SUM(\s$535 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_60_4 (.A(pp_row60_26),
    .B(pp_row60_27),
    .CIN(pp_row60_28),
    .COUT(\c$536 ),
    .SUM(\s$537 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_60_5 (.A(pp_row60_29),
    .B(pp_row60_30),
    .CIN(pp_row60_31),
    .COUT(\c$538 ),
    .SUM(\s$539 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_60_6 (.A(pp_row60_32),
    .B(\c$32 ),
    .CIN(\c$34 ),
    .COUT(\c$540 ),
    .SUM(\s$541 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_60_7 (.A(\c$36 ),
    .B(\c$38 ),
    .CIN(\s$41 ),
    .COUT(\c$542 ),
    .SUM(\s$543 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_60_8 (.A(\s$43 ),
    .B(\s$45 ),
    .CIN(\s$47 ),
    .COUT(\c$544 ),
    .SUM(\s$545 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_61_0 (.A(pp_row61_14),
    .B(pp_row61_15),
    .CIN(pp_row61_16),
    .COUT(\c$546 ),
    .SUM(\s$547 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_61_1 (.A(pp_row61_17),
    .B(pp_row61_18),
    .CIN(pp_row61_19),
    .COUT(\c$548 ),
    .SUM(\s$549 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_61_2 (.A(pp_row61_20),
    .B(pp_row61_21),
    .CIN(pp_row61_22),
    .COUT(\c$550 ),
    .SUM(\s$551 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_61_3 (.A(pp_row61_23),
    .B(pp_row61_24),
    .CIN(pp_row61_25),
    .COUT(\c$552 ),
    .SUM(\s$553 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_61_4 (.A(pp_row61_26),
    .B(pp_row61_27),
    .CIN(pp_row61_28),
    .COUT(\c$554 ),
    .SUM(\s$555 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_61_5 (.A(pp_row61_29),
    .B(pp_row61_30),
    .CIN(pp_row61_31),
    .COUT(\c$556 ),
    .SUM(\s$557 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_61_6 (.A(\c$40 ),
    .B(\c$42 ),
    .CIN(\c$44 ),
    .COUT(\c$558 ),
    .SUM(\s$559 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_61_7 (.A(\c$46 ),
    .B(\c$48 ),
    .CIN(\s$51 ),
    .COUT(\c$560 ),
    .SUM(\s$561 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_61_8 (.A(\s$53 ),
    .B(\s$55 ),
    .CIN(\s$57 ),
    .COUT(\c$562 ),
    .SUM(\s$563 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_62_0 (.A(pp_row62_17),
    .B(pp_row62_18),
    .CIN(pp_row62_19),
    .COUT(\c$564 ),
    .SUM(\s$565 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_62_1 (.A(pp_row62_20),
    .B(pp_row62_21),
    .CIN(pp_row62_22),
    .COUT(\c$566 ),
    .SUM(\s$567 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_62_2 (.A(pp_row62_23),
    .B(pp_row62_24),
    .CIN(pp_row62_25),
    .COUT(\c$568 ),
    .SUM(\s$569 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_62_3 (.A(pp_row62_26),
    .B(pp_row62_27),
    .CIN(pp_row62_28),
    .COUT(\c$570 ),
    .SUM(\s$571 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_62_4 (.A(pp_row62_29),
    .B(pp_row62_30),
    .CIN(pp_row62_31),
    .COUT(\c$572 ),
    .SUM(\s$573 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_62_5 (.A(pp_row62_32),
    .B(pp_row62_33),
    .CIN(\c$50 ),
    .COUT(\c$574 ),
    .SUM(\s$575 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_62_6 (.A(\c$52 ),
    .B(\c$54 ),
    .CIN(\c$56 ),
    .COUT(\c$576 ),
    .SUM(\s$577 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_62_7 (.A(\c$58 ),
    .B(\s$61 ),
    .CIN(\s$63 ),
    .COUT(\c$578 ),
    .SUM(\s$579 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_62_8 (.A(\s$65 ),
    .B(\s$67 ),
    .CIN(\s$69 ),
    .COUT(\c$580 ),
    .SUM(\s$581 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_63_0 (.A(pp_row63_17),
    .B(pp_row63_18),
    .CIN(pp_row63_19),
    .COUT(\c$582 ),
    .SUM(\s$583 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_63_1 (.A(pp_row63_20),
    .B(pp_row63_21),
    .CIN(pp_row63_22),
    .COUT(\c$584 ),
    .SUM(\s$585 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_63_2 (.A(pp_row63_23),
    .B(pp_row63_24),
    .CIN(pp_row63_25),
    .COUT(\c$586 ),
    .SUM(\s$587 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_63_3 (.A(pp_row63_26),
    .B(pp_row63_27),
    .CIN(pp_row63_28),
    .COUT(\c$588 ),
    .SUM(\s$589 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_63_4 (.A(pp_row63_29),
    .B(pp_row63_30),
    .CIN(pp_row63_31),
    .COUT(\c$590 ),
    .SUM(\s$591 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_63_5 (.A(pp_row63_32),
    .B(\c$60 ),
    .CIN(\c$62 ),
    .COUT(\c$592 ),
    .SUM(\s$593 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_63_6 (.A(\c$64 ),
    .B(\c$66 ),
    .CIN(\c$68 ),
    .COUT(\c$594 ),
    .SUM(\s$595 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_63_7 (.A(\c$70 ),
    .B(\s$73 ),
    .CIN(\s$75 ),
    .COUT(\c$596 ),
    .SUM(\s$597 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_63_8 (.A(\s$77 ),
    .B(\s$79 ),
    .CIN(\s$81 ),
    .COUT(\c$598 ),
    .SUM(\s$599 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_64_0 (.A(pp_row64_18),
    .B(pp_row64_19),
    .CIN(pp_row64_20),
    .COUT(\c$600 ),
    .SUM(\s$601 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_64_1 (.A(pp_row64_21),
    .B(pp_row64_22),
    .CIN(pp_row64_23),
    .COUT(\c$602 ),
    .SUM(\s$603 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_64_2 (.A(pp_row64_24),
    .B(pp_row64_25),
    .CIN(pp_row64_26),
    .COUT(\c$604 ),
    .SUM(\s$605 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_64_3 (.A(pp_row64_27),
    .B(pp_row64_28),
    .CIN(pp_row64_29),
    .COUT(\c$606 ),
    .SUM(\s$607 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_64_4 (.A(pp_row64_30),
    .B(pp_row64_31),
    .CIN(pp_row64_32),
    .COUT(\c$608 ),
    .SUM(\s$609 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_64_5 (.A(pp_row64_33),
    .B(\c$72 ),
    .CIN(\c$74 ),
    .COUT(\c$610 ),
    .SUM(\s$611 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_64_6 (.A(\c$76 ),
    .B(\c$78 ),
    .CIN(\c$80 ),
    .COUT(\c$612 ),
    .SUM(\s$613 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_64_7 (.A(\c$82 ),
    .B(\s$85 ),
    .CIN(\s$87 ),
    .COUT(\c$614 ),
    .SUM(\s$615 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_64_8 (.A(\s$89 ),
    .B(\s$91 ),
    .CIN(\s$93 ),
    .COUT(\c$616 ),
    .SUM(\s$617 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_65_0 (.A(pp_row65_18),
    .B(pp_row65_19),
    .CIN(pp_row65_20),
    .COUT(\c$618 ),
    .SUM(\s$619 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_65_1 (.A(pp_row65_21),
    .B(pp_row65_22),
    .CIN(pp_row65_23),
    .COUT(\c$620 ),
    .SUM(\s$621 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_65_2 (.A(pp_row65_24),
    .B(pp_row65_25),
    .CIN(pp_row65_26),
    .COUT(\c$622 ),
    .SUM(\s$623 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_65_3 (.A(pp_row65_27),
    .B(pp_row65_28),
    .CIN(pp_row65_29),
    .COUT(\c$624 ),
    .SUM(\s$625 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_65_4 (.A(pp_row65_30),
    .B(pp_row65_31),
    .CIN(pp_row65_32),
    .COUT(\c$626 ),
    .SUM(\s$627 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_65_5 (.A(pp_row65_33),
    .B(\c$84 ),
    .CIN(\c$86 ),
    .COUT(\c$628 ),
    .SUM(\s$629 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_65_6 (.A(\c$88 ),
    .B(\c$90 ),
    .CIN(\c$92 ),
    .COUT(\c$630 ),
    .SUM(\s$631 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_65_7 (.A(\c$94 ),
    .B(\s$97 ),
    .CIN(\s$99 ),
    .COUT(\c$632 ),
    .SUM(\s$633 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_65_8 (.A(\s$101 ),
    .B(\s$103 ),
    .CIN(\s$105 ),
    .COUT(\c$634 ),
    .SUM(\s$635 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_66_0 (.A(pp_row66_18),
    .B(pp_row66_19),
    .CIN(pp_row66_20),
    .COUT(\c$636 ),
    .SUM(\s$637 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_66_1 (.A(pp_row66_21),
    .B(pp_row66_22),
    .CIN(pp_row66_23),
    .COUT(\c$638 ),
    .SUM(\s$639 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_66_2 (.A(pp_row66_24),
    .B(pp_row66_25),
    .CIN(pp_row66_26),
    .COUT(\c$640 ),
    .SUM(\s$641 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_66_3 (.A(pp_row66_27),
    .B(pp_row66_28),
    .CIN(pp_row66_29),
    .COUT(\c$642 ),
    .SUM(\s$643 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_66_4 (.A(pp_row66_30),
    .B(pp_row66_31),
    .CIN(pp_row66_32),
    .COUT(\c$644 ),
    .SUM(\s$645 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_66_5 (.A(pp_row66_33),
    .B(\c$96 ),
    .CIN(\c$98 ),
    .COUT(\c$646 ),
    .SUM(\s$647 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_66_6 (.A(\c$100 ),
    .B(\c$102 ),
    .CIN(\c$104 ),
    .COUT(\c$648 ),
    .SUM(\s$649 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_66_7 (.A(\c$106 ),
    .B(\s$109 ),
    .CIN(\s$111 ),
    .COUT(\c$650 ),
    .SUM(\s$651 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_66_8 (.A(\s$113 ),
    .B(\s$115 ),
    .CIN(\s$117 ),
    .COUT(\c$652 ),
    .SUM(\s$653 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_67_0 (.A(pp_row67_18),
    .B(pp_row67_19),
    .CIN(pp_row67_20),
    .COUT(\c$654 ),
    .SUM(\s$655 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_67_1 (.A(pp_row67_21),
    .B(pp_row67_22),
    .CIN(pp_row67_23),
    .COUT(\c$656 ),
    .SUM(\s$657 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_67_2 (.A(pp_row67_24),
    .B(pp_row67_25),
    .CIN(pp_row67_26),
    .COUT(\c$658 ),
    .SUM(\s$659 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_67_3 (.A(pp_row67_27),
    .B(pp_row67_28),
    .CIN(pp_row67_29),
    .COUT(\c$660 ),
    .SUM(\s$661 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_67_4 (.A(pp_row67_30),
    .B(pp_row67_31),
    .CIN(pp_row67_32),
    .COUT(\c$662 ),
    .SUM(\s$663 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_67_5 (.A(pp_row67_33),
    .B(\c$108 ),
    .CIN(\c$110 ),
    .COUT(\c$664 ),
    .SUM(\s$665 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_67_6 (.A(\c$112 ),
    .B(\c$114 ),
    .CIN(\c$116 ),
    .COUT(\c$666 ),
    .SUM(\s$667 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_67_7 (.A(\c$118 ),
    .B(\s$121 ),
    .CIN(\s$123 ),
    .COUT(\c$668 ),
    .SUM(\s$669 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_67_8 (.A(\s$125 ),
    .B(\s$127 ),
    .CIN(\s$129 ),
    .COUT(\c$670 ),
    .SUM(\s$671 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_68_0 (.A(pp_row68_17),
    .B(pp_row68_18),
    .CIN(pp_row68_19),
    .COUT(\c$672 ),
    .SUM(\s$673 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_68_1 (.A(pp_row68_20),
    .B(pp_row68_21),
    .CIN(pp_row68_22),
    .COUT(\c$674 ),
    .SUM(\s$675 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_68_2 (.A(pp_row68_23),
    .B(pp_row68_24),
    .CIN(pp_row68_25),
    .COUT(\c$676 ),
    .SUM(\s$677 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_68_3 (.A(pp_row68_26),
    .B(pp_row68_27),
    .CIN(pp_row68_28),
    .COUT(\c$678 ),
    .SUM(\s$679 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_68_4 (.A(pp_row68_29),
    .B(pp_row68_30),
    .CIN(pp_row68_31),
    .COUT(\c$680 ),
    .SUM(\s$681 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_68_5 (.A(pp_row68_32),
    .B(\c$120 ),
    .CIN(\c$122 ),
    .COUT(\c$682 ),
    .SUM(\s$683 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_68_6 (.A(\c$124 ),
    .B(\c$126 ),
    .CIN(\c$128 ),
    .COUT(\c$684 ),
    .SUM(\s$685 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_68_7 (.A(\c$130 ),
    .B(\s$133 ),
    .CIN(\s$135 ),
    .COUT(\c$686 ),
    .SUM(\s$687 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_68_8 (.A(\s$137 ),
    .B(\s$139 ),
    .CIN(\s$141 ),
    .COUT(\c$688 ),
    .SUM(\s$689 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_69_0 (.A(pp_row69_15),
    .B(pp_row69_16),
    .CIN(pp_row69_17),
    .COUT(\c$690 ),
    .SUM(\s$691 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_69_1 (.A(pp_row69_18),
    .B(pp_row69_19),
    .CIN(pp_row69_20),
    .COUT(\c$692 ),
    .SUM(\s$693 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_69_2 (.A(pp_row69_21),
    .B(pp_row69_22),
    .CIN(pp_row69_23),
    .COUT(\c$694 ),
    .SUM(\s$695 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_69_3 (.A(pp_row69_24),
    .B(pp_row69_25),
    .CIN(pp_row69_26),
    .COUT(\c$696 ),
    .SUM(\s$697 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_69_4 (.A(pp_row69_27),
    .B(pp_row69_28),
    .CIN(pp_row69_29),
    .COUT(\c$698 ),
    .SUM(\s$699 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_69_5 (.A(pp_row69_30),
    .B(pp_row69_31),
    .CIN(\c$132 ),
    .COUT(\c$700 ),
    .SUM(\s$701 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_69_6 (.A(\c$134 ),
    .B(\c$136 ),
    .CIN(\c$138 ),
    .COUT(\c$702 ),
    .SUM(\s$703 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_69_7 (.A(\c$140 ),
    .B(\c$142 ),
    .CIN(\s$145 ),
    .COUT(\c$704 ),
    .SUM(\s$705 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_69_8 (.A(\s$147 ),
    .B(\s$149 ),
    .CIN(\s$151 ),
    .COUT(\c$706 ),
    .SUM(\s$707 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_70_0 (.A(pp_row70_14),
    .B(pp_row70_15),
    .CIN(pp_row70_16),
    .COUT(\c$708 ),
    .SUM(\s$709 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_70_1 (.A(pp_row70_17),
    .B(pp_row70_18),
    .CIN(pp_row70_19),
    .COUT(\c$710 ),
    .SUM(\s$711 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_70_2 (.A(pp_row70_20),
    .B(pp_row70_21),
    .CIN(pp_row70_22),
    .COUT(\c$712 ),
    .SUM(\s$713 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_70_3 (.A(pp_row70_23),
    .B(pp_row70_24),
    .CIN(pp_row70_25),
    .COUT(\c$714 ),
    .SUM(\s$715 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_70_4 (.A(pp_row70_26),
    .B(pp_row70_27),
    .CIN(pp_row70_28),
    .COUT(\c$716 ),
    .SUM(\s$717 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_70_5 (.A(pp_row70_29),
    .B(pp_row70_30),
    .CIN(pp_row70_31),
    .COUT(\c$718 ),
    .SUM(\s$719 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_70_6 (.A(\c$144 ),
    .B(\c$146 ),
    .CIN(\c$148 ),
    .COUT(\c$720 ),
    .SUM(\s$721 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_70_7 (.A(\c$150 ),
    .B(\c$152 ),
    .CIN(\s$155 ),
    .COUT(\c$722 ),
    .SUM(\s$723 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_70_8 (.A(\s$157 ),
    .B(\s$159 ),
    .CIN(\s$161 ),
    .COUT(\c$724 ),
    .SUM(\s$725 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_71_0 (.A(pp_row71_12),
    .B(pp_row71_13),
    .CIN(pp_row71_14),
    .COUT(\c$726 ),
    .SUM(\s$727 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_71_1 (.A(pp_row71_15),
    .B(pp_row71_16),
    .CIN(pp_row71_17),
    .COUT(\c$728 ),
    .SUM(\s$729 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_71_2 (.A(pp_row71_18),
    .B(pp_row71_19),
    .CIN(pp_row71_20),
    .COUT(\c$730 ),
    .SUM(\s$731 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_71_3 (.A(pp_row71_21),
    .B(pp_row71_22),
    .CIN(pp_row71_23),
    .COUT(\c$732 ),
    .SUM(\s$733 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_71_4 (.A(pp_row71_24),
    .B(pp_row71_25),
    .CIN(pp_row71_26),
    .COUT(\c$734 ),
    .SUM(\s$735 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_71_5 (.A(pp_row71_27),
    .B(pp_row71_28),
    .CIN(pp_row71_29),
    .COUT(\c$736 ),
    .SUM(\s$737 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_71_6 (.A(pp_row71_30),
    .B(\c$154 ),
    .CIN(\c$156 ),
    .COUT(\c$738 ),
    .SUM(\s$739 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_71_7 (.A(\c$158 ),
    .B(\c$160 ),
    .CIN(\c$162 ),
    .COUT(\c$740 ),
    .SUM(\s$741 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_71_8 (.A(\s$165 ),
    .B(\s$167 ),
    .CIN(\s$169 ),
    .COUT(\c$742 ),
    .SUM(\s$743 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_72_0 (.A(pp_row72_11),
    .B(pp_row72_12),
    .CIN(pp_row72_13),
    .COUT(\c$744 ),
    .SUM(\s$745 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_72_1 (.A(pp_row72_14),
    .B(pp_row72_15),
    .CIN(pp_row72_16),
    .COUT(\c$746 ),
    .SUM(\s$747 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_72_2 (.A(pp_row72_17),
    .B(pp_row72_18),
    .CIN(pp_row72_19),
    .COUT(\c$748 ),
    .SUM(\s$749 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_72_3 (.A(pp_row72_20),
    .B(pp_row72_21),
    .CIN(pp_row72_22),
    .COUT(\c$750 ),
    .SUM(\s$751 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_72_4 (.A(pp_row72_23),
    .B(pp_row72_24),
    .CIN(pp_row72_25),
    .COUT(\c$752 ),
    .SUM(\s$753 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_72_5 (.A(pp_row72_26),
    .B(pp_row72_27),
    .CIN(pp_row72_28),
    .COUT(\c$754 ),
    .SUM(\s$755 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_72_6 (.A(pp_row72_29),
    .B(pp_row72_30),
    .CIN(\c$164 ),
    .COUT(\c$756 ),
    .SUM(\s$757 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_72_7 (.A(\c$166 ),
    .B(\c$168 ),
    .CIN(\c$170 ),
    .COUT(\c$758 ),
    .SUM(\s$759 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_72_8 (.A(\s$173 ),
    .B(\s$175 ),
    .CIN(\s$177 ),
    .COUT(\c$760 ),
    .SUM(\s$761 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_73_0 (.A(pp_row73_9),
    .B(pp_row73_10),
    .CIN(pp_row73_11),
    .COUT(\c$762 ),
    .SUM(\s$763 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_73_1 (.A(pp_row73_12),
    .B(pp_row73_13),
    .CIN(pp_row73_14),
    .COUT(\c$764 ),
    .SUM(\s$765 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_73_2 (.A(pp_row73_15),
    .B(pp_row73_16),
    .CIN(pp_row73_17),
    .COUT(\c$766 ),
    .SUM(\s$767 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_73_3 (.A(pp_row73_18),
    .B(pp_row73_19),
    .CIN(pp_row73_20),
    .COUT(\c$768 ),
    .SUM(\s$769 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_73_4 (.A(pp_row73_21),
    .B(pp_row73_22),
    .CIN(pp_row73_23),
    .COUT(\c$770 ),
    .SUM(\s$771 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_73_5 (.A(pp_row73_24),
    .B(pp_row73_25),
    .CIN(pp_row73_26),
    .COUT(\c$772 ),
    .SUM(\s$773 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_73_6 (.A(pp_row73_27),
    .B(pp_row73_28),
    .CIN(pp_row73_29),
    .COUT(\c$774 ),
    .SUM(\s$775 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_73_7 (.A(\c$172 ),
    .B(\c$174 ),
    .CIN(\c$176 ),
    .COUT(\c$776 ),
    .SUM(\s$777 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_73_8 (.A(\c$178 ),
    .B(\s$181 ),
    .CIN(\s$183 ),
    .COUT(\c$778 ),
    .SUM(\s$779 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_74_0 (.A(pp_row74_8),
    .B(pp_row74_9),
    .CIN(pp_row74_10),
    .COUT(\c$780 ),
    .SUM(\s$781 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_74_1 (.A(pp_row74_11),
    .B(pp_row74_12),
    .CIN(pp_row74_13),
    .COUT(\c$782 ),
    .SUM(\s$783 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_74_2 (.A(pp_row74_14),
    .B(pp_row74_15),
    .CIN(pp_row74_16),
    .COUT(\c$784 ),
    .SUM(\s$785 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_74_3 (.A(pp_row74_17),
    .B(pp_row74_18),
    .CIN(pp_row74_19),
    .COUT(\c$786 ),
    .SUM(\s$787 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_74_4 (.A(pp_row74_20),
    .B(pp_row74_21),
    .CIN(pp_row74_22),
    .COUT(\c$788 ),
    .SUM(\s$789 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_74_5 (.A(pp_row74_23),
    .B(pp_row74_24),
    .CIN(pp_row74_25),
    .COUT(\c$790 ),
    .SUM(\s$791 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_74_6 (.A(pp_row74_26),
    .B(pp_row74_27),
    .CIN(pp_row74_28),
    .COUT(\c$792 ),
    .SUM(\s$793 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_74_7 (.A(pp_row74_29),
    .B(\c$180 ),
    .CIN(\c$182 ),
    .COUT(\c$794 ),
    .SUM(\s$795 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_74_8 (.A(\c$184 ),
    .B(\s$187 ),
    .CIN(\s$189 ),
    .COUT(\c$796 ),
    .SUM(\s$797 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_75_0 (.A(pp_row75_6),
    .B(pp_row75_7),
    .CIN(pp_row75_8),
    .COUT(\c$798 ),
    .SUM(\s$799 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_75_1 (.A(pp_row75_9),
    .B(pp_row75_10),
    .CIN(pp_row75_11),
    .COUT(\c$800 ),
    .SUM(\s$801 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_75_2 (.A(pp_row75_12),
    .B(pp_row75_13),
    .CIN(pp_row75_14),
    .COUT(\c$802 ),
    .SUM(\s$803 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_75_3 (.A(pp_row75_15),
    .B(pp_row75_16),
    .CIN(pp_row75_17),
    .COUT(\c$804 ),
    .SUM(\s$805 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_75_4 (.A(pp_row75_18),
    .B(pp_row75_19),
    .CIN(pp_row75_20),
    .COUT(\c$806 ),
    .SUM(\s$807 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_75_5 (.A(pp_row75_21),
    .B(pp_row75_22),
    .CIN(pp_row75_23),
    .COUT(\c$808 ),
    .SUM(\s$809 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_75_6 (.A(pp_row75_24),
    .B(pp_row75_25),
    .CIN(pp_row75_26),
    .COUT(\c$810 ),
    .SUM(\s$811 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_75_7 (.A(pp_row75_27),
    .B(pp_row75_28),
    .CIN(\c$186 ),
    .COUT(\c$812 ),
    .SUM(\s$813 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_75_8 (.A(\c$188 ),
    .B(\c$190 ),
    .CIN(\s$193 ),
    .COUT(\c$814 ),
    .SUM(\s$815 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_76_0 (.A(pp_row76_5),
    .B(pp_row76_6),
    .CIN(pp_row76_7),
    .COUT(\c$816 ),
    .SUM(\s$817 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_76_1 (.A(pp_row76_8),
    .B(pp_row76_9),
    .CIN(pp_row76_10),
    .COUT(\c$818 ),
    .SUM(\s$819 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_76_2 (.A(pp_row76_11),
    .B(pp_row76_12),
    .CIN(pp_row76_13),
    .COUT(\c$820 ),
    .SUM(\s$821 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_76_3 (.A(pp_row76_14),
    .B(pp_row76_15),
    .CIN(pp_row76_16),
    .COUT(\c$822 ),
    .SUM(\s$823 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_76_4 (.A(pp_row76_17),
    .B(pp_row76_18),
    .CIN(pp_row76_19),
    .COUT(\c$824 ),
    .SUM(\s$825 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_76_5 (.A(pp_row76_20),
    .B(pp_row76_21),
    .CIN(pp_row76_22),
    .COUT(\c$826 ),
    .SUM(\s$827 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_76_6 (.A(pp_row76_23),
    .B(pp_row76_24),
    .CIN(pp_row76_25),
    .COUT(\c$828 ),
    .SUM(\s$829 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_76_7 (.A(pp_row76_26),
    .B(pp_row76_27),
    .CIN(pp_row76_28),
    .COUT(\c$830 ),
    .SUM(\s$831 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_76_8 (.A(\c$192 ),
    .B(\c$194 ),
    .CIN(\s$197 ),
    .COUT(\c$832 ),
    .SUM(\s$833 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_77_0 (.A(pp_row77_3),
    .B(pp_row77_4),
    .CIN(pp_row77_5),
    .COUT(\c$834 ),
    .SUM(\s$835 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_77_1 (.A(pp_row77_6),
    .B(pp_row77_7),
    .CIN(pp_row77_8),
    .COUT(\c$836 ),
    .SUM(\s$837 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_77_2 (.A(pp_row77_9),
    .B(pp_row77_10),
    .CIN(pp_row77_11),
    .COUT(\c$838 ),
    .SUM(\s$839 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_77_3 (.A(pp_row77_12),
    .B(pp_row77_13),
    .CIN(pp_row77_14),
    .COUT(\c$840 ),
    .SUM(\s$841 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_77_4 (.A(pp_row77_15),
    .B(pp_row77_16),
    .CIN(pp_row77_17),
    .COUT(\c$842 ),
    .SUM(\s$843 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_77_5 (.A(pp_row77_18),
    .B(pp_row77_19),
    .CIN(pp_row77_20),
    .COUT(\c$844 ),
    .SUM(\s$845 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_77_6 (.A(pp_row77_21),
    .B(pp_row77_22),
    .CIN(pp_row77_23),
    .COUT(\c$846 ),
    .SUM(\s$847 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_77_7 (.A(pp_row77_24),
    .B(pp_row77_25),
    .CIN(pp_row77_26),
    .COUT(\c$848 ),
    .SUM(\s$849 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_77_8 (.A(pp_row77_27),
    .B(\c$196 ),
    .CIN(\c$198 ),
    .COUT(\c$850 ),
    .SUM(\s$851 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_78_0 (.A(pp_row78_2),
    .B(pp_row78_3),
    .CIN(pp_row78_4),
    .COUT(\c$852 ),
    .SUM(\s$853 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_78_1 (.A(pp_row78_5),
    .B(pp_row78_6),
    .CIN(pp_row78_7),
    .COUT(\c$854 ),
    .SUM(\s$855 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_78_2 (.A(pp_row78_8),
    .B(pp_row78_9),
    .CIN(pp_row78_10),
    .COUT(\c$856 ),
    .SUM(\s$857 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_78_3 (.A(pp_row78_11),
    .B(pp_row78_12),
    .CIN(pp_row78_13),
    .COUT(\c$858 ),
    .SUM(\s$859 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_78_4 (.A(pp_row78_14),
    .B(pp_row78_15),
    .CIN(pp_row78_16),
    .COUT(\c$860 ),
    .SUM(\s$861 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_78_5 (.A(pp_row78_17),
    .B(pp_row78_18),
    .CIN(pp_row78_19),
    .COUT(\c$862 ),
    .SUM(\s$863 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_78_6 (.A(pp_row78_20),
    .B(pp_row78_21),
    .CIN(pp_row78_22),
    .COUT(\c$864 ),
    .SUM(\s$865 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_78_7 (.A(pp_row78_23),
    .B(pp_row78_24),
    .CIN(pp_row78_25),
    .COUT(\c$866 ),
    .SUM(\s$867 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_78_8 (.A(pp_row78_26),
    .B(pp_row78_27),
    .CIN(\c$200 ),
    .COUT(\c$868 ),
    .SUM(\s$869 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_79_0 (.A(pp_row79_0),
    .B(pp_row79_1),
    .CIN(pp_row79_2),
    .COUT(\c$870 ),
    .SUM(\s$871 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_79_1 (.A(pp_row79_3),
    .B(pp_row79_4),
    .CIN(pp_row79_5),
    .COUT(\c$872 ),
    .SUM(\s$873 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_79_2 (.A(pp_row79_6),
    .B(pp_row79_7),
    .CIN(pp_row79_8),
    .COUT(\c$874 ),
    .SUM(\s$875 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_79_3 (.A(pp_row79_9),
    .B(pp_row79_10),
    .CIN(pp_row79_11),
    .COUT(\c$876 ),
    .SUM(\s$877 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_79_4 (.A(pp_row79_12),
    .B(pp_row79_13),
    .CIN(pp_row79_14),
    .COUT(\c$878 ),
    .SUM(\s$879 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_79_5 (.A(pp_row79_15),
    .B(pp_row79_16),
    .CIN(pp_row79_17),
    .COUT(\c$880 ),
    .SUM(\s$881 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_79_6 (.A(pp_row79_18),
    .B(pp_row79_19),
    .CIN(pp_row79_20),
    .COUT(\c$882 ),
    .SUM(\s$883 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_79_7 (.A(pp_row79_21),
    .B(pp_row79_22),
    .CIN(pp_row79_23),
    .COUT(\c$884 ),
    .SUM(\s$885 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_79_8 (.A(pp_row79_24),
    .B(pp_row79_25),
    .CIN(pp_row79_26),
    .COUT(\c$886 ),
    .SUM(\s$887 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_80_0 (.A(net1896),
    .B(pp_row80_1),
    .CIN(pp_row80_2),
    .COUT(\c$888 ),
    .SUM(\s$889 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_80_1 (.A(pp_row80_3),
    .B(pp_row80_4),
    .CIN(pp_row80_5),
    .COUT(\c$890 ),
    .SUM(\s$891 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_80_2 (.A(pp_row80_6),
    .B(pp_row80_7),
    .CIN(pp_row80_8),
    .COUT(\c$892 ),
    .SUM(\s$893 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_80_3 (.A(pp_row80_9),
    .B(pp_row80_10),
    .CIN(pp_row80_11),
    .COUT(\c$894 ),
    .SUM(\s$895 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_80_4 (.A(pp_row80_12),
    .B(pp_row80_13),
    .CIN(pp_row80_14),
    .COUT(\c$896 ),
    .SUM(\s$897 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_80_5 (.A(pp_row80_15),
    .B(pp_row80_16),
    .CIN(pp_row80_17),
    .COUT(\c$898 ),
    .SUM(\s$899 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_80_6 (.A(pp_row80_18),
    .B(pp_row80_19),
    .CIN(pp_row80_20),
    .COUT(\c$900 ),
    .SUM(\s$901 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_80_7 (.A(pp_row80_21),
    .B(pp_row80_22),
    .CIN(pp_row80_23),
    .COUT(\c$902 ),
    .SUM(\s$903 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_81_0 (.A(pp_row81_0),
    .B(pp_row81_1),
    .CIN(pp_row81_2),
    .COUT(\c$906 ),
    .SUM(\s$907 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_81_1 (.A(pp_row81_3),
    .B(pp_row81_4),
    .CIN(pp_row81_5),
    .COUT(\c$908 ),
    .SUM(\s$909 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_81_2 (.A(pp_row81_6),
    .B(pp_row81_7),
    .CIN(pp_row81_8),
    .COUT(\c$910 ),
    .SUM(\s$911 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_81_3 (.A(pp_row81_9),
    .B(pp_row81_10),
    .CIN(pp_row81_11),
    .COUT(\c$912 ),
    .SUM(\s$913 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_81_4 (.A(pp_row81_12),
    .B(pp_row81_13),
    .CIN(pp_row81_14),
    .COUT(\c$914 ),
    .SUM(\s$915 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_81_5 (.A(pp_row81_15),
    .B(pp_row81_16),
    .CIN(pp_row81_17),
    .COUT(\c$916 ),
    .SUM(\s$917 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_81_6 (.A(pp_row81_18),
    .B(pp_row81_19),
    .CIN(pp_row81_20),
    .COUT(\c$918 ),
    .SUM(\s$919 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_81_7 (.A(pp_row81_21),
    .B(pp_row81_22),
    .CIN(pp_row81_23),
    .COUT(\c$920 ),
    .SUM(\s$921 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_82_0 (.A(net1897),
    .B(pp_row82_1),
    .CIN(pp_row82_2),
    .COUT(\c$922 ),
    .SUM(\s$923 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_82_1 (.A(pp_row82_3),
    .B(pp_row82_4),
    .CIN(pp_row82_5),
    .COUT(\c$924 ),
    .SUM(\s$925 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_82_2 (.A(pp_row82_6),
    .B(pp_row82_7),
    .CIN(pp_row82_8),
    .COUT(\c$926 ),
    .SUM(\s$927 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_82_3 (.A(pp_row82_9),
    .B(pp_row82_10),
    .CIN(pp_row82_11),
    .COUT(\c$928 ),
    .SUM(\s$929 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_82_4 (.A(pp_row82_12),
    .B(pp_row82_13),
    .CIN(pp_row82_14),
    .COUT(\c$930 ),
    .SUM(\s$931 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_82_5 (.A(pp_row82_15),
    .B(pp_row82_16),
    .CIN(pp_row82_17),
    .COUT(\c$932 ),
    .SUM(\s$933 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_82_6 (.A(pp_row82_18),
    .B(pp_row82_19),
    .CIN(pp_row82_20),
    .COUT(\c$934 ),
    .SUM(\s$935 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_83_0 (.A(pp_row83_0),
    .B(pp_row83_1),
    .CIN(pp_row83_2),
    .COUT(\c$938 ),
    .SUM(\s$939 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_83_1 (.A(pp_row83_3),
    .B(pp_row83_4),
    .CIN(pp_row83_5),
    .COUT(\c$940 ),
    .SUM(\s$941 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_83_2 (.A(pp_row83_6),
    .B(pp_row83_7),
    .CIN(pp_row83_8),
    .COUT(\c$942 ),
    .SUM(\s$943 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_83_3 (.A(pp_row83_9),
    .B(pp_row83_10),
    .CIN(pp_row83_11),
    .COUT(\c$944 ),
    .SUM(\s$945 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_83_4 (.A(pp_row83_12),
    .B(pp_row83_13),
    .CIN(pp_row83_14),
    .COUT(\c$946 ),
    .SUM(\s$947 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_83_5 (.A(pp_row83_15),
    .B(pp_row83_16),
    .CIN(pp_row83_17),
    .COUT(\c$948 ),
    .SUM(\s$949 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_83_6 (.A(pp_row83_18),
    .B(pp_row83_19),
    .CIN(pp_row83_20),
    .COUT(\c$950 ),
    .SUM(\s$951 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_84_0 (.A(net1898),
    .B(pp_row84_1),
    .CIN(pp_row84_2),
    .COUT(\c$952 ),
    .SUM(\s$953 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_84_1 (.A(pp_row84_3),
    .B(pp_row84_4),
    .CIN(pp_row84_5),
    .COUT(\c$954 ),
    .SUM(\s$955 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_84_2 (.A(pp_row84_6),
    .B(pp_row84_7),
    .CIN(pp_row84_8),
    .COUT(\c$956 ),
    .SUM(\s$957 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_84_3 (.A(pp_row84_9),
    .B(pp_row84_10),
    .CIN(pp_row84_11),
    .COUT(\c$958 ),
    .SUM(\s$959 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_84_4 (.A(pp_row84_12),
    .B(pp_row84_13),
    .CIN(pp_row84_14),
    .COUT(\c$960 ),
    .SUM(\s$961 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_84_5 (.A(pp_row84_15),
    .B(pp_row84_16),
    .CIN(pp_row84_17),
    .COUT(\c$962 ),
    .SUM(\s$963 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_85_0 (.A(pp_row85_0),
    .B(pp_row85_1),
    .CIN(pp_row85_2),
    .COUT(\c$966 ),
    .SUM(\s$967 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_85_1 (.A(pp_row85_3),
    .B(pp_row85_4),
    .CIN(pp_row85_5),
    .COUT(\c$968 ),
    .SUM(\s$969 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_85_2 (.A(pp_row85_6),
    .B(pp_row85_7),
    .CIN(pp_row85_8),
    .COUT(\c$970 ),
    .SUM(\s$971 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_85_3 (.A(pp_row85_9),
    .B(pp_row85_10),
    .CIN(pp_row85_11),
    .COUT(\c$972 ),
    .SUM(\s$973 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_85_4 (.A(pp_row85_12),
    .B(pp_row85_13),
    .CIN(pp_row85_14),
    .COUT(\c$974 ),
    .SUM(\s$975 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_85_5 (.A(pp_row85_15),
    .B(pp_row85_16),
    .CIN(pp_row85_17),
    .COUT(\c$976 ),
    .SUM(\s$977 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_86_0 (.A(net1899),
    .B(pp_row86_1),
    .CIN(pp_row86_2),
    .COUT(\c$978 ),
    .SUM(\s$979 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_86_1 (.A(pp_row86_3),
    .B(pp_row86_4),
    .CIN(pp_row86_5),
    .COUT(\c$980 ),
    .SUM(\s$981 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_86_2 (.A(pp_row86_6),
    .B(pp_row86_7),
    .CIN(pp_row86_8),
    .COUT(\c$982 ),
    .SUM(\s$983 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_86_3 (.A(pp_row86_9),
    .B(pp_row86_10),
    .CIN(pp_row86_11),
    .COUT(\c$984 ),
    .SUM(\s$985 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_86_4 (.A(pp_row86_12),
    .B(pp_row86_13),
    .CIN(pp_row86_14),
    .COUT(\c$986 ),
    .SUM(\s$987 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_87_0 (.A(pp_row87_0),
    .B(pp_row87_1),
    .CIN(pp_row87_2),
    .COUT(\c$990 ),
    .SUM(\s$991 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_87_1 (.A(pp_row87_3),
    .B(pp_row87_4),
    .CIN(pp_row87_5),
    .COUT(\c$992 ),
    .SUM(\s$993 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_87_2 (.A(pp_row87_6),
    .B(pp_row87_7),
    .CIN(pp_row87_8),
    .COUT(\c$994 ),
    .SUM(\s$995 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_87_3 (.A(pp_row87_9),
    .B(pp_row87_10),
    .CIN(pp_row87_11),
    .COUT(\c$996 ),
    .SUM(\s$997 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_87_4 (.A(pp_row87_12),
    .B(pp_row87_13),
    .CIN(pp_row87_14),
    .COUT(\c$998 ),
    .SUM(\s$999 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_88_0 (.A(net1900),
    .B(pp_row88_1),
    .CIN(pp_row88_2),
    .COUT(\c$1000 ),
    .SUM(\s$1001 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_88_1 (.A(pp_row88_3),
    .B(pp_row88_4),
    .CIN(pp_row88_5),
    .COUT(\c$1002 ),
    .SUM(\s$1003 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_88_2 (.A(pp_row88_6),
    .B(pp_row88_7),
    .CIN(pp_row88_8),
    .COUT(\c$1004 ),
    .SUM(\s$1005 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_88_3 (.A(pp_row88_9),
    .B(pp_row88_10),
    .CIN(pp_row88_11),
    .COUT(\c$1006 ),
    .SUM(\s$1007 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_1_89_0 (.A(pp_row89_0),
    .B(pp_row89_1),
    .CIN(pp_row89_2),
    .COUT(\c$1010 ),
    .SUM(\s$1011 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_89_1 (.A(pp_row89_3),
    .B(pp_row89_4),
    .CIN(pp_row89_5),
    .COUT(\c$1012 ),
    .SUM(\s$1013 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_89_2 (.A(pp_row89_6),
    .B(pp_row89_7),
    .CIN(pp_row89_8),
    .COUT(\c$1014 ),
    .SUM(\s$1015 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_89_3 (.A(pp_row89_9),
    .B(pp_row89_10),
    .CIN(pp_row89_11),
    .COUT(\c$1016 ),
    .SUM(\s$1017 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_90_0 (.A(net1901),
    .B(pp_row90_1),
    .CIN(pp_row90_2),
    .COUT(\c$1018 ),
    .SUM(\s$1019 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_90_1 (.A(pp_row90_3),
    .B(pp_row90_4),
    .CIN(pp_row90_5),
    .COUT(\c$1020 ),
    .SUM(\s$1021 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_90_2 (.A(pp_row90_6),
    .B(pp_row90_7),
    .CIN(pp_row90_8),
    .COUT(\c$1022 ),
    .SUM(\s$1023 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_91_0 (.A(pp_row91_0),
    .B(pp_row91_1),
    .CIN(pp_row91_2),
    .COUT(\c$1026 ),
    .SUM(\s$1027 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_91_1 (.A(pp_row91_3),
    .B(pp_row91_4),
    .CIN(pp_row91_5),
    .COUT(\c$1028 ),
    .SUM(\s$1029 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_91_2 (.A(pp_row91_6),
    .B(pp_row91_7),
    .CIN(pp_row91_8),
    .COUT(\c$1030 ),
    .SUM(\s$1031 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_92_0 (.A(net1902),
    .B(pp_row92_1),
    .CIN(pp_row92_2),
    .COUT(\c$1032 ),
    .SUM(\s$1033 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_92_1 (.A(pp_row92_3),
    .B(pp_row92_4),
    .CIN(pp_row92_5),
    .COUT(\c$1034 ),
    .SUM(\s$1035 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_93_0 (.A(pp_row93_0),
    .B(pp_row93_1),
    .CIN(pp_row93_2),
    .COUT(\c$1038 ),
    .SUM(\s$1039 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_93_1 (.A(pp_row93_3),
    .B(pp_row93_4),
    .CIN(pp_row93_5),
    .COUT(\c$1040 ),
    .SUM(\s$1041 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_94_0 (.A(net1903),
    .B(pp_row94_1),
    .CIN(pp_row94_2),
    .COUT(\c$1042 ),
    .SUM(\s$1043 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_1_95_0 (.A(pp_row95_0),
    .B(pp_row95_1),
    .CIN(pp_row95_2),
    .COUT(\c$1046 ),
    .SUM(\s$1047 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_100_0 (.A(net1904),
    .B(pp_row100_1),
    .CIN(pp_row100_2),
    .COUT(\c$1924 ),
    .SUM(\s$1925 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_100_1 (.A(pp_row100_3),
    .B(pp_row100_4),
    .CIN(pp_row100_5),
    .COUT(\c$1926 ),
    .SUM(\s$1927 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_100_2 (.A(pp_row100_6),
    .B(pp_row100_7),
    .CIN(pp_row100_8),
    .COUT(\c$1928 ),
    .SUM(\s$1929 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_100_3 (.A(pp_row100_9),
    .B(pp_row100_10),
    .CIN(pp_row100_11),
    .COUT(\c$1930 ),
    .SUM(\s$1931 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_101_0 (.A(pp_row101_0),
    .B(pp_row101_1),
    .CIN(pp_row101_2),
    .COUT(\c$1934 ),
    .SUM(\s$1935 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_101_1 (.A(pp_row101_3),
    .B(pp_row101_4),
    .CIN(pp_row101_5),
    .COUT(\c$1936 ),
    .SUM(\s$1937 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_101_2 (.A(pp_row101_6),
    .B(pp_row101_7),
    .CIN(pp_row101_8),
    .COUT(\c$1938 ),
    .SUM(\s$1939 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_101_3 (.A(pp_row101_9),
    .B(pp_row101_10),
    .CIN(pp_row101_11),
    .COUT(\c$1940 ),
    .SUM(\s$1941 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_102_0 (.A(net1905),
    .B(pp_row102_1),
    .CIN(pp_row102_2),
    .COUT(\c$1942 ),
    .SUM(\s$1943 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_102_1 (.A(pp_row102_3),
    .B(pp_row102_4),
    .CIN(pp_row102_5),
    .COUT(\c$1944 ),
    .SUM(\s$1945 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_102_2 (.A(pp_row102_6),
    .B(pp_row102_7),
    .CIN(pp_row102_8),
    .COUT(\c$1946 ),
    .SUM(\s$1947 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_103_0 (.A(pp_row103_0),
    .B(pp_row103_1),
    .CIN(pp_row103_2),
    .COUT(\c$1950 ),
    .SUM(\s$1951 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_103_1 (.A(pp_row103_3),
    .B(pp_row103_4),
    .CIN(pp_row103_5),
    .COUT(\c$1952 ),
    .SUM(\s$1953 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_103_2 (.A(pp_row103_6),
    .B(pp_row103_7),
    .CIN(pp_row103_8),
    .COUT(\c$1954 ),
    .SUM(\s$1955 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_104_0 (.A(net1906),
    .B(pp_row104_1),
    .CIN(pp_row104_2),
    .COUT(\c$1956 ),
    .SUM(\s$1957 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_104_1 (.A(pp_row104_3),
    .B(pp_row104_4),
    .CIN(pp_row104_5),
    .COUT(\c$1958 ),
    .SUM(\s$1959 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_105_0 (.A(pp_row105_0),
    .B(pp_row105_1),
    .CIN(pp_row105_2),
    .COUT(\c$1962 ),
    .SUM(\s$1963 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_105_1 (.A(pp_row105_3),
    .B(pp_row105_4),
    .CIN(pp_row105_5),
    .COUT(\c$1964 ),
    .SUM(\s$1965 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_106_0 (.A(net1907),
    .B(pp_row106_1),
    .CIN(pp_row106_2),
    .COUT(\c$1966 ),
    .SUM(\s$1967 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_107_0 (.A(pp_row107_0),
    .B(pp_row107_1),
    .CIN(pp_row107_2),
    .COUT(\c$1970 ),
    .SUM(\s$1971 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_24_0 (.A(pp_row24_0),
    .B(pp_row24_1),
    .CIN(pp_row24_2),
    .COUT(\c$1054 ),
    .SUM(\s$1055 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_25_0 (.A(pp_row25_0),
    .B(pp_row25_1),
    .CIN(pp_row25_2),
    .COUT(\c$1058 ),
    .SUM(\s$1059 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_26_0 (.A(pp_row26_0),
    .B(pp_row26_1),
    .CIN(pp_row26_2),
    .COUT(\c$1062 ),
    .SUM(\s$1063 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_26_1 (.A(pp_row26_3),
    .B(pp_row26_4),
    .CIN(pp_row26_5),
    .COUT(\c$1064 ),
    .SUM(\s$1065 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_27_0 (.A(pp_row27_0),
    .B(pp_row27_1),
    .CIN(pp_row27_2),
    .COUT(\c$1068 ),
    .SUM(\s$1069 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_27_1 (.A(pp_row27_3),
    .B(pp_row27_4),
    .CIN(pp_row27_5),
    .COUT(\c$1070 ),
    .SUM(\s$1071 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_28_0 (.A(pp_row28_0),
    .B(pp_row28_1),
    .CIN(pp_row28_2),
    .COUT(\c$1074 ),
    .SUM(\s$1075 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_28_1 (.A(pp_row28_3),
    .B(pp_row28_4),
    .CIN(pp_row28_5),
    .COUT(\c$1076 ),
    .SUM(\s$1077 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_28_2 (.A(pp_row28_6),
    .B(pp_row28_7),
    .CIN(pp_row28_8),
    .COUT(\c$1078 ),
    .SUM(\s$1079 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_29_0 (.A(pp_row29_0),
    .B(pp_row29_1),
    .CIN(pp_row29_2),
    .COUT(\c$1082 ),
    .SUM(\s$1083 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_29_1 (.A(pp_row29_3),
    .B(pp_row29_4),
    .CIN(pp_row29_5),
    .COUT(\c$1084 ),
    .SUM(\s$1085 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_29_2 (.A(pp_row29_6),
    .B(pp_row29_7),
    .CIN(pp_row29_8),
    .COUT(\c$1086 ),
    .SUM(\s$1087 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_30_0 (.A(pp_row30_0),
    .B(pp_row30_1),
    .CIN(pp_row30_2),
    .COUT(\c$1090 ),
    .SUM(\s$1091 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_30_1 (.A(pp_row30_3),
    .B(pp_row30_4),
    .CIN(pp_row30_5),
    .COUT(\c$1092 ),
    .SUM(\s$1093 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_30_2 (.A(pp_row30_6),
    .B(pp_row30_7),
    .CIN(pp_row30_8),
    .COUT(\c$1094 ),
    .SUM(\s$1095 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_30_3 (.A(pp_row30_9),
    .B(pp_row30_10),
    .CIN(pp_row30_11),
    .COUT(\c$1096 ),
    .SUM(\s$1097 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_31_0 (.A(pp_row31_0),
    .B(pp_row31_1),
    .CIN(pp_row31_2),
    .COUT(\c$1100 ),
    .SUM(\s$1101 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_31_1 (.A(pp_row31_3),
    .B(pp_row31_4),
    .CIN(pp_row31_5),
    .COUT(\c$1102 ),
    .SUM(\s$1103 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_31_2 (.A(pp_row31_6),
    .B(pp_row31_7),
    .CIN(pp_row31_8),
    .COUT(\c$1104 ),
    .SUM(\s$1105 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_31_3 (.A(pp_row31_9),
    .B(pp_row31_10),
    .CIN(pp_row31_11),
    .COUT(\c$1106 ),
    .SUM(\s$1107 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_32_0 (.A(pp_row32_0),
    .B(pp_row32_1),
    .CIN(pp_row32_2),
    .COUT(\c$1110 ),
    .SUM(\s$1111 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_32_1 (.A(pp_row32_3),
    .B(pp_row32_4),
    .CIN(pp_row32_5),
    .COUT(\c$1112 ),
    .SUM(\s$1113 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_32_2 (.A(pp_row32_6),
    .B(pp_row32_7),
    .CIN(pp_row32_8),
    .COUT(\c$1114 ),
    .SUM(\s$1115 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_32_3 (.A(pp_row32_9),
    .B(pp_row32_10),
    .CIN(pp_row32_11),
    .COUT(\c$1116 ),
    .SUM(\s$1117 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_32_4 (.A(pp_row32_12),
    .B(pp_row32_13),
    .CIN(pp_row32_14),
    .COUT(\c$1118 ),
    .SUM(\s$1119 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_33_0 (.A(pp_row33_0),
    .B(pp_row33_1),
    .CIN(pp_row33_2),
    .COUT(\c$1122 ),
    .SUM(\s$1123 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_33_1 (.A(pp_row33_3),
    .B(pp_row33_4),
    .CIN(pp_row33_5),
    .COUT(\c$1124 ),
    .SUM(\s$1125 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_33_2 (.A(pp_row33_6),
    .B(pp_row33_7),
    .CIN(pp_row33_8),
    .COUT(\c$1126 ),
    .SUM(\s$1127 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_33_3 (.A(pp_row33_9),
    .B(pp_row33_10),
    .CIN(pp_row33_11),
    .COUT(\c$1128 ),
    .SUM(\s$1129 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_33_4 (.A(pp_row33_12),
    .B(pp_row33_13),
    .CIN(pp_row33_14),
    .COUT(\c$1130 ),
    .SUM(\s$1131 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_34_0 (.A(pp_row34_2),
    .B(pp_row34_3),
    .CIN(pp_row34_4),
    .COUT(\c$1134 ),
    .SUM(\s$1135 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_34_1 (.A(pp_row34_5),
    .B(pp_row34_6),
    .CIN(pp_row34_7),
    .COUT(\c$1136 ),
    .SUM(\s$1137 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_34_2 (.A(pp_row34_8),
    .B(pp_row34_9),
    .CIN(pp_row34_10),
    .COUT(\c$1138 ),
    .SUM(\s$1139 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_34_3 (.A(pp_row34_11),
    .B(pp_row34_12),
    .CIN(pp_row34_13),
    .COUT(\c$1140 ),
    .SUM(\s$1141 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_34_4 (.A(pp_row34_14),
    .B(pp_row34_15),
    .CIN(pp_row34_16),
    .COUT(\c$1142 ),
    .SUM(\s$1143 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_34_5 (.A(pp_row34_17),
    .B(pp_row34_18),
    .CIN(pp_row34_19),
    .COUT(\c$1144 ),
    .SUM(\s$1145 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_35_0 (.A(pp_row35_2),
    .B(pp_row35_3),
    .CIN(pp_row35_4),
    .COUT(\c$1146 ),
    .SUM(\s$1147 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_35_1 (.A(pp_row35_5),
    .B(pp_row35_6),
    .CIN(pp_row35_7),
    .COUT(\c$1148 ),
    .SUM(\s$1149 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_35_2 (.A(pp_row35_8),
    .B(pp_row35_9),
    .CIN(pp_row35_10),
    .COUT(\c$1150 ),
    .SUM(\s$1151 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_35_3 (.A(pp_row35_11),
    .B(pp_row35_12),
    .CIN(pp_row35_13),
    .COUT(\c$1152 ),
    .SUM(\s$1153 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_35_4 (.A(pp_row35_14),
    .B(pp_row35_15),
    .CIN(pp_row35_16),
    .COUT(\c$1154 ),
    .SUM(\s$1155 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_35_5 (.A(pp_row35_17),
    .B(pp_row35_18),
    .CIN(\c$204 ),
    .COUT(\c$1156 ),
    .SUM(\s$1157 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_36_0 (.A(pp_row36_5),
    .B(pp_row36_6),
    .CIN(pp_row36_7),
    .COUT(\c$1158 ),
    .SUM(\s$1159 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_36_1 (.A(pp_row36_8),
    .B(pp_row36_9),
    .CIN(pp_row36_10),
    .COUT(\c$1160 ),
    .SUM(\s$1161 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_36_2 (.A(pp_row36_11),
    .B(pp_row36_12),
    .CIN(pp_row36_13),
    .COUT(\c$1162 ),
    .SUM(\s$1163 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_36_3 (.A(pp_row36_14),
    .B(pp_row36_15),
    .CIN(pp_row36_16),
    .COUT(\c$1164 ),
    .SUM(\s$1165 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_36_4 (.A(pp_row36_17),
    .B(pp_row36_18),
    .CIN(pp_row36_19),
    .COUT(\c$1166 ),
    .SUM(\s$1167 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_36_5 (.A(pp_row36_20),
    .B(\c$206 ),
    .CIN(\s$209 ),
    .COUT(\c$1168 ),
    .SUM(\s$1169 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_37_0 (.A(pp_row37_5),
    .B(pp_row37_6),
    .CIN(pp_row37_7),
    .COUT(\c$1170 ),
    .SUM(\s$1171 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_37_1 (.A(pp_row37_8),
    .B(pp_row37_9),
    .CIN(pp_row37_10),
    .COUT(\c$1172 ),
    .SUM(\s$1173 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_37_2 (.A(pp_row37_11),
    .B(pp_row37_12),
    .CIN(pp_row37_13),
    .COUT(\c$1174 ),
    .SUM(\s$1175 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_37_3 (.A(pp_row37_14),
    .B(pp_row37_15),
    .CIN(pp_row37_16),
    .COUT(\c$1176 ),
    .SUM(\s$1177 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_37_4 (.A(pp_row37_17),
    .B(pp_row37_18),
    .CIN(pp_row37_19),
    .COUT(\c$1178 ),
    .SUM(\s$1179 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_37_5 (.A(\c$208 ),
    .B(\c$210 ),
    .CIN(\s$213 ),
    .COUT(\c$1180 ),
    .SUM(\s$1181 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_38_0 (.A(pp_row38_8),
    .B(pp_row38_9),
    .CIN(pp_row38_10),
    .COUT(\c$1182 ),
    .SUM(\s$1183 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_38_1 (.A(pp_row38_11),
    .B(pp_row38_12),
    .CIN(pp_row38_13),
    .COUT(\c$1184 ),
    .SUM(\s$1185 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_38_2 (.A(pp_row38_14),
    .B(pp_row38_15),
    .CIN(pp_row38_16),
    .COUT(\c$1186 ),
    .SUM(\s$1187 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_38_3 (.A(pp_row38_17),
    .B(pp_row38_18),
    .CIN(pp_row38_19),
    .COUT(\c$1188 ),
    .SUM(\s$1189 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_38_4 (.A(pp_row38_20),
    .B(pp_row38_21),
    .CIN(\c$212 ),
    .COUT(\c$1190 ),
    .SUM(\s$1191 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_38_5 (.A(\c$214 ),
    .B(\s$217 ),
    .CIN(\s$219 ),
    .COUT(\c$1192 ),
    .SUM(\s$1193 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_39_0 (.A(pp_row39_8),
    .B(pp_row39_9),
    .CIN(pp_row39_10),
    .COUT(\c$1194 ),
    .SUM(\s$1195 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_39_1 (.A(pp_row39_11),
    .B(pp_row39_12),
    .CIN(pp_row39_13),
    .COUT(\c$1196 ),
    .SUM(\s$1197 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_39_2 (.A(pp_row39_14),
    .B(pp_row39_15),
    .CIN(pp_row39_16),
    .COUT(\c$1198 ),
    .SUM(\s$1199 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_39_3 (.A(pp_row39_17),
    .B(pp_row39_18),
    .CIN(pp_row39_19),
    .COUT(\c$1200 ),
    .SUM(\s$1201 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_39_4 (.A(pp_row39_20),
    .B(\c$216 ),
    .CIN(\c$218 ),
    .COUT(\c$1202 ),
    .SUM(\s$1203 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_39_5 (.A(\c$220 ),
    .B(\s$223 ),
    .CIN(\s$225 ),
    .COUT(\c$1204 ),
    .SUM(\s$1205 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_40_0 (.A(pp_row40_11),
    .B(pp_row40_12),
    .CIN(pp_row40_13),
    .COUT(\c$1206 ),
    .SUM(\s$1207 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_40_1 (.A(pp_row40_14),
    .B(pp_row40_15),
    .CIN(pp_row40_16),
    .COUT(\c$1208 ),
    .SUM(\s$1209 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_40_2 (.A(pp_row40_17),
    .B(pp_row40_18),
    .CIN(pp_row40_19),
    .COUT(\c$1210 ),
    .SUM(\s$1211 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_40_3 (.A(pp_row40_20),
    .B(pp_row40_21),
    .CIN(pp_row40_22),
    .COUT(\c$1212 ),
    .SUM(\s$1213 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_40_4 (.A(\c$222 ),
    .B(\c$224 ),
    .CIN(\c$226 ),
    .COUT(\c$1214 ),
    .SUM(\s$1215 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_40_5 (.A(\s$229 ),
    .B(\s$231 ),
    .CIN(\s$233 ),
    .COUT(\c$1216 ),
    .SUM(\s$1217 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_41_0 (.A(pp_row41_11),
    .B(pp_row41_12),
    .CIN(pp_row41_13),
    .COUT(\c$1218 ),
    .SUM(\s$1219 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_41_1 (.A(pp_row41_14),
    .B(pp_row41_15),
    .CIN(pp_row41_16),
    .COUT(\c$1220 ),
    .SUM(\s$1221 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_41_2 (.A(pp_row41_17),
    .B(pp_row41_18),
    .CIN(pp_row41_19),
    .COUT(\c$1222 ),
    .SUM(\s$1223 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_41_3 (.A(pp_row41_20),
    .B(pp_row41_21),
    .CIN(\c$228 ),
    .COUT(\c$1224 ),
    .SUM(\s$1225 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_41_4 (.A(\c$230 ),
    .B(\c$232 ),
    .CIN(\c$234 ),
    .COUT(\c$1226 ),
    .SUM(\s$1227 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_41_5 (.A(\s$237 ),
    .B(\s$239 ),
    .CIN(\s$241 ),
    .COUT(\c$1228 ),
    .SUM(\s$1229 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_42_0 (.A(pp_row42_14),
    .B(pp_row42_15),
    .CIN(pp_row42_16),
    .COUT(\c$1230 ),
    .SUM(\s$1231 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_42_1 (.A(pp_row42_17),
    .B(pp_row42_18),
    .CIN(pp_row42_19),
    .COUT(\c$1232 ),
    .SUM(\s$1233 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_42_2 (.A(pp_row42_20),
    .B(pp_row42_21),
    .CIN(pp_row42_22),
    .COUT(\c$1234 ),
    .SUM(\s$1235 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_42_3 (.A(pp_row42_23),
    .B(\c$236 ),
    .CIN(\c$238 ),
    .COUT(\c$1236 ),
    .SUM(\s$1237 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_42_4 (.A(\c$240 ),
    .B(\c$242 ),
    .CIN(\s$245 ),
    .COUT(\c$1238 ),
    .SUM(\s$1239 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_42_5 (.A(\s$247 ),
    .B(\s$249 ),
    .CIN(\s$251 ),
    .COUT(\c$1240 ),
    .SUM(\s$1241 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_43_0 (.A(pp_row43_14),
    .B(pp_row43_15),
    .CIN(pp_row43_16),
    .COUT(\c$1242 ),
    .SUM(\s$1243 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_43_1 (.A(pp_row43_17),
    .B(pp_row43_18),
    .CIN(pp_row43_19),
    .COUT(\c$1244 ),
    .SUM(\s$1245 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_43_2 (.A(pp_row43_20),
    .B(pp_row43_21),
    .CIN(pp_row43_22),
    .COUT(\c$1246 ),
    .SUM(\s$1247 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_43_3 (.A(\c$244 ),
    .B(\c$246 ),
    .CIN(\c$248 ),
    .COUT(\c$1248 ),
    .SUM(\s$1249 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_43_4 (.A(\c$250 ),
    .B(\c$252 ),
    .CIN(\s$255 ),
    .COUT(\c$1250 ),
    .SUM(\s$1251 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_43_5 (.A(\s$257 ),
    .B(\s$259 ),
    .CIN(\s$261 ),
    .COUT(\c$1252 ),
    .SUM(\s$1253 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_44_0 (.A(pp_row44_17),
    .B(pp_row44_18),
    .CIN(pp_row44_19),
    .COUT(\c$1254 ),
    .SUM(\s$1255 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_44_1 (.A(pp_row44_20),
    .B(pp_row44_21),
    .CIN(pp_row44_22),
    .COUT(\c$1256 ),
    .SUM(\s$1257 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_44_2 (.A(pp_row44_23),
    .B(pp_row44_24),
    .CIN(\c$254 ),
    .COUT(\c$1258 ),
    .SUM(\s$1259 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_44_3 (.A(\c$256 ),
    .B(\c$258 ),
    .CIN(\c$260 ),
    .COUT(\c$1260 ),
    .SUM(\s$1261 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_44_4 (.A(\c$262 ),
    .B(\s$265 ),
    .CIN(\s$267 ),
    .COUT(\c$1262 ),
    .SUM(\s$1263 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_44_5 (.A(\s$269 ),
    .B(\s$271 ),
    .CIN(\s$273 ),
    .COUT(\c$1264 ),
    .SUM(\s$1265 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_45_0 (.A(pp_row45_17),
    .B(pp_row45_18),
    .CIN(pp_row45_19),
    .COUT(\c$1266 ),
    .SUM(\s$1267 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_45_1 (.A(pp_row45_20),
    .B(pp_row45_21),
    .CIN(pp_row45_22),
    .COUT(\c$1268 ),
    .SUM(\s$1269 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_45_2 (.A(pp_row45_23),
    .B(\c$264 ),
    .CIN(\c$266 ),
    .COUT(\c$1270 ),
    .SUM(\s$1271 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_45_3 (.A(\c$268 ),
    .B(\c$270 ),
    .CIN(\c$272 ),
    .COUT(\c$1272 ),
    .SUM(\s$1273 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_45_4 (.A(\c$274 ),
    .B(\s$277 ),
    .CIN(\s$279 ),
    .COUT(\c$1274 ),
    .SUM(\s$1275 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_45_5 (.A(\s$281 ),
    .B(\s$283 ),
    .CIN(\s$285 ),
    .COUT(\c$1276 ),
    .SUM(\s$1277 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_46_0 (.A(pp_row46_20),
    .B(pp_row46_21),
    .CIN(pp_row46_22),
    .COUT(\c$1278 ),
    .SUM(\s$1279 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_46_1 (.A(pp_row46_23),
    .B(pp_row46_24),
    .CIN(pp_row46_25),
    .COUT(\c$1280 ),
    .SUM(\s$1281 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_46_2 (.A(\c$276 ),
    .B(\c$278 ),
    .CIN(\c$280 ),
    .COUT(\c$1282 ),
    .SUM(\s$1283 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_46_3 (.A(\c$282 ),
    .B(\c$284 ),
    .CIN(\c$286 ),
    .COUT(\c$1284 ),
    .SUM(\s$1285 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_46_4 (.A(\s$289 ),
    .B(\s$291 ),
    .CIN(\s$293 ),
    .COUT(\c$1286 ),
    .SUM(\s$1287 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_46_5 (.A(\s$295 ),
    .B(\s$297 ),
    .CIN(\s$299 ),
    .COUT(\c$1288 ),
    .SUM(\s$1289 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_47_0 (.A(pp_row47_20),
    .B(pp_row47_21),
    .CIN(pp_row47_22),
    .COUT(\c$1290 ),
    .SUM(\s$1291 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_47_1 (.A(pp_row47_23),
    .B(pp_row47_24),
    .CIN(\c$288 ),
    .COUT(\c$1292 ),
    .SUM(\s$1293 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_47_2 (.A(\c$290 ),
    .B(\c$292 ),
    .CIN(\c$294 ),
    .COUT(\c$1294 ),
    .SUM(\s$1295 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_47_3 (.A(\c$296 ),
    .B(\c$298 ),
    .CIN(\c$300 ),
    .COUT(\c$1296 ),
    .SUM(\s$1297 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_47_4 (.A(\s$303 ),
    .B(\s$305 ),
    .CIN(\s$307 ),
    .COUT(\c$1298 ),
    .SUM(\s$1299 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_47_5 (.A(\s$309 ),
    .B(\s$311 ),
    .CIN(\s$313 ),
    .COUT(\c$1300 ),
    .SUM(\s$1301 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_48_0 (.A(pp_row48_23),
    .B(pp_row48_24),
    .CIN(pp_row48_25),
    .COUT(\c$1302 ),
    .SUM(\s$1303 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_48_1 (.A(pp_row48_26),
    .B(\c$302 ),
    .CIN(\c$304 ),
    .COUT(\c$1304 ),
    .SUM(\s$1305 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_48_2 (.A(\c$306 ),
    .B(\c$308 ),
    .CIN(\c$310 ),
    .COUT(\c$1306 ),
    .SUM(\s$1307 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_48_3 (.A(\c$312 ),
    .B(\c$314 ),
    .CIN(\s$317 ),
    .COUT(\c$1308 ),
    .SUM(\s$1309 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_48_4 (.A(\s$319 ),
    .B(\s$321 ),
    .CIN(\s$323 ),
    .COUT(\c$1310 ),
    .SUM(\s$1311 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_48_5 (.A(\s$325 ),
    .B(\s$327 ),
    .CIN(\s$329 ),
    .COUT(\c$1312 ),
    .SUM(\s$1313 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_49_0 (.A(pp_row49_23),
    .B(pp_row49_24),
    .CIN(pp_row49_25),
    .COUT(\c$1314 ),
    .SUM(\s$1315 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_49_1 (.A(\c$316 ),
    .B(\c$318 ),
    .CIN(\c$320 ),
    .COUT(\c$1316 ),
    .SUM(\s$1317 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_49_2 (.A(\c$322 ),
    .B(\c$324 ),
    .CIN(\c$326 ),
    .COUT(\c$1318 ),
    .SUM(\s$1319 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_49_3 (.A(\c$328 ),
    .B(\c$330 ),
    .CIN(\s$333 ),
    .COUT(\c$1320 ),
    .SUM(\s$1321 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_49_4 (.A(\s$335 ),
    .B(\s$337 ),
    .CIN(\s$339 ),
    .COUT(\c$1322 ),
    .SUM(\s$1323 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_49_5 (.A(\s$341 ),
    .B(\s$343 ),
    .CIN(\s$345 ),
    .COUT(\c$1324 ),
    .SUM(\s$1325 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_50_0 (.A(pp_row50_26),
    .B(pp_row50_27),
    .CIN(\c$332 ),
    .COUT(\c$1326 ),
    .SUM(\s$1327 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_50_1 (.A(\c$334 ),
    .B(\c$336 ),
    .CIN(\c$338 ),
    .COUT(\c$1328 ),
    .SUM(\s$1329 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_50_2 (.A(\c$340 ),
    .B(\c$342 ),
    .CIN(\c$344 ),
    .COUT(\c$1330 ),
    .SUM(\s$1331 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_50_3 (.A(\c$346 ),
    .B(\s$349 ),
    .CIN(\s$351 ),
    .COUT(\c$1332 ),
    .SUM(\s$1333 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_50_4 (.A(\s$353 ),
    .B(\s$355 ),
    .CIN(\s$357 ),
    .COUT(\c$1334 ),
    .SUM(\s$1335 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_50_5 (.A(\s$359 ),
    .B(\s$361 ),
    .CIN(\s$363 ),
    .COUT(\c$1336 ),
    .SUM(\s$1337 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_51_0 (.A(pp_row51_26),
    .B(\c$348 ),
    .CIN(\c$350 ),
    .COUT(\c$1338 ),
    .SUM(\s$1339 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_51_1 (.A(\c$352 ),
    .B(\c$354 ),
    .CIN(\c$356 ),
    .COUT(\c$1340 ),
    .SUM(\s$1341 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_51_2 (.A(\c$358 ),
    .B(\c$360 ),
    .CIN(\c$362 ),
    .COUT(\c$1342 ),
    .SUM(\s$1343 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_51_3 (.A(\c$364 ),
    .B(\s$367 ),
    .CIN(\s$369 ),
    .COUT(\c$1344 ),
    .SUM(\s$1345 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_51_4 (.A(\s$371 ),
    .B(\s$373 ),
    .CIN(\s$375 ),
    .COUT(\c$1346 ),
    .SUM(\s$1347 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_51_5 (.A(\s$377 ),
    .B(\s$379 ),
    .CIN(\s$381 ),
    .COUT(\c$1348 ),
    .SUM(\s$1349 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_52_0 (.A(s),
    .B(\c$366 ),
    .CIN(\c$368 ),
    .COUT(\c$1350 ),
    .SUM(\s$1351 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_52_1 (.A(\c$370 ),
    .B(\c$372 ),
    .CIN(\c$374 ),
    .COUT(\c$1352 ),
    .SUM(\s$1353 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_52_2 (.A(\c$376 ),
    .B(\c$378 ),
    .CIN(\c$380 ),
    .COUT(\c$1354 ),
    .SUM(\s$1355 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_52_3 (.A(\c$382 ),
    .B(\s$385 ),
    .CIN(\s$387 ),
    .COUT(\c$1356 ),
    .SUM(\s$1357 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_52_4 (.A(\s$389 ),
    .B(\s$391 ),
    .CIN(\s$393 ),
    .COUT(\c$1358 ),
    .SUM(\s$1359 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_52_5 (.A(\s$395 ),
    .B(\s$397 ),
    .CIN(\s$399 ),
    .COUT(\c$1360 ),
    .SUM(\s$1361 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_53_0 (.A(\s$3 ),
    .B(\c$384 ),
    .CIN(\c$386 ),
    .COUT(\c$1362 ),
    .SUM(\s$1363 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_53_1 (.A(\c$388 ),
    .B(\c$390 ),
    .CIN(\c$392 ),
    .COUT(\c$1364 ),
    .SUM(\s$1365 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_53_2 (.A(\c$394 ),
    .B(\c$396 ),
    .CIN(\c$398 ),
    .COUT(\c$1366 ),
    .SUM(\s$1367 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_53_3 (.A(\c$400 ),
    .B(\s$403 ),
    .CIN(\s$405 ),
    .COUT(\c$1368 ),
    .SUM(\s$1369 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_53_4 (.A(\s$407 ),
    .B(\s$409 ),
    .CIN(\s$411 ),
    .COUT(\c$1370 ),
    .SUM(\s$1371 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_53_5 (.A(\s$413 ),
    .B(\s$415 ),
    .CIN(\s$417 ),
    .COUT(\c$1372 ),
    .SUM(\s$1373 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_54_0 (.A(\s$7 ),
    .B(\c$402 ),
    .CIN(\c$404 ),
    .COUT(\c$1374 ),
    .SUM(\s$1375 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_54_1 (.A(\c$406 ),
    .B(\c$408 ),
    .CIN(\c$410 ),
    .COUT(\c$1376 ),
    .SUM(\s$1377 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_54_2 (.A(\c$412 ),
    .B(\c$414 ),
    .CIN(\c$416 ),
    .COUT(\c$1378 ),
    .SUM(\s$1379 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_54_3 (.A(\c$418 ),
    .B(\s$421 ),
    .CIN(\s$423 ),
    .COUT(\c$1380 ),
    .SUM(\s$1381 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_54_4 (.A(\s$425 ),
    .B(\s$427 ),
    .CIN(\s$429 ),
    .COUT(\c$1382 ),
    .SUM(\s$1383 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_54_5 (.A(\s$431 ),
    .B(\s$433 ),
    .CIN(\s$435 ),
    .COUT(\c$1384 ),
    .SUM(\s$1385 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_55_0 (.A(\s$11 ),
    .B(\c$420 ),
    .CIN(\c$422 ),
    .COUT(\c$1386 ),
    .SUM(\s$1387 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_55_1 (.A(\c$424 ),
    .B(\c$426 ),
    .CIN(\c$428 ),
    .COUT(\c$1388 ),
    .SUM(\s$1389 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_55_2 (.A(\c$430 ),
    .B(\c$432 ),
    .CIN(\c$434 ),
    .COUT(\c$1390 ),
    .SUM(\s$1391 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_55_3 (.A(\c$436 ),
    .B(\s$439 ),
    .CIN(\s$441 ),
    .COUT(\c$1392 ),
    .SUM(\s$1393 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_55_4 (.A(\s$443 ),
    .B(\s$445 ),
    .CIN(\s$447 ),
    .COUT(\c$1394 ),
    .SUM(\s$1395 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_55_5 (.A(\s$449 ),
    .B(\s$451 ),
    .CIN(\s$453 ),
    .COUT(\c$1396 ),
    .SUM(\s$1397 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_56_0 (.A(\s$17 ),
    .B(\c$438 ),
    .CIN(\c$440 ),
    .COUT(\c$1398 ),
    .SUM(\s$1399 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_56_1 (.A(\c$442 ),
    .B(\c$444 ),
    .CIN(\c$446 ),
    .COUT(\c$1400 ),
    .SUM(\s$1401 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_56_2 (.A(\c$448 ),
    .B(\c$450 ),
    .CIN(\c$452 ),
    .COUT(\c$1402 ),
    .SUM(\s$1403 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_56_3 (.A(\c$454 ),
    .B(\s$457 ),
    .CIN(\s$459 ),
    .COUT(\c$1404 ),
    .SUM(\s$1405 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_56_4 (.A(\s$461 ),
    .B(\s$463 ),
    .CIN(\s$465 ),
    .COUT(\c$1406 ),
    .SUM(\s$1407 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_56_5 (.A(\s$467 ),
    .B(\s$469 ),
    .CIN(\s$471 ),
    .COUT(\c$1408 ),
    .SUM(\s$1409 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_57_0 (.A(\s$23 ),
    .B(\c$456 ),
    .CIN(\c$458 ),
    .COUT(\c$1410 ),
    .SUM(\s$1411 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_57_1 (.A(\c$460 ),
    .B(\c$462 ),
    .CIN(\c$464 ),
    .COUT(\c$1412 ),
    .SUM(\s$1413 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_57_2 (.A(\c$466 ),
    .B(\c$468 ),
    .CIN(\c$470 ),
    .COUT(\c$1414 ),
    .SUM(\s$1415 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_57_3 (.A(\c$472 ),
    .B(\s$475 ),
    .CIN(\s$477 ),
    .COUT(\c$1416 ),
    .SUM(\s$1417 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_57_4 (.A(\s$479 ),
    .B(\s$481 ),
    .CIN(\s$483 ),
    .COUT(\c$1418 ),
    .SUM(\s$1419 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_57_5 (.A(\s$485 ),
    .B(\s$487 ),
    .CIN(\s$489 ),
    .COUT(\c$1420 ),
    .SUM(\s$1421 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_58_0 (.A(\s$31 ),
    .B(\c$474 ),
    .CIN(\c$476 ),
    .COUT(\c$1422 ),
    .SUM(\s$1423 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_58_1 (.A(\c$478 ),
    .B(\c$480 ),
    .CIN(\c$482 ),
    .COUT(\c$1424 ),
    .SUM(\s$1425 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_58_2 (.A(\c$484 ),
    .B(\c$486 ),
    .CIN(\c$488 ),
    .COUT(\c$1426 ),
    .SUM(\s$1427 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_58_3 (.A(\c$490 ),
    .B(\s$493 ),
    .CIN(\s$495 ),
    .COUT(\c$1428 ),
    .SUM(\s$1429 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_58_4 (.A(\s$497 ),
    .B(\s$499 ),
    .CIN(\s$501 ),
    .COUT(\c$1430 ),
    .SUM(\s$1431 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_58_5 (.A(\s$503 ),
    .B(\s$505 ),
    .CIN(\s$507 ),
    .COUT(\c$1432 ),
    .SUM(\s$1433 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_59_0 (.A(\s$39 ),
    .B(\c$492 ),
    .CIN(\c$494 ),
    .COUT(\c$1434 ),
    .SUM(\s$1435 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_59_1 (.A(\c$496 ),
    .B(\c$498 ),
    .CIN(\c$500 ),
    .COUT(\c$1436 ),
    .SUM(\s$1437 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_59_2 (.A(\c$502 ),
    .B(\c$504 ),
    .CIN(\c$506 ),
    .COUT(\c$1438 ),
    .SUM(\s$1439 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_59_3 (.A(\c$508 ),
    .B(\s$511 ),
    .CIN(\s$513 ),
    .COUT(\c$1440 ),
    .SUM(\s$1441 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_59_4 (.A(\s$515 ),
    .B(\s$517 ),
    .CIN(\s$519 ),
    .COUT(\c$1442 ),
    .SUM(\s$1443 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_59_5 (.A(\s$521 ),
    .B(\s$523 ),
    .CIN(\s$525 ),
    .COUT(\c$1444 ),
    .SUM(\s$1445 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_60_0 (.A(\s$49 ),
    .B(\c$510 ),
    .CIN(\c$512 ),
    .COUT(\c$1446 ),
    .SUM(\s$1447 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_60_1 (.A(\c$514 ),
    .B(\c$516 ),
    .CIN(\c$518 ),
    .COUT(\c$1448 ),
    .SUM(\s$1449 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_60_2 (.A(\c$520 ),
    .B(\c$522 ),
    .CIN(\c$524 ),
    .COUT(\c$1450 ),
    .SUM(\s$1451 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_60_3 (.A(\c$526 ),
    .B(\s$529 ),
    .CIN(\s$531 ),
    .COUT(\c$1452 ),
    .SUM(\s$1453 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_60_4 (.A(\s$533 ),
    .B(\s$535 ),
    .CIN(\s$537 ),
    .COUT(\c$1454 ),
    .SUM(\s$1455 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_60_5 (.A(\s$539 ),
    .B(\s$541 ),
    .CIN(\s$543 ),
    .COUT(\c$1456 ),
    .SUM(\s$1457 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_61_0 (.A(\s$59 ),
    .B(\c$528 ),
    .CIN(\c$530 ),
    .COUT(\c$1458 ),
    .SUM(\s$1459 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_61_1 (.A(\c$532 ),
    .B(\c$534 ),
    .CIN(\c$536 ),
    .COUT(\c$1460 ),
    .SUM(\s$1461 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_61_2 (.A(\c$538 ),
    .B(\c$540 ),
    .CIN(\c$542 ),
    .COUT(\c$1462 ),
    .SUM(\s$1463 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_61_3 (.A(\c$544 ),
    .B(\s$547 ),
    .CIN(\s$549 ),
    .COUT(\c$1464 ),
    .SUM(\s$1465 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_61_4 (.A(\s$551 ),
    .B(\s$553 ),
    .CIN(\s$555 ),
    .COUT(\c$1466 ),
    .SUM(\s$1467 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_61_5 (.A(\s$557 ),
    .B(\s$559 ),
    .CIN(\s$561 ),
    .COUT(\c$1468 ),
    .SUM(\s$1469 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_62_0 (.A(\s$71 ),
    .B(\c$546 ),
    .CIN(\c$548 ),
    .COUT(\c$1470 ),
    .SUM(\s$1471 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_62_1 (.A(\c$550 ),
    .B(\c$552 ),
    .CIN(\c$554 ),
    .COUT(\c$1472 ),
    .SUM(\s$1473 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_62_2 (.A(\c$556 ),
    .B(\c$558 ),
    .CIN(\c$560 ),
    .COUT(\c$1474 ),
    .SUM(\s$1475 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_62_3 (.A(\c$562 ),
    .B(\s$565 ),
    .CIN(\s$567 ),
    .COUT(\c$1476 ),
    .SUM(\s$1477 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_62_4 (.A(\s$569 ),
    .B(\s$571 ),
    .CIN(\s$573 ),
    .COUT(\c$1478 ),
    .SUM(\s$1479 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_62_5 (.A(\s$575 ),
    .B(\s$577 ),
    .CIN(\s$579 ),
    .COUT(\c$1480 ),
    .SUM(\s$1481 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_63_0 (.A(\s$83 ),
    .B(\c$564 ),
    .CIN(\c$566 ),
    .COUT(\c$1482 ),
    .SUM(\s$1483 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_63_1 (.A(\c$568 ),
    .B(\c$570 ),
    .CIN(\c$572 ),
    .COUT(\c$1484 ),
    .SUM(\s$1485 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_63_2 (.A(\c$574 ),
    .B(\c$576 ),
    .CIN(\c$578 ),
    .COUT(\c$1486 ),
    .SUM(\s$1487 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_63_3 (.A(\c$580 ),
    .B(\s$583 ),
    .CIN(\s$585 ),
    .COUT(\c$1488 ),
    .SUM(\s$1489 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_63_4 (.A(\s$587 ),
    .B(\s$589 ),
    .CIN(\s$591 ),
    .COUT(\c$1490 ),
    .SUM(\s$1491 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_63_5 (.A(\s$593 ),
    .B(\s$595 ),
    .CIN(\s$597 ),
    .COUT(\c$1492 ),
    .SUM(\s$1493 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_64_0 (.A(\s$95 ),
    .B(\c$582 ),
    .CIN(\c$584 ),
    .COUT(\c$1494 ),
    .SUM(\s$1495 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_64_1 (.A(\c$586 ),
    .B(\c$588 ),
    .CIN(\c$590 ),
    .COUT(\c$1496 ),
    .SUM(\s$1497 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_64_2 (.A(\c$592 ),
    .B(\c$594 ),
    .CIN(\c$596 ),
    .COUT(\c$1498 ),
    .SUM(\s$1499 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_64_3 (.A(\c$598 ),
    .B(\s$601 ),
    .CIN(\s$603 ),
    .COUT(\c$1500 ),
    .SUM(\s$1501 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_64_4 (.A(\s$605 ),
    .B(\s$607 ),
    .CIN(\s$609 ),
    .COUT(\c$1502 ),
    .SUM(\s$1503 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_64_5 (.A(\s$611 ),
    .B(\s$613 ),
    .CIN(\s$615 ),
    .COUT(\c$1504 ),
    .SUM(\s$1505 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_65_0 (.A(\s$107 ),
    .B(\c$600 ),
    .CIN(\c$602 ),
    .COUT(\c$1506 ),
    .SUM(\s$1507 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_65_1 (.A(\c$604 ),
    .B(\c$606 ),
    .CIN(\c$608 ),
    .COUT(\c$1508 ),
    .SUM(\s$1509 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_65_2 (.A(\c$610 ),
    .B(\c$612 ),
    .CIN(\c$614 ),
    .COUT(\c$1510 ),
    .SUM(\s$1511 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_65_3 (.A(\c$616 ),
    .B(\s$619 ),
    .CIN(\s$621 ),
    .COUT(\c$1512 ),
    .SUM(\s$1513 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_65_4 (.A(\s$623 ),
    .B(\s$625 ),
    .CIN(\s$627 ),
    .COUT(\c$1514 ),
    .SUM(\s$1515 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_65_5 (.A(\s$629 ),
    .B(\s$631 ),
    .CIN(\s$633 ),
    .COUT(\c$1516 ),
    .SUM(\s$1517 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_66_0 (.A(\s$119 ),
    .B(\c$618 ),
    .CIN(\c$620 ),
    .COUT(\c$1518 ),
    .SUM(\s$1519 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_66_1 (.A(\c$622 ),
    .B(\c$624 ),
    .CIN(\c$626 ),
    .COUT(\c$1520 ),
    .SUM(\s$1521 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_66_2 (.A(\c$628 ),
    .B(\c$630 ),
    .CIN(\c$632 ),
    .COUT(\c$1522 ),
    .SUM(\s$1523 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_66_3 (.A(\c$634 ),
    .B(\s$637 ),
    .CIN(\s$639 ),
    .COUT(\c$1524 ),
    .SUM(\s$1525 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_66_4 (.A(\s$641 ),
    .B(\s$643 ),
    .CIN(\s$645 ),
    .COUT(\c$1526 ),
    .SUM(\s$1527 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_66_5 (.A(\s$647 ),
    .B(\s$649 ),
    .CIN(\s$651 ),
    .COUT(\c$1528 ),
    .SUM(\s$1529 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_67_0 (.A(\s$131 ),
    .B(\c$636 ),
    .CIN(\c$638 ),
    .COUT(\c$1530 ),
    .SUM(\s$1531 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_67_1 (.A(\c$640 ),
    .B(\c$642 ),
    .CIN(\c$644 ),
    .COUT(\c$1532 ),
    .SUM(\s$1533 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_67_2 (.A(\c$646 ),
    .B(\c$648 ),
    .CIN(\c$650 ),
    .COUT(\c$1534 ),
    .SUM(\s$1535 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_67_3 (.A(\c$652 ),
    .B(\s$655 ),
    .CIN(\s$657 ),
    .COUT(\c$1536 ),
    .SUM(\s$1537 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_67_4 (.A(\s$659 ),
    .B(\s$661 ),
    .CIN(\s$663 ),
    .COUT(\c$1538 ),
    .SUM(\s$1539 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_67_5 (.A(\s$665 ),
    .B(\s$667 ),
    .CIN(\s$669 ),
    .COUT(\c$1540 ),
    .SUM(\s$1541 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_68_0 (.A(\s$143 ),
    .B(\c$654 ),
    .CIN(\c$656 ),
    .COUT(\c$1542 ),
    .SUM(\s$1543 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_68_1 (.A(\c$658 ),
    .B(\c$660 ),
    .CIN(\c$662 ),
    .COUT(\c$1544 ),
    .SUM(\s$1545 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_68_2 (.A(\c$664 ),
    .B(\c$666 ),
    .CIN(\c$668 ),
    .COUT(\c$1546 ),
    .SUM(\s$1547 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_68_3 (.A(\c$670 ),
    .B(\s$673 ),
    .CIN(\s$675 ),
    .COUT(\c$1548 ),
    .SUM(\s$1549 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_68_4 (.A(\s$677 ),
    .B(\s$679 ),
    .CIN(\s$681 ),
    .COUT(\c$1550 ),
    .SUM(\s$1551 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_68_5 (.A(\s$683 ),
    .B(\s$685 ),
    .CIN(\s$687 ),
    .COUT(\c$1552 ),
    .SUM(\s$1553 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_69_0 (.A(\s$153 ),
    .B(\c$672 ),
    .CIN(\c$674 ),
    .COUT(\c$1554 ),
    .SUM(\s$1555 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_69_1 (.A(\c$676 ),
    .B(\c$678 ),
    .CIN(\c$680 ),
    .COUT(\c$1556 ),
    .SUM(\s$1557 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_69_2 (.A(\c$682 ),
    .B(\c$684 ),
    .CIN(\c$686 ),
    .COUT(\c$1558 ),
    .SUM(\s$1559 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_69_3 (.A(\c$688 ),
    .B(\s$691 ),
    .CIN(\s$693 ),
    .COUT(\c$1560 ),
    .SUM(\s$1561 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_69_4 (.A(\s$695 ),
    .B(\s$697 ),
    .CIN(\s$699 ),
    .COUT(\c$1562 ),
    .SUM(\s$1563 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_69_5 (.A(\s$701 ),
    .B(\s$703 ),
    .CIN(\s$705 ),
    .COUT(\c$1564 ),
    .SUM(\s$1565 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_70_0 (.A(\s$163 ),
    .B(\c$690 ),
    .CIN(\c$692 ),
    .COUT(\c$1566 ),
    .SUM(\s$1567 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_70_1 (.A(\c$694 ),
    .B(\c$696 ),
    .CIN(\c$698 ),
    .COUT(\c$1568 ),
    .SUM(\s$1569 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_70_2 (.A(\c$700 ),
    .B(\c$702 ),
    .CIN(\c$704 ),
    .COUT(\c$1570 ),
    .SUM(\s$1571 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_70_3 (.A(\c$706 ),
    .B(\s$709 ),
    .CIN(\s$711 ),
    .COUT(\c$1572 ),
    .SUM(\s$1573 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_70_4 (.A(\s$713 ),
    .B(\s$715 ),
    .CIN(\s$717 ),
    .COUT(\c$1574 ),
    .SUM(\s$1575 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_70_5 (.A(\s$719 ),
    .B(\s$721 ),
    .CIN(\s$723 ),
    .COUT(\c$1576 ),
    .SUM(\s$1577 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_71_0 (.A(\s$171 ),
    .B(\c$708 ),
    .CIN(\c$710 ),
    .COUT(\c$1578 ),
    .SUM(\s$1579 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_71_1 (.A(\c$712 ),
    .B(\c$714 ),
    .CIN(\c$716 ),
    .COUT(\c$1580 ),
    .SUM(\s$1581 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_71_2 (.A(\c$718 ),
    .B(\c$720 ),
    .CIN(\c$722 ),
    .COUT(\c$1582 ),
    .SUM(\s$1583 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_71_3 (.A(\c$724 ),
    .B(\s$727 ),
    .CIN(\s$729 ),
    .COUT(\c$1584 ),
    .SUM(\s$1585 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_71_4 (.A(\s$731 ),
    .B(\s$733 ),
    .CIN(\s$735 ),
    .COUT(\c$1586 ),
    .SUM(\s$1587 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_71_5 (.A(\s$737 ),
    .B(\s$739 ),
    .CIN(\s$741 ),
    .COUT(\c$1588 ),
    .SUM(\s$1589 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_72_0 (.A(\s$179 ),
    .B(\c$726 ),
    .CIN(\c$728 ),
    .COUT(\c$1590 ),
    .SUM(\s$1591 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_72_1 (.A(\c$730 ),
    .B(\c$732 ),
    .CIN(\c$734 ),
    .COUT(\c$1592 ),
    .SUM(\s$1593 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_72_2 (.A(\c$736 ),
    .B(\c$738 ),
    .CIN(\c$740 ),
    .COUT(\c$1594 ),
    .SUM(\s$1595 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_72_3 (.A(\c$742 ),
    .B(\s$745 ),
    .CIN(\s$747 ),
    .COUT(\c$1596 ),
    .SUM(\s$1597 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_72_4 (.A(\s$749 ),
    .B(\s$751 ),
    .CIN(\s$753 ),
    .COUT(\c$1598 ),
    .SUM(\s$1599 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_72_5 (.A(\s$755 ),
    .B(\s$757 ),
    .CIN(\s$759 ),
    .COUT(\c$1600 ),
    .SUM(\s$1601 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_73_0 (.A(\s$185 ),
    .B(\c$744 ),
    .CIN(\c$746 ),
    .COUT(\c$1602 ),
    .SUM(\s$1603 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_73_1 (.A(\c$748 ),
    .B(\c$750 ),
    .CIN(\c$752 ),
    .COUT(\c$1604 ),
    .SUM(\s$1605 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_73_2 (.A(\c$754 ),
    .B(\c$756 ),
    .CIN(\c$758 ),
    .COUT(\c$1606 ),
    .SUM(\s$1607 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_73_3 (.A(\c$760 ),
    .B(\s$763 ),
    .CIN(\s$765 ),
    .COUT(\c$1608 ),
    .SUM(\s$1609 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_73_4 (.A(\s$767 ),
    .B(\s$769 ),
    .CIN(\s$771 ),
    .COUT(\c$1610 ),
    .SUM(\s$1611 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_73_5 (.A(\s$773 ),
    .B(\s$775 ),
    .CIN(\s$777 ),
    .COUT(\c$1612 ),
    .SUM(\s$1613 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_74_0 (.A(\s$191 ),
    .B(\c$762 ),
    .CIN(\c$764 ),
    .COUT(\c$1614 ),
    .SUM(\s$1615 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_74_1 (.A(\c$766 ),
    .B(\c$768 ),
    .CIN(\c$770 ),
    .COUT(\c$1616 ),
    .SUM(\s$1617 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_74_2 (.A(\c$772 ),
    .B(\c$774 ),
    .CIN(\c$776 ),
    .COUT(\c$1618 ),
    .SUM(\s$1619 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_74_3 (.A(\c$778 ),
    .B(\s$781 ),
    .CIN(\s$783 ),
    .COUT(\c$1620 ),
    .SUM(\s$1621 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_74_4 (.A(\s$785 ),
    .B(\s$787 ),
    .CIN(\s$789 ),
    .COUT(\c$1622 ),
    .SUM(\s$1623 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_74_5 (.A(\s$791 ),
    .B(\s$793 ),
    .CIN(\s$795 ),
    .COUT(\c$1624 ),
    .SUM(\s$1625 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_75_0 (.A(\s$195 ),
    .B(\c$780 ),
    .CIN(\c$782 ),
    .COUT(\c$1626 ),
    .SUM(\s$1627 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_75_1 (.A(\c$784 ),
    .B(\c$786 ),
    .CIN(\c$788 ),
    .COUT(\c$1628 ),
    .SUM(\s$1629 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_75_2 (.A(\c$790 ),
    .B(\c$792 ),
    .CIN(\c$794 ),
    .COUT(\c$1630 ),
    .SUM(\s$1631 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_75_3 (.A(\c$796 ),
    .B(\s$799 ),
    .CIN(\s$801 ),
    .COUT(\c$1632 ),
    .SUM(\s$1633 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_75_4 (.A(\s$803 ),
    .B(\s$805 ),
    .CIN(\s$807 ),
    .COUT(\c$1634 ),
    .SUM(\s$1635 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_75_5 (.A(\s$809 ),
    .B(\s$811 ),
    .CIN(\s$813 ),
    .COUT(\c$1636 ),
    .SUM(\s$1637 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_76_0 (.A(\s$199 ),
    .B(\c$798 ),
    .CIN(\c$800 ),
    .COUT(\c$1638 ),
    .SUM(\s$1639 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_76_1 (.A(\c$802 ),
    .B(\c$804 ),
    .CIN(\c$806 ),
    .COUT(\c$1640 ),
    .SUM(\s$1641 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_76_2 (.A(\c$808 ),
    .B(\c$810 ),
    .CIN(\c$812 ),
    .COUT(\c$1642 ),
    .SUM(\s$1643 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_76_3 (.A(\c$814 ),
    .B(\s$817 ),
    .CIN(\s$819 ),
    .COUT(\c$1644 ),
    .SUM(\s$1645 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_76_4 (.A(\s$821 ),
    .B(\s$823 ),
    .CIN(\s$825 ),
    .COUT(\c$1646 ),
    .SUM(\s$1647 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_76_5 (.A(\s$827 ),
    .B(\s$829 ),
    .CIN(\s$831 ),
    .COUT(\c$1648 ),
    .SUM(\s$1649 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_77_0 (.A(\s$201 ),
    .B(\c$816 ),
    .CIN(\c$818 ),
    .COUT(\c$1650 ),
    .SUM(\s$1651 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_77_1 (.A(\c$820 ),
    .B(\c$822 ),
    .CIN(\c$824 ),
    .COUT(\c$1652 ),
    .SUM(\s$1653 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_77_2 (.A(\c$826 ),
    .B(\c$828 ),
    .CIN(\c$830 ),
    .COUT(\c$1654 ),
    .SUM(\s$1655 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_77_3 (.A(\c$832 ),
    .B(\s$835 ),
    .CIN(\s$837 ),
    .COUT(\c$1656 ),
    .SUM(\s$1657 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_77_4 (.A(\s$839 ),
    .B(\s$841 ),
    .CIN(\s$843 ),
    .COUT(\c$1658 ),
    .SUM(\s$1659 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_77_5 (.A(\s$845 ),
    .B(\s$847 ),
    .CIN(\s$849 ),
    .COUT(\c$1660 ),
    .SUM(\s$1661 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_78_0 (.A(\s$203 ),
    .B(\c$834 ),
    .CIN(\c$836 ),
    .COUT(\c$1662 ),
    .SUM(\s$1663 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_78_1 (.A(\c$838 ),
    .B(\c$840 ),
    .CIN(\c$842 ),
    .COUT(\c$1664 ),
    .SUM(\s$1665 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_78_2 (.A(\c$844 ),
    .B(\c$846 ),
    .CIN(\c$848 ),
    .COUT(\c$1666 ),
    .SUM(\s$1667 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_78_3 (.A(\c$850 ),
    .B(\s$853 ),
    .CIN(\s$855 ),
    .COUT(\c$1668 ),
    .SUM(\s$1669 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_78_4 (.A(\s$857 ),
    .B(\s$859 ),
    .CIN(\s$861 ),
    .COUT(\c$1670 ),
    .SUM(\s$1671 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_78_5 (.A(\s$863 ),
    .B(\s$865 ),
    .CIN(\s$867 ),
    .COUT(\c$1672 ),
    .SUM(\s$1673 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_79_0 (.A(\c$202 ),
    .B(\c$852 ),
    .CIN(\c$854 ),
    .COUT(\c$1674 ),
    .SUM(\s$1675 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_79_1 (.A(\c$856 ),
    .B(\c$858 ),
    .CIN(\c$860 ),
    .COUT(\c$1676 ),
    .SUM(\s$1677 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_79_2 (.A(\c$862 ),
    .B(\c$864 ),
    .CIN(\c$866 ),
    .COUT(\c$1678 ),
    .SUM(\s$1679 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_79_3 (.A(\c$868 ),
    .B(\s$871 ),
    .CIN(\s$873 ),
    .COUT(\c$1680 ),
    .SUM(\s$1681 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_79_4 (.A(\s$875 ),
    .B(\s$877 ),
    .CIN(\s$879 ),
    .COUT(\c$1682 ),
    .SUM(\s$1683 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_79_5 (.A(\s$881 ),
    .B(\s$883 ),
    .CIN(\s$885 ),
    .COUT(\c$1684 ),
    .SUM(\s$1685 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_80_0 (.A(pp_row80_26),
    .B(\c$870 ),
    .CIN(\c$872 ),
    .COUT(\c$1686 ),
    .SUM(\s$1687 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_80_1 (.A(\c$874 ),
    .B(\c$876 ),
    .CIN(\c$878 ),
    .COUT(\c$1688 ),
    .SUM(\s$1689 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_80_2 (.A(\c$880 ),
    .B(\c$882 ),
    .CIN(\c$884 ),
    .COUT(\c$1690 ),
    .SUM(\s$1691 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_80_3 (.A(\c$886 ),
    .B(\s$889 ),
    .CIN(\s$891 ),
    .COUT(\c$1692 ),
    .SUM(\s$1693 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_80_4 (.A(\s$893 ),
    .B(\s$895 ),
    .CIN(\s$897 ),
    .COUT(\c$1694 ),
    .SUM(\s$1695 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_80_5 (.A(\s$899 ),
    .B(\s$901 ),
    .CIN(\s$903 ),
    .COUT(\c$1696 ),
    .SUM(\s$1697 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_81_0 (.A(pp_row81_24),
    .B(pp_row81_25),
    .CIN(\c$888 ),
    .COUT(\c$1698 ),
    .SUM(\s$1699 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_81_1 (.A(\c$890 ),
    .B(\c$892 ),
    .CIN(\c$894 ),
    .COUT(\c$1700 ),
    .SUM(\s$1701 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_81_2 (.A(\c$896 ),
    .B(\c$898 ),
    .CIN(\c$900 ),
    .COUT(\c$1702 ),
    .SUM(\s$1703 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_81_3 (.A(\c$902 ),
    .B(\c$904 ),
    .CIN(\s$907 ),
    .COUT(\c$1704 ),
    .SUM(\s$1705 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_81_4 (.A(\s$909 ),
    .B(\s$911 ),
    .CIN(\s$913 ),
    .COUT(\c$1706 ),
    .SUM(\s$1707 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_81_5 (.A(\s$915 ),
    .B(\s$917 ),
    .CIN(\s$919 ),
    .COUT(\c$1708 ),
    .SUM(\s$1709 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_82_0 (.A(pp_row82_23),
    .B(pp_row82_24),
    .CIN(pp_row82_25),
    .COUT(\c$1710 ),
    .SUM(\s$1711 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_82_1 (.A(\c$906 ),
    .B(\c$908 ),
    .CIN(\c$910 ),
    .COUT(\c$1712 ),
    .SUM(\s$1713 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_82_2 (.A(\c$912 ),
    .B(\c$914 ),
    .CIN(\c$916 ),
    .COUT(\c$1714 ),
    .SUM(\s$1715 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_82_3 (.A(\c$918 ),
    .B(\c$920 ),
    .CIN(\s$923 ),
    .COUT(\c$1716 ),
    .SUM(\s$1717 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_82_4 (.A(\s$925 ),
    .B(\s$927 ),
    .CIN(\s$929 ),
    .COUT(\c$1718 ),
    .SUM(\s$1719 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_82_5 (.A(\s$931 ),
    .B(\s$933 ),
    .CIN(\s$935 ),
    .COUT(\c$1720 ),
    .SUM(\s$1721 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_83_0 (.A(pp_row83_21),
    .B(pp_row83_22),
    .CIN(pp_row83_23),
    .COUT(\c$1722 ),
    .SUM(\s$1723 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_83_1 (.A(pp_row83_24),
    .B(\c$922 ),
    .CIN(\c$924 ),
    .COUT(\c$1724 ),
    .SUM(\s$1725 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_83_2 (.A(\c$926 ),
    .B(\c$928 ),
    .CIN(\c$930 ),
    .COUT(\c$1726 ),
    .SUM(\s$1727 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_83_3 (.A(\c$932 ),
    .B(\c$934 ),
    .CIN(\c$936 ),
    .COUT(\c$1728 ),
    .SUM(\s$1729 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_83_4 (.A(\s$939 ),
    .B(\s$941 ),
    .CIN(\s$943 ),
    .COUT(\c$1730 ),
    .SUM(\s$1731 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_83_5 (.A(\s$945 ),
    .B(\s$947 ),
    .CIN(\s$949 ),
    .COUT(\c$1732 ),
    .SUM(\s$1733 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_84_0 (.A(pp_row84_20),
    .B(pp_row84_21),
    .CIN(pp_row84_22),
    .COUT(\c$1734 ),
    .SUM(\s$1735 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_84_1 (.A(pp_row84_23),
    .B(pp_row84_24),
    .CIN(\c$938 ),
    .COUT(\c$1736 ),
    .SUM(\s$1737 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_84_2 (.A(\c$940 ),
    .B(\c$942 ),
    .CIN(\c$944 ),
    .COUT(\c$1738 ),
    .SUM(\s$1739 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_84_3 (.A(\c$946 ),
    .B(\c$948 ),
    .CIN(\c$950 ),
    .COUT(\c$1740 ),
    .SUM(\s$1741 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_84_4 (.A(\s$953 ),
    .B(\s$955 ),
    .CIN(\s$957 ),
    .COUT(\c$1742 ),
    .SUM(\s$1743 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_84_5 (.A(\s$959 ),
    .B(\s$961 ),
    .CIN(\s$963 ),
    .COUT(\c$1744 ),
    .SUM(\s$1745 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_85_0 (.A(pp_row85_18),
    .B(pp_row85_19),
    .CIN(pp_row85_20),
    .COUT(\c$1746 ),
    .SUM(\s$1747 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_85_1 (.A(pp_row85_21),
    .B(pp_row85_22),
    .CIN(pp_row85_23),
    .COUT(\c$1748 ),
    .SUM(\s$1749 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_85_2 (.A(\c$952 ),
    .B(\c$954 ),
    .CIN(\c$956 ),
    .COUT(\c$1750 ),
    .SUM(\s$1751 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_85_3 (.A(\c$958 ),
    .B(\c$960 ),
    .CIN(\c$962 ),
    .COUT(\c$1752 ),
    .SUM(\s$1753 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_85_4 (.A(\c$964 ),
    .B(\s$967 ),
    .CIN(\s$969 ),
    .COUT(\c$1754 ),
    .SUM(\s$1755 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_85_5 (.A(\s$971 ),
    .B(\s$973 ),
    .CIN(\s$975 ),
    .COUT(\c$1756 ),
    .SUM(\s$1757 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_86_0 (.A(pp_row86_17),
    .B(pp_row86_18),
    .CIN(pp_row86_19),
    .COUT(\c$1758 ),
    .SUM(\s$1759 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_86_1 (.A(pp_row86_20),
    .B(pp_row86_21),
    .CIN(pp_row86_22),
    .COUT(\c$1760 ),
    .SUM(\s$1761 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_86_2 (.A(pp_row86_23),
    .B(\c$966 ),
    .CIN(\c$968 ),
    .COUT(\c$1762 ),
    .SUM(\s$1763 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_86_3 (.A(\c$970 ),
    .B(\c$972 ),
    .CIN(\c$974 ),
    .COUT(\c$1764 ),
    .SUM(\s$1765 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_86_4 (.A(\c$976 ),
    .B(\s$979 ),
    .CIN(\s$981 ),
    .COUT(\c$1766 ),
    .SUM(\s$1767 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_86_5 (.A(\s$983 ),
    .B(\s$985 ),
    .CIN(\s$987 ),
    .COUT(\c$1768 ),
    .SUM(\s$1769 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_87_0 (.A(pp_row87_15),
    .B(pp_row87_16),
    .CIN(pp_row87_17),
    .COUT(\c$1770 ),
    .SUM(\s$1771 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_87_1 (.A(pp_row87_18),
    .B(pp_row87_19),
    .CIN(pp_row87_20),
    .COUT(\c$1772 ),
    .SUM(\s$1773 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_87_2 (.A(pp_row87_21),
    .B(pp_row87_22),
    .CIN(\c$978 ),
    .COUT(\c$1774 ),
    .SUM(\s$1775 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_87_3 (.A(\c$980 ),
    .B(\c$982 ),
    .CIN(\c$984 ),
    .COUT(\c$1776 ),
    .SUM(\s$1777 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_87_4 (.A(\c$986 ),
    .B(\c$988 ),
    .CIN(\s$991 ),
    .COUT(\c$1778 ),
    .SUM(\s$1779 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_87_5 (.A(\s$993 ),
    .B(\s$995 ),
    .CIN(\s$997 ),
    .COUT(\c$1780 ),
    .SUM(\s$1781 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_88_0 (.A(pp_row88_14),
    .B(pp_row88_15),
    .CIN(pp_row88_16),
    .COUT(\c$1782 ),
    .SUM(\s$1783 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_88_1 (.A(pp_row88_17),
    .B(pp_row88_18),
    .CIN(pp_row88_19),
    .COUT(\c$1784 ),
    .SUM(\s$1785 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_88_2 (.A(pp_row88_20),
    .B(pp_row88_21),
    .CIN(pp_row88_22),
    .COUT(\c$1786 ),
    .SUM(\s$1787 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_88_3 (.A(\c$990 ),
    .B(\c$992 ),
    .CIN(\c$994 ),
    .COUT(\c$1788 ),
    .SUM(\s$1789 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_88_4 (.A(\c$996 ),
    .B(\c$998 ),
    .CIN(\s$1001 ),
    .COUT(\c$1790 ),
    .SUM(\s$1791 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_88_5 (.A(\s$1003 ),
    .B(\s$1005 ),
    .CIN(\s$1007 ),
    .COUT(\c$1792 ),
    .SUM(\s$1793 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_89_0 (.A(pp_row89_12),
    .B(pp_row89_13),
    .CIN(pp_row89_14),
    .COUT(\c$1794 ),
    .SUM(\s$1795 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_89_1 (.A(pp_row89_15),
    .B(pp_row89_16),
    .CIN(pp_row89_17),
    .COUT(\c$1796 ),
    .SUM(\s$1797 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_89_2 (.A(pp_row89_18),
    .B(pp_row89_19),
    .CIN(pp_row89_20),
    .COUT(\c$1798 ),
    .SUM(\s$1799 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_89_3 (.A(pp_row89_21),
    .B(\c$1000 ),
    .CIN(\c$1002 ),
    .COUT(\c$1800 ),
    .SUM(\s$1801 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_89_4 (.A(\c$1004 ),
    .B(\c$1006 ),
    .CIN(\c$1008 ),
    .COUT(\c$1802 ),
    .SUM(\s$1803 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_89_5 (.A(\s$1011 ),
    .B(\s$1013 ),
    .CIN(\s$1015 ),
    .COUT(\c$1804 ),
    .SUM(\s$1805 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_90_0 (.A(pp_row90_11),
    .B(pp_row90_12),
    .CIN(pp_row90_13),
    .COUT(\c$1806 ),
    .SUM(\s$1807 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_90_1 (.A(pp_row90_14),
    .B(pp_row90_15),
    .CIN(pp_row90_16),
    .COUT(\c$1808 ),
    .SUM(\s$1809 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_90_2 (.A(pp_row90_17),
    .B(pp_row90_18),
    .CIN(pp_row90_19),
    .COUT(\c$1810 ),
    .SUM(\s$1811 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_90_3 (.A(pp_row90_20),
    .B(pp_row90_21),
    .CIN(\c$1010 ),
    .COUT(\c$1812 ),
    .SUM(\s$1813 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_90_4 (.A(\c$1012 ),
    .B(\c$1014 ),
    .CIN(\c$1016 ),
    .COUT(\c$1814 ),
    .SUM(\s$1815 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_90_5 (.A(\s$1019 ),
    .B(\s$1021 ),
    .CIN(\s$1023 ),
    .COUT(\c$1816 ),
    .SUM(\s$1817 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_91_0 (.A(pp_row91_9),
    .B(pp_row91_10),
    .CIN(pp_row91_11),
    .COUT(\c$1818 ),
    .SUM(\s$1819 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_91_1 (.A(pp_row91_12),
    .B(pp_row91_13),
    .CIN(pp_row91_14),
    .COUT(\c$1820 ),
    .SUM(\s$1821 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_91_2 (.A(pp_row91_15),
    .B(pp_row91_16),
    .CIN(pp_row91_17),
    .COUT(\c$1822 ),
    .SUM(\s$1823 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_91_3 (.A(pp_row91_18),
    .B(pp_row91_19),
    .CIN(pp_row91_20),
    .COUT(\c$1824 ),
    .SUM(\s$1825 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_91_4 (.A(\c$1018 ),
    .B(\c$1020 ),
    .CIN(\c$1022 ),
    .COUT(\c$1826 ),
    .SUM(\s$1827 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_91_5 (.A(\c$1024 ),
    .B(\s$1027 ),
    .CIN(\s$1029 ),
    .COUT(\c$1828 ),
    .SUM(\s$1829 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_92_0 (.A(pp_row92_8),
    .B(pp_row92_9),
    .CIN(pp_row92_10),
    .COUT(\c$1830 ),
    .SUM(\s$1831 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_92_1 (.A(pp_row92_11),
    .B(pp_row92_12),
    .CIN(pp_row92_13),
    .COUT(\c$1832 ),
    .SUM(\s$1833 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_92_2 (.A(pp_row92_14),
    .B(pp_row92_15),
    .CIN(pp_row92_16),
    .COUT(\c$1834 ),
    .SUM(\s$1835 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_92_3 (.A(pp_row92_17),
    .B(pp_row92_18),
    .CIN(pp_row92_19),
    .COUT(\c$1836 ),
    .SUM(\s$1837 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_92_4 (.A(pp_row92_20),
    .B(\c$1026 ),
    .CIN(\c$1028 ),
    .COUT(\c$1838 ),
    .SUM(\s$1839 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_92_5 (.A(\c$1030 ),
    .B(\s$1033 ),
    .CIN(\s$1035 ),
    .COUT(\c$1840 ),
    .SUM(\s$1841 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_93_0 (.A(pp_row93_6),
    .B(pp_row93_7),
    .CIN(pp_row93_8),
    .COUT(\c$1842 ),
    .SUM(\s$1843 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_93_1 (.A(pp_row93_9),
    .B(pp_row93_10),
    .CIN(pp_row93_11),
    .COUT(\c$1844 ),
    .SUM(\s$1845 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_93_2 (.A(pp_row93_12),
    .B(pp_row93_13),
    .CIN(pp_row93_14),
    .COUT(\c$1846 ),
    .SUM(\s$1847 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_93_3 (.A(pp_row93_15),
    .B(pp_row93_16),
    .CIN(pp_row93_17),
    .COUT(\c$1848 ),
    .SUM(\s$1849 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_93_4 (.A(pp_row93_18),
    .B(pp_row93_19),
    .CIN(\c$1032 ),
    .COUT(\c$1850 ),
    .SUM(\s$1851 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_93_5 (.A(\c$1034 ),
    .B(\c$1036 ),
    .CIN(\s$1039 ),
    .COUT(\c$1852 ),
    .SUM(\s$1853 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_94_0 (.A(pp_row94_5),
    .B(pp_row94_6),
    .CIN(pp_row94_7),
    .COUT(\c$1854 ),
    .SUM(\s$1855 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_94_1 (.A(pp_row94_8),
    .B(pp_row94_9),
    .CIN(pp_row94_10),
    .COUT(\c$1856 ),
    .SUM(\s$1857 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_94_2 (.A(pp_row94_11),
    .B(pp_row94_12),
    .CIN(pp_row94_13),
    .COUT(\c$1858 ),
    .SUM(\s$1859 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_94_3 (.A(pp_row94_14),
    .B(pp_row94_15),
    .CIN(pp_row94_16),
    .COUT(\c$1860 ),
    .SUM(\s$1861 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_94_4 (.A(pp_row94_17),
    .B(pp_row94_18),
    .CIN(pp_row94_19),
    .COUT(\c$1862 ),
    .SUM(\s$1863 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_94_5 (.A(\c$1038 ),
    .B(\c$1040 ),
    .CIN(\s$1043 ),
    .COUT(\c$1864 ),
    .SUM(\s$1865 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_95_0 (.A(pp_row95_3),
    .B(pp_row95_4),
    .CIN(pp_row95_5),
    .COUT(\c$1866 ),
    .SUM(\s$1867 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_95_1 (.A(pp_row95_6),
    .B(pp_row95_7),
    .CIN(pp_row95_8),
    .COUT(\c$1868 ),
    .SUM(\s$1869 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_95_2 (.A(pp_row95_9),
    .B(pp_row95_10),
    .CIN(pp_row95_11),
    .COUT(\c$1870 ),
    .SUM(\s$1871 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_95_3 (.A(pp_row95_12),
    .B(pp_row95_13),
    .CIN(pp_row95_14),
    .COUT(\c$1872 ),
    .SUM(\s$1873 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_95_4 (.A(pp_row95_15),
    .B(pp_row95_16),
    .CIN(pp_row95_17),
    .COUT(\c$1874 ),
    .SUM(\s$1875 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_95_5 (.A(pp_row95_18),
    .B(\c$1042 ),
    .CIN(\c$1044 ),
    .COUT(\c$1876 ),
    .SUM(\s$1877 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_96_0 (.A(pp_row96_2),
    .B(pp_row96_3),
    .CIN(pp_row96_4),
    .COUT(\c$1878 ),
    .SUM(\s$1879 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_96_1 (.A(pp_row96_5),
    .B(pp_row96_6),
    .CIN(pp_row96_7),
    .COUT(\c$1880 ),
    .SUM(\s$1881 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_96_2 (.A(pp_row96_8),
    .B(pp_row96_9),
    .CIN(pp_row96_10),
    .COUT(\c$1882 ),
    .SUM(\s$1883 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_96_3 (.A(pp_row96_11),
    .B(pp_row96_12),
    .CIN(pp_row96_13),
    .COUT(\c$1884 ),
    .SUM(\s$1885 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_96_4 (.A(pp_row96_14),
    .B(pp_row96_15),
    .CIN(pp_row96_16),
    .COUT(\c$1886 ),
    .SUM(\s$1887 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_96_5 (.A(pp_row96_17),
    .B(pp_row96_18),
    .CIN(\c$1046 ),
    .COUT(\c$1888 ),
    .SUM(\s$1889 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_97_0 (.A(pp_row97_0),
    .B(pp_row97_1),
    .CIN(pp_row97_2),
    .COUT(\c$1890 ),
    .SUM(\s$1891 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_97_1 (.A(pp_row97_3),
    .B(pp_row97_4),
    .CIN(pp_row97_5),
    .COUT(\c$1892 ),
    .SUM(\s$1893 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_97_2 (.A(pp_row97_6),
    .B(pp_row97_7),
    .CIN(pp_row97_8),
    .COUT(\c$1894 ),
    .SUM(\s$1895 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_97_3 (.A(pp_row97_9),
    .B(pp_row97_10),
    .CIN(pp_row97_11),
    .COUT(\c$1896 ),
    .SUM(\s$1897 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_97_4 (.A(pp_row97_12),
    .B(pp_row97_13),
    .CIN(pp_row97_14),
    .COUT(\c$1898 ),
    .SUM(\s$1899 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_97_5 (.A(pp_row97_15),
    .B(pp_row97_16),
    .CIN(pp_row97_17),
    .COUT(\c$1900 ),
    .SUM(\s$1901 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_98_0 (.A(net1908),
    .B(pp_row98_1),
    .CIN(pp_row98_2),
    .COUT(\c$1902 ),
    .SUM(\s$1903 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_98_1 (.A(pp_row98_3),
    .B(pp_row98_4),
    .CIN(pp_row98_5),
    .COUT(\c$1904 ),
    .SUM(\s$1905 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_98_2 (.A(pp_row98_6),
    .B(pp_row98_7),
    .CIN(pp_row98_8),
    .COUT(\c$1906 ),
    .SUM(\s$1907 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_98_3 (.A(pp_row98_9),
    .B(pp_row98_10),
    .CIN(pp_row98_11),
    .COUT(\c$1908 ),
    .SUM(\s$1909 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_98_4 (.A(pp_row98_12),
    .B(pp_row98_13),
    .CIN(pp_row98_14),
    .COUT(\c$1910 ),
    .SUM(\s$1911 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_99_0 (.A(pp_row99_0),
    .B(pp_row99_1),
    .CIN(pp_row99_2),
    .COUT(\c$1914 ),
    .SUM(\s$1915 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_99_1 (.A(pp_row99_3),
    .B(pp_row99_4),
    .CIN(pp_row99_5),
    .COUT(\c$1916 ),
    .SUM(\s$1917 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_99_2 (.A(pp_row99_6),
    .B(pp_row99_7),
    .CIN(pp_row99_8),
    .COUT(\c$1918 ),
    .SUM(\s$1919 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_2_99_3 (.A(pp_row99_9),
    .B(pp_row99_10),
    .CIN(pp_row99_11),
    .COUT(\c$1920 ),
    .SUM(\s$1921 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_2_99_4 (.A(pp_row99_12),
    .B(pp_row99_13),
    .CIN(pp_row99_14),
    .COUT(\c$1922 ),
    .SUM(\s$1923 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_100_0 (.A(pp_row100_14),
    .B(pp_row100_15),
    .CIN(pp_row100_16),
    .COUT(\c$2638 ),
    .SUM(\s$2639 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_100_1 (.A(\c$1914 ),
    .B(\c$1916 ),
    .CIN(\c$1918 ),
    .COUT(\c$2640 ),
    .SUM(\s$2641 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_100_2 (.A(\c$1920 ),
    .B(\c$1922 ),
    .CIN(\s$1925 ),
    .COUT(\c$2642 ),
    .SUM(\s$2643 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_100_3 (.A(\s$1927 ),
    .B(\s$1929 ),
    .CIN(\s$1931 ),
    .COUT(\c$2644 ),
    .SUM(\s$2645 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_101_0 (.A(pp_row101_12),
    .B(pp_row101_13),
    .CIN(pp_row101_14),
    .COUT(\c$2646 ),
    .SUM(\s$2647 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_101_1 (.A(pp_row101_15),
    .B(\c$1924 ),
    .CIN(\c$1926 ),
    .COUT(\c$2648 ),
    .SUM(\s$2649 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_101_2 (.A(\c$1928 ),
    .B(\c$1930 ),
    .CIN(\c$1932 ),
    .COUT(\c$2650 ),
    .SUM(\s$2651 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_101_3 (.A(\s$1935 ),
    .B(\s$1937 ),
    .CIN(\s$1939 ),
    .COUT(\c$2652 ),
    .SUM(\s$2653 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_102_0 (.A(pp_row102_11),
    .B(pp_row102_12),
    .CIN(pp_row102_13),
    .COUT(\c$2654 ),
    .SUM(\s$2655 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_102_1 (.A(pp_row102_14),
    .B(pp_row102_15),
    .CIN(\c$1934 ),
    .COUT(\c$2656 ),
    .SUM(\s$2657 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_102_2 (.A(\c$1936 ),
    .B(\c$1938 ),
    .CIN(\c$1940 ),
    .COUT(\c$2658 ),
    .SUM(\s$2659 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_102_3 (.A(\s$1943 ),
    .B(\s$1945 ),
    .CIN(\s$1947 ),
    .COUT(\c$2660 ),
    .SUM(\s$2661 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_103_0 (.A(pp_row103_9),
    .B(pp_row103_10),
    .CIN(pp_row103_11),
    .COUT(\c$2662 ),
    .SUM(\s$2663 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_103_1 (.A(pp_row103_12),
    .B(pp_row103_13),
    .CIN(pp_row103_14),
    .COUT(\c$2664 ),
    .SUM(\s$2665 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_103_2 (.A(\c$1942 ),
    .B(\c$1944 ),
    .CIN(\c$1946 ),
    .COUT(\c$2666 ),
    .SUM(\s$2667 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_103_3 (.A(\c$1948 ),
    .B(\s$1951 ),
    .CIN(\s$1953 ),
    .COUT(\c$2668 ),
    .SUM(\s$2669 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_104_0 (.A(pp_row104_8),
    .B(pp_row104_9),
    .CIN(pp_row104_10),
    .COUT(\c$2670 ),
    .SUM(\s$2671 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_104_1 (.A(pp_row104_11),
    .B(pp_row104_12),
    .CIN(pp_row104_13),
    .COUT(\c$2672 ),
    .SUM(\s$2673 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_104_2 (.A(pp_row104_14),
    .B(\c$1950 ),
    .CIN(\c$1952 ),
    .COUT(\c$2674 ),
    .SUM(\s$2675 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_104_3 (.A(\c$1954 ),
    .B(\s$1957 ),
    .CIN(\s$1959 ),
    .COUT(\c$2676 ),
    .SUM(\s$2677 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_105_0 (.A(pp_row105_6),
    .B(pp_row105_7),
    .CIN(pp_row105_8),
    .COUT(\c$2678 ),
    .SUM(\s$2679 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_105_1 (.A(pp_row105_9),
    .B(pp_row105_10),
    .CIN(pp_row105_11),
    .COUT(\c$2680 ),
    .SUM(\s$2681 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_105_2 (.A(pp_row105_12),
    .B(pp_row105_13),
    .CIN(\c$1956 ),
    .COUT(\c$2682 ),
    .SUM(\s$2683 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_105_3 (.A(\c$1958 ),
    .B(\c$1960 ),
    .CIN(\s$1963 ),
    .COUT(\c$2684 ),
    .SUM(\s$2685 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_106_0 (.A(pp_row106_5),
    .B(pp_row106_6),
    .CIN(pp_row106_7),
    .COUT(\c$2686 ),
    .SUM(\s$2687 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_106_1 (.A(pp_row106_8),
    .B(pp_row106_9),
    .CIN(pp_row106_10),
    .COUT(\c$2688 ),
    .SUM(\s$2689 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_106_2 (.A(pp_row106_11),
    .B(pp_row106_12),
    .CIN(pp_row106_13),
    .COUT(\c$2690 ),
    .SUM(\s$2691 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_106_3 (.A(\c$1962 ),
    .B(\c$1964 ),
    .CIN(\s$1967 ),
    .COUT(\c$2692 ),
    .SUM(\s$2693 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_107_0 (.A(pp_row107_3),
    .B(pp_row107_4),
    .CIN(pp_row107_5),
    .COUT(\c$2694 ),
    .SUM(\s$2695 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_107_1 (.A(pp_row107_6),
    .B(pp_row107_7),
    .CIN(pp_row107_8),
    .COUT(\c$2696 ),
    .SUM(\s$2697 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_107_2 (.A(pp_row107_9),
    .B(pp_row107_10),
    .CIN(pp_row107_11),
    .COUT(\c$2698 ),
    .SUM(\s$2699 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_107_3 (.A(pp_row107_12),
    .B(\c$1966 ),
    .CIN(\c$1968 ),
    .COUT(\c$2700 ),
    .SUM(\s$2701 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_108_0 (.A(pp_row108_2),
    .B(pp_row108_3),
    .CIN(pp_row108_4),
    .COUT(\c$2702 ),
    .SUM(\s$2703 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_108_1 (.A(pp_row108_5),
    .B(pp_row108_6),
    .CIN(pp_row108_7),
    .COUT(\c$2704 ),
    .SUM(\s$2705 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_108_2 (.A(pp_row108_8),
    .B(pp_row108_9),
    .CIN(pp_row108_10),
    .COUT(\c$2706 ),
    .SUM(\s$2707 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_108_3 (.A(pp_row108_11),
    .B(pp_row108_12),
    .CIN(\c$1970 ),
    .COUT(\c$2708 ),
    .SUM(\s$2709 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_109_0 (.A(pp_row109_0),
    .B(pp_row109_1),
    .CIN(pp_row109_2),
    .COUT(\c$2710 ),
    .SUM(\s$2711 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_109_1 (.A(pp_row109_3),
    .B(pp_row109_4),
    .CIN(pp_row109_5),
    .COUT(\c$2712 ),
    .SUM(\s$2713 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_109_2 (.A(pp_row109_6),
    .B(pp_row109_7),
    .CIN(pp_row109_8),
    .COUT(\c$2714 ),
    .SUM(\s$2715 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_109_3 (.A(pp_row109_9),
    .B(pp_row109_10),
    .CIN(pp_row109_11),
    .COUT(\c$2716 ),
    .SUM(\s$2717 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_110_0 (.A(net1909),
    .B(pp_row110_1),
    .CIN(pp_row110_2),
    .COUT(\c$2718 ),
    .SUM(\s$2719 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_110_1 (.A(pp_row110_3),
    .B(pp_row110_4),
    .CIN(pp_row110_5),
    .COUT(\c$2720 ),
    .SUM(\s$2721 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_110_2 (.A(pp_row110_6),
    .B(pp_row110_7),
    .CIN(pp_row110_8),
    .COUT(\c$2722 ),
    .SUM(\s$2723 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_111_0 (.A(pp_row111_0),
    .B(pp_row111_1),
    .CIN(pp_row111_2),
    .COUT(\c$2726 ),
    .SUM(\s$2727 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_111_1 (.A(pp_row111_3),
    .B(pp_row111_4),
    .CIN(pp_row111_5),
    .COUT(\c$2728 ),
    .SUM(\s$2729 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_111_2 (.A(pp_row111_6),
    .B(pp_row111_7),
    .CIN(pp_row111_8),
    .COUT(\c$2730 ),
    .SUM(\s$2731 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_112_0 (.A(net1910),
    .B(pp_row112_1),
    .CIN(pp_row112_2),
    .COUT(\c$2732 ),
    .SUM(\s$2733 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_112_1 (.A(pp_row112_3),
    .B(pp_row112_4),
    .CIN(pp_row112_5),
    .COUT(\c$2734 ),
    .SUM(\s$2735 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_113_0 (.A(pp_row113_0),
    .B(pp_row113_1),
    .CIN(pp_row113_2),
    .COUT(\c$2738 ),
    .SUM(\s$2739 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_113_1 (.A(pp_row113_3),
    .B(pp_row113_4),
    .CIN(pp_row113_5),
    .COUT(\c$2740 ),
    .SUM(\s$2741 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_114_0 (.A(net1911),
    .B(pp_row114_1),
    .CIN(pp_row114_2),
    .COUT(\c$2742 ),
    .SUM(\s$2743 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_115_0 (.A(pp_row115_0),
    .B(pp_row115_1),
    .CIN(pp_row115_2),
    .COUT(\c$2746 ),
    .SUM(\s$2747 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_16_0 (.A(pp_row16_0),
    .B(pp_row16_1),
    .CIN(pp_row16_2),
    .COUT(\c$1978 ),
    .SUM(\s$1979 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_17_0 (.A(pp_row17_0),
    .B(pp_row17_1),
    .CIN(pp_row17_2),
    .COUT(\c$1982 ),
    .SUM(\s$1983 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_18_0 (.A(pp_row18_0),
    .B(pp_row18_1),
    .CIN(pp_row18_2),
    .COUT(\c$1986 ),
    .SUM(\s$1987 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_18_1 (.A(pp_row18_3),
    .B(pp_row18_4),
    .CIN(pp_row18_5),
    .COUT(\c$1988 ),
    .SUM(\s$1989 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_19_0 (.A(pp_row19_0),
    .B(pp_row19_1),
    .CIN(pp_row19_2),
    .COUT(\c$1992 ),
    .SUM(\s$1993 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_19_1 (.A(pp_row19_3),
    .B(pp_row19_4),
    .CIN(pp_row19_5),
    .COUT(\c$1994 ),
    .SUM(\s$1995 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_20_0 (.A(pp_row20_0),
    .B(pp_row20_1),
    .CIN(pp_row20_2),
    .COUT(\c$1998 ),
    .SUM(\s$1999 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_20_1 (.A(pp_row20_3),
    .B(pp_row20_4),
    .CIN(pp_row20_5),
    .COUT(\c$2000 ),
    .SUM(\s$2001 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_20_2 (.A(pp_row20_6),
    .B(pp_row20_7),
    .CIN(pp_row20_8),
    .COUT(\c$2002 ),
    .SUM(\s$2003 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_21_0 (.A(pp_row21_0),
    .B(pp_row21_1),
    .CIN(pp_row21_2),
    .COUT(\c$2006 ),
    .SUM(\s$2007 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_21_1 (.A(pp_row21_3),
    .B(pp_row21_4),
    .CIN(pp_row21_5),
    .COUT(\c$2008 ),
    .SUM(\s$2009 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_21_2 (.A(pp_row21_6),
    .B(pp_row21_7),
    .CIN(pp_row21_8),
    .COUT(\c$2010 ),
    .SUM(\s$2011 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_22_0 (.A(pp_row22_2),
    .B(pp_row22_3),
    .CIN(pp_row22_4),
    .COUT(\c$2014 ),
    .SUM(\s$2015 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_22_1 (.A(pp_row22_5),
    .B(pp_row22_6),
    .CIN(pp_row22_7),
    .COUT(\c$2016 ),
    .SUM(\s$2017 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_22_2 (.A(pp_row22_8),
    .B(pp_row22_9),
    .CIN(pp_row22_10),
    .COUT(\c$2018 ),
    .SUM(\s$2019 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_22_3 (.A(pp_row22_11),
    .B(pp_row22_12),
    .CIN(pp_row22_13),
    .COUT(\c$2020 ),
    .SUM(\s$2021 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_23_0 (.A(pp_row23_2),
    .B(pp_row23_3),
    .CIN(pp_row23_4),
    .COUT(\c$2022 ),
    .SUM(\s$2023 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_23_1 (.A(pp_row23_5),
    .B(pp_row23_6),
    .CIN(pp_row23_7),
    .COUT(\c$2024 ),
    .SUM(\s$2025 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_23_2 (.A(pp_row23_8),
    .B(pp_row23_9),
    .CIN(pp_row23_10),
    .COUT(\c$2026 ),
    .SUM(\s$2027 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_23_3 (.A(pp_row23_11),
    .B(pp_row23_12),
    .CIN(\c$1050 ),
    .COUT(\c$2028 ),
    .SUM(\s$2029 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_24_0 (.A(pp_row24_5),
    .B(pp_row24_6),
    .CIN(pp_row24_7),
    .COUT(\c$2030 ),
    .SUM(\s$2031 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_24_1 (.A(pp_row24_8),
    .B(pp_row24_9),
    .CIN(pp_row24_10),
    .COUT(\c$2032 ),
    .SUM(\s$2033 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_24_2 (.A(pp_row24_11),
    .B(pp_row24_12),
    .CIN(pp_row24_13),
    .COUT(\c$2034 ),
    .SUM(\s$2035 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_24_3 (.A(pp_row24_14),
    .B(\c$1052 ),
    .CIN(\s$1055 ),
    .COUT(\c$2036 ),
    .SUM(\s$2037 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_25_0 (.A(pp_row25_5),
    .B(pp_row25_6),
    .CIN(pp_row25_7),
    .COUT(\c$2038 ),
    .SUM(\s$2039 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_25_1 (.A(pp_row25_8),
    .B(pp_row25_9),
    .CIN(pp_row25_10),
    .COUT(\c$2040 ),
    .SUM(\s$2041 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_25_2 (.A(pp_row25_11),
    .B(pp_row25_12),
    .CIN(pp_row25_13),
    .COUT(\c$2042 ),
    .SUM(\s$2043 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_25_3 (.A(\c$1054 ),
    .B(\c$1056 ),
    .CIN(\s$1059 ),
    .COUT(\c$2044 ),
    .SUM(\s$2045 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_26_0 (.A(pp_row26_8),
    .B(pp_row26_9),
    .CIN(pp_row26_10),
    .COUT(\c$2046 ),
    .SUM(\s$2047 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_26_1 (.A(pp_row26_11),
    .B(pp_row26_12),
    .CIN(pp_row26_13),
    .COUT(\c$2048 ),
    .SUM(\s$2049 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_26_2 (.A(pp_row26_14),
    .B(pp_row26_15),
    .CIN(\c$1058 ),
    .COUT(\c$2050 ),
    .SUM(\s$2051 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_26_3 (.A(\c$1060 ),
    .B(\s$1063 ),
    .CIN(\s$1065 ),
    .COUT(\c$2052 ),
    .SUM(\s$2053 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_27_0 (.A(pp_row27_8),
    .B(pp_row27_9),
    .CIN(pp_row27_10),
    .COUT(\c$2054 ),
    .SUM(\s$2055 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_27_1 (.A(pp_row27_11),
    .B(pp_row27_12),
    .CIN(pp_row27_13),
    .COUT(\c$2056 ),
    .SUM(\s$2057 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_27_2 (.A(pp_row27_14),
    .B(\c$1062 ),
    .CIN(\c$1064 ),
    .COUT(\c$2058 ),
    .SUM(\s$2059 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_27_3 (.A(\c$1066 ),
    .B(\s$1069 ),
    .CIN(\s$1071 ),
    .COUT(\c$2060 ),
    .SUM(\s$2061 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_28_0 (.A(pp_row28_11),
    .B(pp_row28_12),
    .CIN(pp_row28_13),
    .COUT(\c$2062 ),
    .SUM(\s$2063 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_28_1 (.A(pp_row28_14),
    .B(pp_row28_15),
    .CIN(pp_row28_16),
    .COUT(\c$2064 ),
    .SUM(\s$2065 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_28_2 (.A(\c$1068 ),
    .B(\c$1070 ),
    .CIN(\c$1072 ),
    .COUT(\c$2066 ),
    .SUM(\s$2067 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_28_3 (.A(\s$1075 ),
    .B(\s$1077 ),
    .CIN(\s$1079 ),
    .COUT(\c$2068 ),
    .SUM(\s$2069 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_29_0 (.A(pp_row29_11),
    .B(pp_row29_12),
    .CIN(pp_row29_13),
    .COUT(\c$2070 ),
    .SUM(\s$2071 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_29_1 (.A(pp_row29_14),
    .B(pp_row29_15),
    .CIN(\c$1074 ),
    .COUT(\c$2072 ),
    .SUM(\s$2073 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_29_2 (.A(\c$1076 ),
    .B(\c$1078 ),
    .CIN(\c$1080 ),
    .COUT(\c$2074 ),
    .SUM(\s$2075 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_29_3 (.A(\s$1083 ),
    .B(\s$1085 ),
    .CIN(\s$1087 ),
    .COUT(\c$2076 ),
    .SUM(\s$2077 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_30_0 (.A(pp_row30_14),
    .B(pp_row30_15),
    .CIN(pp_row30_16),
    .COUT(\c$2078 ),
    .SUM(\s$2079 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_30_1 (.A(pp_row30_17),
    .B(\c$1082 ),
    .CIN(\c$1084 ),
    .COUT(\c$2080 ),
    .SUM(\s$2081 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_30_2 (.A(\c$1086 ),
    .B(\c$1088 ),
    .CIN(\s$1091 ),
    .COUT(\c$2082 ),
    .SUM(\s$2083 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_30_3 (.A(\s$1093 ),
    .B(\s$1095 ),
    .CIN(\s$1097 ),
    .COUT(\c$2084 ),
    .SUM(\s$2085 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_31_0 (.A(pp_row31_14),
    .B(pp_row31_15),
    .CIN(pp_row31_16),
    .COUT(\c$2086 ),
    .SUM(\s$2087 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_31_1 (.A(\c$1090 ),
    .B(\c$1092 ),
    .CIN(\c$1094 ),
    .COUT(\c$2088 ),
    .SUM(\s$2089 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_31_2 (.A(\c$1096 ),
    .B(\c$1098 ),
    .CIN(\s$1101 ),
    .COUT(\c$2090 ),
    .SUM(\s$2091 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_31_3 (.A(\s$1103 ),
    .B(\s$1105 ),
    .CIN(\s$1107 ),
    .COUT(\c$2092 ),
    .SUM(\s$2093 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_32_0 (.A(pp_row32_17),
    .B(pp_row32_18),
    .CIN(\c$1100 ),
    .COUT(\c$2094 ),
    .SUM(\s$2095 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_32_1 (.A(\c$1102 ),
    .B(\c$1104 ),
    .CIN(\c$1106 ),
    .COUT(\c$2096 ),
    .SUM(\s$2097 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_32_2 (.A(\c$1108 ),
    .B(\s$1111 ),
    .CIN(\s$1113 ),
    .COUT(\c$2098 ),
    .SUM(\s$2099 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_32_3 (.A(\s$1115 ),
    .B(\s$1117 ),
    .CIN(\s$1119 ),
    .COUT(\c$2100 ),
    .SUM(\s$2101 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_33_0 (.A(pp_row33_17),
    .B(\c$1110 ),
    .CIN(\c$1112 ),
    .COUT(\c$2102 ),
    .SUM(\s$2103 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_33_1 (.A(\c$1114 ),
    .B(\c$1116 ),
    .CIN(\c$1118 ),
    .COUT(\c$2104 ),
    .SUM(\s$2105 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_33_2 (.A(\c$1120 ),
    .B(\s$1123 ),
    .CIN(\s$1125 ),
    .COUT(\c$2106 ),
    .SUM(\s$2107 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_33_3 (.A(\s$1127 ),
    .B(\s$1129 ),
    .CIN(\s$1131 ),
    .COUT(\c$2108 ),
    .SUM(\s$2109 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_34_0 (.A(\s$205 ),
    .B(\c$1122 ),
    .CIN(\c$1124 ),
    .COUT(\c$2110 ),
    .SUM(\s$2111 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_34_1 (.A(\c$1126 ),
    .B(\c$1128 ),
    .CIN(\c$1130 ),
    .COUT(\c$2112 ),
    .SUM(\s$2113 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_34_2 (.A(\c$1132 ),
    .B(\s$1135 ),
    .CIN(\s$1137 ),
    .COUT(\c$2114 ),
    .SUM(\s$2115 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_34_3 (.A(\s$1139 ),
    .B(\s$1141 ),
    .CIN(\s$1143 ),
    .COUT(\c$2116 ),
    .SUM(\s$2117 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_35_0 (.A(\s$207 ),
    .B(\c$1134 ),
    .CIN(\c$1136 ),
    .COUT(\c$2118 ),
    .SUM(\s$2119 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_35_1 (.A(\c$1138 ),
    .B(\c$1140 ),
    .CIN(\c$1142 ),
    .COUT(\c$2120 ),
    .SUM(\s$2121 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_35_2 (.A(\c$1144 ),
    .B(\s$1147 ),
    .CIN(\s$1149 ),
    .COUT(\c$2122 ),
    .SUM(\s$2123 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_35_3 (.A(\s$1151 ),
    .B(\s$1153 ),
    .CIN(\s$1155 ),
    .COUT(\c$2124 ),
    .SUM(\s$2125 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_36_0 (.A(\s$211 ),
    .B(\c$1146 ),
    .CIN(\c$1148 ),
    .COUT(\c$2126 ),
    .SUM(\s$2127 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_36_1 (.A(\c$1150 ),
    .B(\c$1152 ),
    .CIN(\c$1154 ),
    .COUT(\c$2128 ),
    .SUM(\s$2129 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_36_2 (.A(\c$1156 ),
    .B(\s$1159 ),
    .CIN(\s$1161 ),
    .COUT(\c$2130 ),
    .SUM(\s$2131 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_36_3 (.A(\s$1163 ),
    .B(\s$1165 ),
    .CIN(\s$1167 ),
    .COUT(\c$2132 ),
    .SUM(\s$2133 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_37_0 (.A(\s$215 ),
    .B(\c$1158 ),
    .CIN(\c$1160 ),
    .COUT(\c$2134 ),
    .SUM(\s$2135 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_37_1 (.A(\c$1162 ),
    .B(\c$1164 ),
    .CIN(\c$1166 ),
    .COUT(\c$2136 ),
    .SUM(\s$2137 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_37_2 (.A(\c$1168 ),
    .B(\s$1171 ),
    .CIN(\s$1173 ),
    .COUT(\c$2138 ),
    .SUM(\s$2139 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_37_3 (.A(\s$1175 ),
    .B(\s$1177 ),
    .CIN(\s$1179 ),
    .COUT(\c$2140 ),
    .SUM(\s$2141 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_38_0 (.A(\s$221 ),
    .B(\c$1170 ),
    .CIN(\c$1172 ),
    .COUT(\c$2142 ),
    .SUM(\s$2143 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_38_1 (.A(\c$1174 ),
    .B(\c$1176 ),
    .CIN(\c$1178 ),
    .COUT(\c$2144 ),
    .SUM(\s$2145 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_38_2 (.A(\c$1180 ),
    .B(\s$1183 ),
    .CIN(\s$1185 ),
    .COUT(\c$2146 ),
    .SUM(\s$2147 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_38_3 (.A(\s$1187 ),
    .B(\s$1189 ),
    .CIN(\s$1191 ),
    .COUT(\c$2148 ),
    .SUM(\s$2149 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_39_0 (.A(\s$227 ),
    .B(\c$1182 ),
    .CIN(\c$1184 ),
    .COUT(\c$2150 ),
    .SUM(\s$2151 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_39_1 (.A(\c$1186 ),
    .B(\c$1188 ),
    .CIN(\c$1190 ),
    .COUT(\c$2152 ),
    .SUM(\s$2153 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_39_2 (.A(\c$1192 ),
    .B(\s$1195 ),
    .CIN(\s$1197 ),
    .COUT(\c$2154 ),
    .SUM(\s$2155 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_39_3 (.A(\s$1199 ),
    .B(\s$1201 ),
    .CIN(\s$1203 ),
    .COUT(\c$2156 ),
    .SUM(\s$2157 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_40_0 (.A(\s$235 ),
    .B(\c$1194 ),
    .CIN(\c$1196 ),
    .COUT(\c$2158 ),
    .SUM(\s$2159 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_40_1 (.A(\c$1198 ),
    .B(\c$1200 ),
    .CIN(\c$1202 ),
    .COUT(\c$2160 ),
    .SUM(\s$2161 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_40_2 (.A(\c$1204 ),
    .B(\s$1207 ),
    .CIN(\s$1209 ),
    .COUT(\c$2162 ),
    .SUM(\s$2163 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_40_3 (.A(\s$1211 ),
    .B(\s$1213 ),
    .CIN(\s$1215 ),
    .COUT(\c$2164 ),
    .SUM(\s$2165 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_41_0 (.A(\s$243 ),
    .B(\c$1206 ),
    .CIN(\c$1208 ),
    .COUT(\c$2166 ),
    .SUM(\s$2167 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_41_1 (.A(\c$1210 ),
    .B(\c$1212 ),
    .CIN(\c$1214 ),
    .COUT(\c$2168 ),
    .SUM(\s$2169 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_41_2 (.A(\c$1216 ),
    .B(\s$1219 ),
    .CIN(\s$1221 ),
    .COUT(\c$2170 ),
    .SUM(\s$2171 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_41_3 (.A(\s$1223 ),
    .B(\s$1225 ),
    .CIN(\s$1227 ),
    .COUT(\c$2172 ),
    .SUM(\s$2173 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_42_0 (.A(\s$253 ),
    .B(\c$1218 ),
    .CIN(\c$1220 ),
    .COUT(\c$2174 ),
    .SUM(\s$2175 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_42_1 (.A(\c$1222 ),
    .B(\c$1224 ),
    .CIN(\c$1226 ),
    .COUT(\c$2176 ),
    .SUM(\s$2177 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_42_2 (.A(\c$1228 ),
    .B(\s$1231 ),
    .CIN(\s$1233 ),
    .COUT(\c$2178 ),
    .SUM(\s$2179 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_42_3 (.A(\s$1235 ),
    .B(\s$1237 ),
    .CIN(\s$1239 ),
    .COUT(\c$2180 ),
    .SUM(\s$2181 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_43_0 (.A(\s$263 ),
    .B(\c$1230 ),
    .CIN(\c$1232 ),
    .COUT(\c$2182 ),
    .SUM(\s$2183 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_43_1 (.A(\c$1234 ),
    .B(\c$1236 ),
    .CIN(\c$1238 ),
    .COUT(\c$2184 ),
    .SUM(\s$2185 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_43_2 (.A(\c$1240 ),
    .B(\s$1243 ),
    .CIN(\s$1245 ),
    .COUT(\c$2186 ),
    .SUM(\s$2187 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_43_3 (.A(\s$1247 ),
    .B(\s$1249 ),
    .CIN(\s$1251 ),
    .COUT(\c$2188 ),
    .SUM(\s$2189 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_44_0 (.A(\s$275 ),
    .B(\c$1242 ),
    .CIN(\c$1244 ),
    .COUT(\c$2190 ),
    .SUM(\s$2191 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_44_1 (.A(\c$1246 ),
    .B(\c$1248 ),
    .CIN(\c$1250 ),
    .COUT(\c$2192 ),
    .SUM(\s$2193 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_44_2 (.A(\c$1252 ),
    .B(\s$1255 ),
    .CIN(\s$1257 ),
    .COUT(\c$2194 ),
    .SUM(\s$2195 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_44_3 (.A(\s$1259 ),
    .B(\s$1261 ),
    .CIN(\s$1263 ),
    .COUT(\c$2196 ),
    .SUM(\s$2197 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_45_0 (.A(\s$287 ),
    .B(\c$1254 ),
    .CIN(\c$1256 ),
    .COUT(\c$2198 ),
    .SUM(\s$2199 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_45_1 (.A(\c$1258 ),
    .B(\c$1260 ),
    .CIN(\c$1262 ),
    .COUT(\c$2200 ),
    .SUM(\s$2201 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_45_2 (.A(\c$1264 ),
    .B(\s$1267 ),
    .CIN(\s$1269 ),
    .COUT(\c$2202 ),
    .SUM(\s$2203 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_45_3 (.A(\s$1271 ),
    .B(\s$1273 ),
    .CIN(\s$1275 ),
    .COUT(\c$2204 ),
    .SUM(\s$2205 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_46_0 (.A(\s$301 ),
    .B(\c$1266 ),
    .CIN(\c$1268 ),
    .COUT(\c$2206 ),
    .SUM(\s$2207 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_46_1 (.A(\c$1270 ),
    .B(\c$1272 ),
    .CIN(\c$1274 ),
    .COUT(\c$2208 ),
    .SUM(\s$2209 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_46_2 (.A(\c$1276 ),
    .B(\s$1279 ),
    .CIN(\s$1281 ),
    .COUT(\c$2210 ),
    .SUM(\s$2211 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_46_3 (.A(\s$1283 ),
    .B(\s$1285 ),
    .CIN(\s$1287 ),
    .COUT(\c$2212 ),
    .SUM(\s$2213 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_47_0 (.A(\s$315 ),
    .B(\c$1278 ),
    .CIN(\c$1280 ),
    .COUT(\c$2214 ),
    .SUM(\s$2215 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_47_1 (.A(\c$1282 ),
    .B(\c$1284 ),
    .CIN(\c$1286 ),
    .COUT(\c$2216 ),
    .SUM(\s$2217 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_47_2 (.A(\c$1288 ),
    .B(\s$1291 ),
    .CIN(\s$1293 ),
    .COUT(\c$2218 ),
    .SUM(\s$2219 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_47_3 (.A(\s$1295 ),
    .B(\s$1297 ),
    .CIN(\s$1299 ),
    .COUT(\c$2220 ),
    .SUM(\s$2221 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_48_0 (.A(\s$331 ),
    .B(\c$1290 ),
    .CIN(\c$1292 ),
    .COUT(\c$2222 ),
    .SUM(\s$2223 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_48_1 (.A(\c$1294 ),
    .B(\c$1296 ),
    .CIN(\c$1298 ),
    .COUT(\c$2224 ),
    .SUM(\s$2225 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_48_2 (.A(\c$1300 ),
    .B(\s$1303 ),
    .CIN(\s$1305 ),
    .COUT(\c$2226 ),
    .SUM(\s$2227 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_48_3 (.A(\s$1307 ),
    .B(\s$1309 ),
    .CIN(\s$1311 ),
    .COUT(\c$2228 ),
    .SUM(\s$2229 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_49_0 (.A(\s$347 ),
    .B(\c$1302 ),
    .CIN(\c$1304 ),
    .COUT(\c$2230 ),
    .SUM(\s$2231 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_49_1 (.A(\c$1306 ),
    .B(\c$1308 ),
    .CIN(\c$1310 ),
    .COUT(\c$2232 ),
    .SUM(\s$2233 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_49_2 (.A(\c$1312 ),
    .B(\s$1315 ),
    .CIN(\s$1317 ),
    .COUT(\c$2234 ),
    .SUM(\s$2235 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_49_3 (.A(\s$1319 ),
    .B(\s$1321 ),
    .CIN(\s$1323 ),
    .COUT(\c$2236 ),
    .SUM(\s$2237 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_50_0 (.A(\s$365 ),
    .B(\c$1314 ),
    .CIN(\c$1316 ),
    .COUT(\c$2238 ),
    .SUM(\s$2239 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_50_1 (.A(\c$1318 ),
    .B(\c$1320 ),
    .CIN(\c$1322 ),
    .COUT(\c$2240 ),
    .SUM(\s$2241 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_50_2 (.A(\c$1324 ),
    .B(\s$1327 ),
    .CIN(\s$1329 ),
    .COUT(\c$2242 ),
    .SUM(\s$2243 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_50_3 (.A(\s$1331 ),
    .B(\s$1333 ),
    .CIN(\s$1335 ),
    .COUT(\c$2244 ),
    .SUM(\s$2245 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_51_0 (.A(\s$383 ),
    .B(\c$1326 ),
    .CIN(\c$1328 ),
    .COUT(\c$2246 ),
    .SUM(\s$2247 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_51_1 (.A(\c$1330 ),
    .B(\c$1332 ),
    .CIN(\c$1334 ),
    .COUT(\c$2248 ),
    .SUM(\s$2249 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_51_2 (.A(\c$1336 ),
    .B(\s$1339 ),
    .CIN(\s$1341 ),
    .COUT(\c$2250 ),
    .SUM(\s$2251 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_51_3 (.A(\s$1343 ),
    .B(\s$1345 ),
    .CIN(\s$1347 ),
    .COUT(\c$2252 ),
    .SUM(\s$2253 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_52_0 (.A(\s$401 ),
    .B(\c$1338 ),
    .CIN(\c$1340 ),
    .COUT(\c$2254 ),
    .SUM(\s$2255 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_52_1 (.A(\c$1342 ),
    .B(\c$1344 ),
    .CIN(\c$1346 ),
    .COUT(\c$2256 ),
    .SUM(\s$2257 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_52_2 (.A(\c$1348 ),
    .B(\s$1351 ),
    .CIN(\s$1353 ),
    .COUT(\c$2258 ),
    .SUM(\s$2259 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_52_3 (.A(\s$1355 ),
    .B(\s$1357 ),
    .CIN(\s$1359 ),
    .COUT(\c$2260 ),
    .SUM(\s$2261 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_53_0 (.A(\s$419 ),
    .B(\c$1350 ),
    .CIN(\c$1352 ),
    .COUT(\c$2262 ),
    .SUM(\s$2263 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_53_1 (.A(\c$1354 ),
    .B(\c$1356 ),
    .CIN(\c$1358 ),
    .COUT(\c$2264 ),
    .SUM(\s$2265 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_53_2 (.A(\c$1360 ),
    .B(\s$1363 ),
    .CIN(\s$1365 ),
    .COUT(\c$2266 ),
    .SUM(\s$2267 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_53_3 (.A(\s$1367 ),
    .B(\s$1369 ),
    .CIN(\s$1371 ),
    .COUT(\c$2268 ),
    .SUM(\s$2269 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_54_0 (.A(\s$437 ),
    .B(\c$1362 ),
    .CIN(\c$1364 ),
    .COUT(\c$2270 ),
    .SUM(\s$2271 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_54_1 (.A(\c$1366 ),
    .B(\c$1368 ),
    .CIN(\c$1370 ),
    .COUT(\c$2272 ),
    .SUM(\s$2273 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_54_2 (.A(\c$1372 ),
    .B(\s$1375 ),
    .CIN(\s$1377 ),
    .COUT(\c$2274 ),
    .SUM(\s$2275 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_54_3 (.A(\s$1379 ),
    .B(\s$1381 ),
    .CIN(\s$1383 ),
    .COUT(\c$2276 ),
    .SUM(\s$2277 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_55_0 (.A(\s$455 ),
    .B(\c$1374 ),
    .CIN(\c$1376 ),
    .COUT(\c$2278 ),
    .SUM(\s$2279 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_55_1 (.A(\c$1378 ),
    .B(\c$1380 ),
    .CIN(\c$1382 ),
    .COUT(\c$2280 ),
    .SUM(\s$2281 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_55_2 (.A(\c$1384 ),
    .B(\s$1387 ),
    .CIN(\s$1389 ),
    .COUT(\c$2282 ),
    .SUM(\s$2283 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_55_3 (.A(\s$1391 ),
    .B(\s$1393 ),
    .CIN(\s$1395 ),
    .COUT(\c$2284 ),
    .SUM(\s$2285 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_56_0 (.A(\s$473 ),
    .B(\c$1386 ),
    .CIN(\c$1388 ),
    .COUT(\c$2286 ),
    .SUM(\s$2287 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_56_1 (.A(\c$1390 ),
    .B(\c$1392 ),
    .CIN(\c$1394 ),
    .COUT(\c$2288 ),
    .SUM(\s$2289 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_56_2 (.A(\c$1396 ),
    .B(\s$1399 ),
    .CIN(\s$1401 ),
    .COUT(\c$2290 ),
    .SUM(\s$2291 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_56_3 (.A(\s$1403 ),
    .B(\s$1405 ),
    .CIN(\s$1407 ),
    .COUT(\c$2292 ),
    .SUM(\s$2293 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_57_0 (.A(\s$491 ),
    .B(\c$1398 ),
    .CIN(\c$1400 ),
    .COUT(\c$2294 ),
    .SUM(\s$2295 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_57_1 (.A(\c$1402 ),
    .B(\c$1404 ),
    .CIN(\c$1406 ),
    .COUT(\c$2296 ),
    .SUM(\s$2297 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_57_2 (.A(\c$1408 ),
    .B(\s$1411 ),
    .CIN(\s$1413 ),
    .COUT(\c$2298 ),
    .SUM(\s$2299 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_57_3 (.A(\s$1415 ),
    .B(\s$1417 ),
    .CIN(\s$1419 ),
    .COUT(\c$2300 ),
    .SUM(\s$2301 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_58_0 (.A(\s$509 ),
    .B(\c$1410 ),
    .CIN(\c$1412 ),
    .COUT(\c$2302 ),
    .SUM(\s$2303 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_58_1 (.A(\c$1414 ),
    .B(\c$1416 ),
    .CIN(\c$1418 ),
    .COUT(\c$2304 ),
    .SUM(\s$2305 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_58_2 (.A(\c$1420 ),
    .B(\s$1423 ),
    .CIN(\s$1425 ),
    .COUT(\c$2306 ),
    .SUM(\s$2307 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_58_3 (.A(\s$1427 ),
    .B(\s$1429 ),
    .CIN(\s$1431 ),
    .COUT(\c$2308 ),
    .SUM(\s$2309 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_59_0 (.A(\s$527 ),
    .B(\c$1422 ),
    .CIN(\c$1424 ),
    .COUT(\c$2310 ),
    .SUM(\s$2311 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_59_1 (.A(\c$1426 ),
    .B(\c$1428 ),
    .CIN(\c$1430 ),
    .COUT(\c$2312 ),
    .SUM(\s$2313 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_59_2 (.A(\c$1432 ),
    .B(\s$1435 ),
    .CIN(\s$1437 ),
    .COUT(\c$2314 ),
    .SUM(\s$2315 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_59_3 (.A(\s$1439 ),
    .B(\s$1441 ),
    .CIN(\s$1443 ),
    .COUT(\c$2316 ),
    .SUM(\s$2317 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_60_0 (.A(\s$545 ),
    .B(\c$1434 ),
    .CIN(\c$1436 ),
    .COUT(\c$2318 ),
    .SUM(\s$2319 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_60_1 (.A(\c$1438 ),
    .B(\c$1440 ),
    .CIN(\c$1442 ),
    .COUT(\c$2320 ),
    .SUM(\s$2321 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_60_2 (.A(\c$1444 ),
    .B(\s$1447 ),
    .CIN(\s$1449 ),
    .COUT(\c$2322 ),
    .SUM(\s$2323 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_60_3 (.A(\s$1451 ),
    .B(\s$1453 ),
    .CIN(\s$1455 ),
    .COUT(\c$2324 ),
    .SUM(\s$2325 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_61_0 (.A(\s$563 ),
    .B(\c$1446 ),
    .CIN(\c$1448 ),
    .COUT(\c$2326 ),
    .SUM(\s$2327 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_61_1 (.A(\c$1450 ),
    .B(\c$1452 ),
    .CIN(\c$1454 ),
    .COUT(\c$2328 ),
    .SUM(\s$2329 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_61_2 (.A(\c$1456 ),
    .B(\s$1459 ),
    .CIN(\s$1461 ),
    .COUT(\c$2330 ),
    .SUM(\s$2331 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_61_3 (.A(\s$1463 ),
    .B(\s$1465 ),
    .CIN(\s$1467 ),
    .COUT(\c$2332 ),
    .SUM(\s$2333 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_62_0 (.A(\s$581 ),
    .B(\c$1458 ),
    .CIN(\c$1460 ),
    .COUT(\c$2334 ),
    .SUM(\s$2335 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_62_1 (.A(\c$1462 ),
    .B(\c$1464 ),
    .CIN(\c$1466 ),
    .COUT(\c$2336 ),
    .SUM(\s$2337 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_62_2 (.A(\c$1468 ),
    .B(\s$1471 ),
    .CIN(\s$1473 ),
    .COUT(\c$2338 ),
    .SUM(\s$2339 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_62_3 (.A(\s$1475 ),
    .B(\s$1477 ),
    .CIN(\s$1479 ),
    .COUT(\c$2340 ),
    .SUM(\s$2341 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_63_0 (.A(\s$599 ),
    .B(\c$1470 ),
    .CIN(\c$1472 ),
    .COUT(\c$2342 ),
    .SUM(\s$2343 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_63_1 (.A(\c$1474 ),
    .B(\c$1476 ),
    .CIN(\c$1478 ),
    .COUT(\c$2344 ),
    .SUM(\s$2345 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_63_2 (.A(\c$1480 ),
    .B(\s$1483 ),
    .CIN(\s$1485 ),
    .COUT(\c$2346 ),
    .SUM(\s$2347 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_63_3 (.A(\s$1487 ),
    .B(\s$1489 ),
    .CIN(\s$1491 ),
    .COUT(\c$2348 ),
    .SUM(\s$2349 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_64_0 (.A(\s$617 ),
    .B(\c$1482 ),
    .CIN(\c$1484 ),
    .COUT(\c$2350 ),
    .SUM(\s$2351 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_64_1 (.A(\c$1486 ),
    .B(\c$1488 ),
    .CIN(\c$1490 ),
    .COUT(\c$2352 ),
    .SUM(\s$2353 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_64_2 (.A(\c$1492 ),
    .B(\s$1495 ),
    .CIN(\s$1497 ),
    .COUT(\c$2354 ),
    .SUM(\s$2355 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_64_3 (.A(\s$1499 ),
    .B(\s$1501 ),
    .CIN(\s$1503 ),
    .COUT(\c$2356 ),
    .SUM(\s$2357 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_65_0 (.A(\s$635 ),
    .B(\c$1494 ),
    .CIN(\c$1496 ),
    .COUT(\c$2358 ),
    .SUM(\s$2359 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_65_1 (.A(\c$1498 ),
    .B(\c$1500 ),
    .CIN(\c$1502 ),
    .COUT(\c$2360 ),
    .SUM(\s$2361 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_65_2 (.A(\c$1504 ),
    .B(\s$1507 ),
    .CIN(\s$1509 ),
    .COUT(\c$2362 ),
    .SUM(\s$2363 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_65_3 (.A(\s$1511 ),
    .B(\s$1513 ),
    .CIN(\s$1515 ),
    .COUT(\c$2364 ),
    .SUM(\s$2365 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_66_0 (.A(\s$653 ),
    .B(\c$1506 ),
    .CIN(\c$1508 ),
    .COUT(\c$2366 ),
    .SUM(\s$2367 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_66_1 (.A(\c$1510 ),
    .B(\c$1512 ),
    .CIN(\c$1514 ),
    .COUT(\c$2368 ),
    .SUM(\s$2369 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_66_2 (.A(\c$1516 ),
    .B(\s$1519 ),
    .CIN(\s$1521 ),
    .COUT(\c$2370 ),
    .SUM(\s$2371 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_66_3 (.A(\s$1523 ),
    .B(\s$1525 ),
    .CIN(\s$1527 ),
    .COUT(\c$2372 ),
    .SUM(\s$2373 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_67_0 (.A(\s$671 ),
    .B(\c$1518 ),
    .CIN(\c$1520 ),
    .COUT(\c$2374 ),
    .SUM(\s$2375 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_67_1 (.A(\c$1522 ),
    .B(\c$1524 ),
    .CIN(\c$1526 ),
    .COUT(\c$2376 ),
    .SUM(\s$2377 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_67_2 (.A(\c$1528 ),
    .B(\s$1531 ),
    .CIN(\s$1533 ),
    .COUT(\c$2378 ),
    .SUM(\s$2379 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_67_3 (.A(\s$1535 ),
    .B(\s$1537 ),
    .CIN(\s$1539 ),
    .COUT(\c$2380 ),
    .SUM(\s$2381 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_68_0 (.A(\s$689 ),
    .B(\c$1530 ),
    .CIN(\c$1532 ),
    .COUT(\c$2382 ),
    .SUM(\s$2383 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_68_1 (.A(\c$1534 ),
    .B(\c$1536 ),
    .CIN(\c$1538 ),
    .COUT(\c$2384 ),
    .SUM(\s$2385 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_68_2 (.A(\c$1540 ),
    .B(\s$1543 ),
    .CIN(\s$1545 ),
    .COUT(\c$2386 ),
    .SUM(\s$2387 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_68_3 (.A(\s$1547 ),
    .B(\s$1549 ),
    .CIN(\s$1551 ),
    .COUT(\c$2388 ),
    .SUM(\s$2389 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_69_0 (.A(\s$707 ),
    .B(\c$1542 ),
    .CIN(\c$1544 ),
    .COUT(\c$2390 ),
    .SUM(\s$2391 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_69_1 (.A(\c$1546 ),
    .B(\c$1548 ),
    .CIN(\c$1550 ),
    .COUT(\c$2392 ),
    .SUM(\s$2393 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_69_2 (.A(\c$1552 ),
    .B(\s$1555 ),
    .CIN(\s$1557 ),
    .COUT(\c$2394 ),
    .SUM(\s$2395 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_69_3 (.A(\s$1559 ),
    .B(\s$1561 ),
    .CIN(\s$1563 ),
    .COUT(\c$2396 ),
    .SUM(\s$2397 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_70_0 (.A(\s$725 ),
    .B(\c$1554 ),
    .CIN(\c$1556 ),
    .COUT(\c$2398 ),
    .SUM(\s$2399 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_70_1 (.A(\c$1558 ),
    .B(\c$1560 ),
    .CIN(\c$1562 ),
    .COUT(\c$2400 ),
    .SUM(\s$2401 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_70_2 (.A(\c$1564 ),
    .B(\s$1567 ),
    .CIN(\s$1569 ),
    .COUT(\c$2402 ),
    .SUM(\s$2403 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_70_3 (.A(\s$1571 ),
    .B(\s$1573 ),
    .CIN(\s$1575 ),
    .COUT(\c$2404 ),
    .SUM(\s$2405 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_71_0 (.A(\s$743 ),
    .B(\c$1566 ),
    .CIN(\c$1568 ),
    .COUT(\c$2406 ),
    .SUM(\s$2407 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_71_1 (.A(\c$1570 ),
    .B(\c$1572 ),
    .CIN(\c$1574 ),
    .COUT(\c$2408 ),
    .SUM(\s$2409 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_71_2 (.A(\c$1576 ),
    .B(\s$1579 ),
    .CIN(\s$1581 ),
    .COUT(\c$2410 ),
    .SUM(\s$2411 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_71_3 (.A(\s$1583 ),
    .B(\s$1585 ),
    .CIN(\s$1587 ),
    .COUT(\c$2412 ),
    .SUM(\s$2413 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_72_0 (.A(\s$761 ),
    .B(\c$1578 ),
    .CIN(\c$1580 ),
    .COUT(\c$2414 ),
    .SUM(\s$2415 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_72_1 (.A(\c$1582 ),
    .B(\c$1584 ),
    .CIN(\c$1586 ),
    .COUT(\c$2416 ),
    .SUM(\s$2417 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_72_2 (.A(\c$1588 ),
    .B(\s$1591 ),
    .CIN(\s$1593 ),
    .COUT(\c$2418 ),
    .SUM(\s$2419 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_72_3 (.A(\s$1595 ),
    .B(\s$1597 ),
    .CIN(\s$1599 ),
    .COUT(\c$2420 ),
    .SUM(\s$2421 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_73_0 (.A(\s$779 ),
    .B(\c$1590 ),
    .CIN(\c$1592 ),
    .COUT(\c$2422 ),
    .SUM(\s$2423 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_73_1 (.A(\c$1594 ),
    .B(\c$1596 ),
    .CIN(\c$1598 ),
    .COUT(\c$2424 ),
    .SUM(\s$2425 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_73_2 (.A(\c$1600 ),
    .B(\s$1603 ),
    .CIN(\s$1605 ),
    .COUT(\c$2426 ),
    .SUM(\s$2427 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_73_3 (.A(\s$1607 ),
    .B(\s$1609 ),
    .CIN(\s$1611 ),
    .COUT(\c$2428 ),
    .SUM(\s$2429 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_74_0 (.A(\s$797 ),
    .B(\c$1602 ),
    .CIN(\c$1604 ),
    .COUT(\c$2430 ),
    .SUM(\s$2431 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_74_1 (.A(\c$1606 ),
    .B(\c$1608 ),
    .CIN(\c$1610 ),
    .COUT(\c$2432 ),
    .SUM(\s$2433 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_74_2 (.A(\c$1612 ),
    .B(\s$1615 ),
    .CIN(\s$1617 ),
    .COUT(\c$2434 ),
    .SUM(\s$2435 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_74_3 (.A(\s$1619 ),
    .B(\s$1621 ),
    .CIN(\s$1623 ),
    .COUT(\c$2436 ),
    .SUM(\s$2437 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_75_0 (.A(\s$815 ),
    .B(\c$1614 ),
    .CIN(\c$1616 ),
    .COUT(\c$2438 ),
    .SUM(\s$2439 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_75_1 (.A(\c$1618 ),
    .B(\c$1620 ),
    .CIN(\c$1622 ),
    .COUT(\c$2440 ),
    .SUM(\s$2441 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_75_2 (.A(\c$1624 ),
    .B(\s$1627 ),
    .CIN(\s$1629 ),
    .COUT(\c$2442 ),
    .SUM(\s$2443 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_75_3 (.A(\s$1631 ),
    .B(\s$1633 ),
    .CIN(\s$1635 ),
    .COUT(\c$2444 ),
    .SUM(\s$2445 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_76_0 (.A(\s$833 ),
    .B(\c$1626 ),
    .CIN(\c$1628 ),
    .COUT(\c$2446 ),
    .SUM(\s$2447 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_76_1 (.A(\c$1630 ),
    .B(\c$1632 ),
    .CIN(\c$1634 ),
    .COUT(\c$2448 ),
    .SUM(\s$2449 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_76_2 (.A(\c$1636 ),
    .B(\s$1639 ),
    .CIN(\s$1641 ),
    .COUT(\c$2450 ),
    .SUM(\s$2451 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_76_3 (.A(\s$1643 ),
    .B(\s$1645 ),
    .CIN(\s$1647 ),
    .COUT(\c$2452 ),
    .SUM(\s$2453 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_77_0 (.A(\s$851 ),
    .B(\c$1638 ),
    .CIN(\c$1640 ),
    .COUT(\c$2454 ),
    .SUM(\s$2455 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_77_1 (.A(\c$1642 ),
    .B(\c$1644 ),
    .CIN(\c$1646 ),
    .COUT(\c$2456 ),
    .SUM(\s$2457 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_77_2 (.A(\c$1648 ),
    .B(\s$1651 ),
    .CIN(\s$1653 ),
    .COUT(\c$2458 ),
    .SUM(\s$2459 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_77_3 (.A(\s$1655 ),
    .B(\s$1657 ),
    .CIN(\s$1659 ),
    .COUT(\c$2460 ),
    .SUM(\s$2461 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_78_0 (.A(\s$869 ),
    .B(\c$1650 ),
    .CIN(\c$1652 ),
    .COUT(\c$2462 ),
    .SUM(\s$2463 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_78_1 (.A(\c$1654 ),
    .B(\c$1656 ),
    .CIN(\c$1658 ),
    .COUT(\c$2464 ),
    .SUM(\s$2465 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_78_2 (.A(\c$1660 ),
    .B(\s$1663 ),
    .CIN(\s$1665 ),
    .COUT(\c$2466 ),
    .SUM(\s$2467 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_78_3 (.A(\s$1667 ),
    .B(\s$1669 ),
    .CIN(\s$1671 ),
    .COUT(\c$2468 ),
    .SUM(\s$2469 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_79_0 (.A(\s$887 ),
    .B(\c$1662 ),
    .CIN(\c$1664 ),
    .COUT(\c$2470 ),
    .SUM(\s$2471 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_79_1 (.A(\c$1666 ),
    .B(\c$1668 ),
    .CIN(\c$1670 ),
    .COUT(\c$2472 ),
    .SUM(\s$2473 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_79_2 (.A(\c$1672 ),
    .B(\s$1675 ),
    .CIN(\s$1677 ),
    .COUT(\c$2474 ),
    .SUM(\s$2475 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_79_3 (.A(\s$1679 ),
    .B(\s$1681 ),
    .CIN(\s$1683 ),
    .COUT(\c$2476 ),
    .SUM(\s$2477 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_80_0 (.A(\s$905 ),
    .B(\c$1674 ),
    .CIN(\c$1676 ),
    .COUT(\c$2478 ),
    .SUM(\s$2479 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_80_1 (.A(\c$1678 ),
    .B(\c$1680 ),
    .CIN(\c$1682 ),
    .COUT(\c$2480 ),
    .SUM(\s$2481 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_80_2 (.A(\c$1684 ),
    .B(\s$1687 ),
    .CIN(\s$1689 ),
    .COUT(\c$2482 ),
    .SUM(\s$2483 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_80_3 (.A(\s$1691 ),
    .B(\s$1693 ),
    .CIN(\s$1695 ),
    .COUT(\c$2484 ),
    .SUM(\s$2485 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_81_0 (.A(\s$921 ),
    .B(\c$1686 ),
    .CIN(\c$1688 ),
    .COUT(\c$2486 ),
    .SUM(\s$2487 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_81_1 (.A(\c$1690 ),
    .B(\c$1692 ),
    .CIN(\c$1694 ),
    .COUT(\c$2488 ),
    .SUM(\s$2489 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_81_2 (.A(\c$1696 ),
    .B(\s$1699 ),
    .CIN(\s$1701 ),
    .COUT(\c$2490 ),
    .SUM(\s$2491 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_81_3 (.A(\s$1703 ),
    .B(\s$1705 ),
    .CIN(\s$1707 ),
    .COUT(\c$2492 ),
    .SUM(\s$2493 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_82_0 (.A(\s$937 ),
    .B(\c$1698 ),
    .CIN(\c$1700 ),
    .COUT(\c$2494 ),
    .SUM(\s$2495 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_82_1 (.A(\c$1702 ),
    .B(\c$1704 ),
    .CIN(\c$1706 ),
    .COUT(\c$2496 ),
    .SUM(\s$2497 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_82_2 (.A(\c$1708 ),
    .B(\s$1711 ),
    .CIN(\s$1713 ),
    .COUT(\c$2498 ),
    .SUM(\s$2499 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_82_3 (.A(\s$1715 ),
    .B(\s$1717 ),
    .CIN(\s$1719 ),
    .COUT(\c$2500 ),
    .SUM(\s$2501 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_83_0 (.A(\s$951 ),
    .B(\c$1710 ),
    .CIN(\c$1712 ),
    .COUT(\c$2502 ),
    .SUM(\s$2503 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_83_1 (.A(\c$1714 ),
    .B(\c$1716 ),
    .CIN(\c$1718 ),
    .COUT(\c$2504 ),
    .SUM(\s$2505 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_83_2 (.A(\c$1720 ),
    .B(\s$1723 ),
    .CIN(\s$1725 ),
    .COUT(\c$2506 ),
    .SUM(\s$2507 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_83_3 (.A(\s$1727 ),
    .B(\s$1729 ),
    .CIN(\s$1731 ),
    .COUT(\c$2508 ),
    .SUM(\s$2509 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_84_0 (.A(\s$965 ),
    .B(\c$1722 ),
    .CIN(\c$1724 ),
    .COUT(\c$2510 ),
    .SUM(\s$2511 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_84_1 (.A(\c$1726 ),
    .B(\c$1728 ),
    .CIN(\c$1730 ),
    .COUT(\c$2512 ),
    .SUM(\s$2513 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_84_2 (.A(\c$1732 ),
    .B(\s$1735 ),
    .CIN(\s$1737 ),
    .COUT(\c$2514 ),
    .SUM(\s$2515 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_84_3 (.A(\s$1739 ),
    .B(\s$1741 ),
    .CIN(\s$1743 ),
    .COUT(\c$2516 ),
    .SUM(\s$2517 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_85_0 (.A(\s$977 ),
    .B(\c$1734 ),
    .CIN(\c$1736 ),
    .COUT(\c$2518 ),
    .SUM(\s$2519 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_85_1 (.A(\c$1738 ),
    .B(\c$1740 ),
    .CIN(\c$1742 ),
    .COUT(\c$2520 ),
    .SUM(\s$2521 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_85_2 (.A(\c$1744 ),
    .B(\s$1747 ),
    .CIN(\s$1749 ),
    .COUT(\c$2522 ),
    .SUM(\s$2523 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_85_3 (.A(\s$1751 ),
    .B(\s$1753 ),
    .CIN(\s$1755 ),
    .COUT(\c$2524 ),
    .SUM(\s$2525 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_86_0 (.A(\s$989 ),
    .B(\c$1746 ),
    .CIN(\c$1748 ),
    .COUT(\c$2526 ),
    .SUM(\s$2527 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_86_1 (.A(\c$1750 ),
    .B(\c$1752 ),
    .CIN(\c$1754 ),
    .COUT(\c$2528 ),
    .SUM(\s$2529 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_86_2 (.A(\c$1756 ),
    .B(\s$1759 ),
    .CIN(\s$1761 ),
    .COUT(\c$2530 ),
    .SUM(\s$2531 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_86_3 (.A(\s$1763 ),
    .B(\s$1765 ),
    .CIN(\s$1767 ),
    .COUT(\c$2532 ),
    .SUM(\s$2533 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_87_0 (.A(\s$999 ),
    .B(\c$1758 ),
    .CIN(\c$1760 ),
    .COUT(\c$2534 ),
    .SUM(\s$2535 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_87_1 (.A(\c$1762 ),
    .B(\c$1764 ),
    .CIN(\c$1766 ),
    .COUT(\c$2536 ),
    .SUM(\s$2537 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_87_2 (.A(\c$1768 ),
    .B(\s$1771 ),
    .CIN(\s$1773 ),
    .COUT(\c$2538 ),
    .SUM(\s$2539 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_87_3 (.A(\s$1775 ),
    .B(\s$1777 ),
    .CIN(\s$1779 ),
    .COUT(\c$2540 ),
    .SUM(\s$2541 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_88_0 (.A(\s$1009 ),
    .B(\c$1770 ),
    .CIN(\c$1772 ),
    .COUT(\c$2542 ),
    .SUM(\s$2543 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_88_1 (.A(\c$1774 ),
    .B(\c$1776 ),
    .CIN(\c$1778 ),
    .COUT(\c$2544 ),
    .SUM(\s$2545 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_88_2 (.A(\c$1780 ),
    .B(\s$1783 ),
    .CIN(\s$1785 ),
    .COUT(\c$2546 ),
    .SUM(\s$2547 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_88_3 (.A(\s$1787 ),
    .B(\s$1789 ),
    .CIN(\s$1791 ),
    .COUT(\c$2548 ),
    .SUM(\s$2549 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_89_0 (.A(\s$1017 ),
    .B(\c$1782 ),
    .CIN(\c$1784 ),
    .COUT(\c$2550 ),
    .SUM(\s$2551 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_89_1 (.A(\c$1786 ),
    .B(\c$1788 ),
    .CIN(\c$1790 ),
    .COUT(\c$2552 ),
    .SUM(\s$2553 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_89_2 (.A(\c$1792 ),
    .B(\s$1795 ),
    .CIN(\s$1797 ),
    .COUT(\c$2554 ),
    .SUM(\s$2555 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_89_3 (.A(\s$1799 ),
    .B(\s$1801 ),
    .CIN(\s$1803 ),
    .COUT(\c$2556 ),
    .SUM(\s$2557 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_90_0 (.A(\s$1025 ),
    .B(\c$1794 ),
    .CIN(\c$1796 ),
    .COUT(\c$2558 ),
    .SUM(\s$2559 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_90_1 (.A(\c$1798 ),
    .B(\c$1800 ),
    .CIN(\c$1802 ),
    .COUT(\c$2560 ),
    .SUM(\s$2561 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_90_2 (.A(\c$1804 ),
    .B(\s$1807 ),
    .CIN(\s$1809 ),
    .COUT(\c$2562 ),
    .SUM(\s$2563 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_90_3 (.A(\s$1811 ),
    .B(\s$1813 ),
    .CIN(\s$1815 ),
    .COUT(\c$2564 ),
    .SUM(\s$2565 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_91_0 (.A(\s$1031 ),
    .B(\c$1806 ),
    .CIN(\c$1808 ),
    .COUT(\c$2566 ),
    .SUM(\s$2567 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_91_1 (.A(\c$1810 ),
    .B(\c$1812 ),
    .CIN(\c$1814 ),
    .COUT(\c$2568 ),
    .SUM(\s$2569 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_91_2 (.A(\c$1816 ),
    .B(\s$1819 ),
    .CIN(\s$1821 ),
    .COUT(\c$2570 ),
    .SUM(\s$2571 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_91_3 (.A(\s$1823 ),
    .B(\s$1825 ),
    .CIN(\s$1827 ),
    .COUT(\c$2572 ),
    .SUM(\s$2573 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_92_0 (.A(\s$1037 ),
    .B(\c$1818 ),
    .CIN(\c$1820 ),
    .COUT(\c$2574 ),
    .SUM(\s$2575 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_92_1 (.A(\c$1822 ),
    .B(\c$1824 ),
    .CIN(\c$1826 ),
    .COUT(\c$2576 ),
    .SUM(\s$2577 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_92_2 (.A(\c$1828 ),
    .B(\s$1831 ),
    .CIN(\s$1833 ),
    .COUT(\c$2578 ),
    .SUM(\s$2579 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_92_3 (.A(\s$1835 ),
    .B(\s$1837 ),
    .CIN(\s$1839 ),
    .COUT(\c$2580 ),
    .SUM(\s$2581 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_93_0 (.A(\s$1041 ),
    .B(\c$1830 ),
    .CIN(\c$1832 ),
    .COUT(\c$2582 ),
    .SUM(\s$2583 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_93_1 (.A(\c$1834 ),
    .B(\c$1836 ),
    .CIN(\c$1838 ),
    .COUT(\c$2584 ),
    .SUM(\s$2585 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_93_2 (.A(\c$1840 ),
    .B(\s$1843 ),
    .CIN(\s$1845 ),
    .COUT(\c$2586 ),
    .SUM(\s$2587 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_93_3 (.A(\s$1847 ),
    .B(\s$1849 ),
    .CIN(\s$1851 ),
    .COUT(\c$2588 ),
    .SUM(\s$2589 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_94_0 (.A(\s$1045 ),
    .B(\c$1842 ),
    .CIN(\c$1844 ),
    .COUT(\c$2590 ),
    .SUM(\s$2591 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_94_1 (.A(\c$1846 ),
    .B(\c$1848 ),
    .CIN(\c$1850 ),
    .COUT(\c$2592 ),
    .SUM(\s$2593 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_94_2 (.A(\c$1852 ),
    .B(\s$1855 ),
    .CIN(\s$1857 ),
    .COUT(\c$2594 ),
    .SUM(\s$2595 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_94_3 (.A(\s$1859 ),
    .B(\s$1861 ),
    .CIN(\s$1863 ),
    .COUT(\c$2596 ),
    .SUM(\s$2597 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_95_0 (.A(\s$1047 ),
    .B(\c$1854 ),
    .CIN(\c$1856 ),
    .COUT(\c$2598 ),
    .SUM(\s$2599 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_3_95_1 (.A(\c$1858 ),
    .B(\c$1860 ),
    .CIN(\c$1862 ),
    .COUT(\c$2600 ),
    .SUM(\s$2601 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_95_2 (.A(\c$1864 ),
    .B(\s$1867 ),
    .CIN(\s$1869 ),
    .COUT(\c$2602 ),
    .SUM(\s$2603 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_95_3 (.A(\s$1871 ),
    .B(\s$1873 ),
    .CIN(\s$1875 ),
    .COUT(\c$2604 ),
    .SUM(\s$2605 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_96_0 (.A(\s$1049 ),
    .B(\c$1866 ),
    .CIN(\c$1868 ),
    .COUT(\c$2606 ),
    .SUM(\s$2607 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_96_1 (.A(\c$1870 ),
    .B(\c$1872 ),
    .CIN(\c$1874 ),
    .COUT(\c$2608 ),
    .SUM(\s$2609 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_96_2 (.A(\c$1876 ),
    .B(\s$1879 ),
    .CIN(\s$1881 ),
    .COUT(\c$2610 ),
    .SUM(\s$2611 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_96_3 (.A(\s$1883 ),
    .B(\s$1885 ),
    .CIN(\s$1887 ),
    .COUT(\c$2612 ),
    .SUM(\s$2613 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_97_0 (.A(\c$1048 ),
    .B(\c$1878 ),
    .CIN(\c$1880 ),
    .COUT(\c$2614 ),
    .SUM(\s$2615 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_97_1 (.A(\c$1882 ),
    .B(\c$1884 ),
    .CIN(\c$1886 ),
    .COUT(\c$2616 ),
    .SUM(\s$2617 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_97_2 (.A(\c$1888 ),
    .B(\s$1891 ),
    .CIN(\s$1893 ),
    .COUT(\c$2618 ),
    .SUM(\s$2619 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_97_3 (.A(\s$1895 ),
    .B(\s$1897 ),
    .CIN(\s$1899 ),
    .COUT(\c$2620 ),
    .SUM(\s$2621 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_98_0 (.A(pp_row98_17),
    .B(\c$1890 ),
    .CIN(\c$1892 ),
    .COUT(\c$2622 ),
    .SUM(\s$2623 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_98_1 (.A(\c$1894 ),
    .B(\c$1896 ),
    .CIN(\c$1898 ),
    .COUT(\c$2624 ),
    .SUM(\s$2625 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_98_2 (.A(\c$1900 ),
    .B(\s$1903 ),
    .CIN(\s$1905 ),
    .COUT(\c$2626 ),
    .SUM(\s$2627 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_98_3 (.A(\s$1907 ),
    .B(\s$1909 ),
    .CIN(\s$1911 ),
    .COUT(\c$2628 ),
    .SUM(\s$2629 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_99_0 (.A(pp_row99_15),
    .B(pp_row99_16),
    .CIN(\c$1902 ),
    .COUT(\c$2630 ),
    .SUM(\s$2631 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_99_1 (.A(\c$1904 ),
    .B(\c$1906 ),
    .CIN(\c$1908 ),
    .COUT(\c$2632 ),
    .SUM(\s$2633 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_99_2 (.A(\c$1910 ),
    .B(\c$1912 ),
    .CIN(\s$1915 ),
    .COUT(\c$2634 ),
    .SUM(\s$2635 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_3_99_3 (.A(\s$1917 ),
    .B(\s$1919 ),
    .CIN(\s$1921 ),
    .COUT(\c$2636 ),
    .SUM(\s$2637 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_100_0 (.A(\s$1933 ),
    .B(\c$2630 ),
    .CIN(\c$2632 ),
    .COUT(\c$3290 ),
    .SUM(\s$3291 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_100_1 (.A(\c$2634 ),
    .B(\c$2636 ),
    .CIN(\s$2639 ),
    .COUT(\c$3292 ),
    .SUM(\s$3293 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_100_2 (.A(\s$2641 ),
    .B(\s$2643 ),
    .CIN(\s$2645 ),
    .COUT(\c$3294 ),
    .SUM(\s$3295 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_101_0 (.A(\s$1941 ),
    .B(\c$2638 ),
    .CIN(\c$2640 ),
    .COUT(\c$3296 ),
    .SUM(\s$3297 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_101_1 (.A(\c$2642 ),
    .B(\c$2644 ),
    .CIN(\s$2647 ),
    .COUT(\c$3298 ),
    .SUM(\s$3299 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_101_2 (.A(\s$2649 ),
    .B(\s$2651 ),
    .CIN(\s$2653 ),
    .COUT(\c$3300 ),
    .SUM(\s$3301 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_102_0 (.A(\s$1949 ),
    .B(\c$2646 ),
    .CIN(\c$2648 ),
    .COUT(\c$3302 ),
    .SUM(\s$3303 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_102_1 (.A(\c$2650 ),
    .B(\c$2652 ),
    .CIN(\s$2655 ),
    .COUT(\c$3304 ),
    .SUM(\s$3305 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_102_2 (.A(\s$2657 ),
    .B(\s$2659 ),
    .CIN(\s$2661 ),
    .COUT(\c$3306 ),
    .SUM(\s$3307 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_103_0 (.A(\s$1955 ),
    .B(\c$2654 ),
    .CIN(\c$2656 ),
    .COUT(\c$3308 ),
    .SUM(\s$3309 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_103_1 (.A(\c$2658 ),
    .B(\c$2660 ),
    .CIN(\s$2663 ),
    .COUT(\c$3310 ),
    .SUM(\s$3311 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_103_2 (.A(\s$2665 ),
    .B(\s$2667 ),
    .CIN(\s$2669 ),
    .COUT(\c$3312 ),
    .SUM(\s$3313 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_104_0 (.A(\s$1961 ),
    .B(\c$2662 ),
    .CIN(\c$2664 ),
    .COUT(\c$3314 ),
    .SUM(\s$3315 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_104_1 (.A(\c$2666 ),
    .B(\c$2668 ),
    .CIN(\s$2671 ),
    .COUT(\c$3316 ),
    .SUM(\s$3317 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_104_2 (.A(\s$2673 ),
    .B(\s$2675 ),
    .CIN(\s$2677 ),
    .COUT(\c$3318 ),
    .SUM(\s$3319 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_105_0 (.A(\s$1965 ),
    .B(\c$2670 ),
    .CIN(\c$2672 ),
    .COUT(\c$3320 ),
    .SUM(\s$3321 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_105_1 (.A(\c$2674 ),
    .B(\c$2676 ),
    .CIN(\s$2679 ),
    .COUT(\c$3322 ),
    .SUM(\s$3323 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_105_2 (.A(\s$2681 ),
    .B(\s$2683 ),
    .CIN(\s$2685 ),
    .COUT(\c$3324 ),
    .SUM(\s$3325 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_106_0 (.A(\s$1969 ),
    .B(\c$2678 ),
    .CIN(\c$2680 ),
    .COUT(\c$3326 ),
    .SUM(\s$3327 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_106_1 (.A(\c$2682 ),
    .B(\c$2684 ),
    .CIN(\s$2687 ),
    .COUT(\c$3328 ),
    .SUM(\s$3329 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_106_2 (.A(\s$2689 ),
    .B(\s$2691 ),
    .CIN(\s$2693 ),
    .COUT(\c$3330 ),
    .SUM(\s$3331 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_107_0 (.A(\s$1971 ),
    .B(\c$2686 ),
    .CIN(\c$2688 ),
    .COUT(\c$3332 ),
    .SUM(\s$3333 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_107_1 (.A(\c$2690 ),
    .B(\c$2692 ),
    .CIN(\s$2695 ),
    .COUT(\c$3334 ),
    .SUM(\s$3335 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_107_2 (.A(\s$2697 ),
    .B(\s$2699 ),
    .CIN(\s$2701 ),
    .COUT(\c$3336 ),
    .SUM(\s$3337 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_108_0 (.A(\s$1973 ),
    .B(\c$2694 ),
    .CIN(\c$2696 ),
    .COUT(\c$3338 ),
    .SUM(\s$3339 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_108_1 (.A(\c$2698 ),
    .B(\c$2700 ),
    .CIN(\s$2703 ),
    .COUT(\c$3340 ),
    .SUM(\s$3341 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_108_2 (.A(\s$2705 ),
    .B(\s$2707 ),
    .CIN(\s$2709 ),
    .COUT(\c$3342 ),
    .SUM(\s$3343 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_109_0 (.A(\c$1972 ),
    .B(\c$2702 ),
    .CIN(\c$2704 ),
    .COUT(\c$3344 ),
    .SUM(\s$3345 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_109_1 (.A(\c$2706 ),
    .B(\c$2708 ),
    .CIN(\s$2711 ),
    .COUT(\c$3346 ),
    .SUM(\s$3347 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_109_2 (.A(\s$2713 ),
    .B(\s$2715 ),
    .CIN(\s$2717 ),
    .COUT(\c$3348 ),
    .SUM(\s$3349 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_10_0 (.A(pp_row10_0),
    .B(pp_row10_1),
    .CIN(pp_row10_2),
    .COUT(\c$2754 ),
    .SUM(\s$2755 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_110_0 (.A(pp_row110_11),
    .B(\c$2710 ),
    .CIN(\c$2712 ),
    .COUT(\c$3350 ),
    .SUM(\s$3351 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_110_1 (.A(\c$2714 ),
    .B(\c$2716 ),
    .CIN(\s$2719 ),
    .COUT(\c$3352 ),
    .SUM(\s$3353 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_110_2 (.A(\s$2721 ),
    .B(\s$2723 ),
    .CIN(\s$2725 ),
    .COUT(\c$3354 ),
    .SUM(\s$3355 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_111_0 (.A(pp_row111_9),
    .B(pp_row111_10),
    .CIN(\c$2718 ),
    .COUT(\c$3356 ),
    .SUM(\s$3357 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_111_1 (.A(\c$2720 ),
    .B(\c$2722 ),
    .CIN(\c$2724 ),
    .COUT(\c$3358 ),
    .SUM(\s$3359 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_111_2 (.A(\s$2727 ),
    .B(\s$2729 ),
    .CIN(\s$2731 ),
    .COUT(\c$3360 ),
    .SUM(\s$3361 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_4_112_0 (.A(pp_row112_8),
    .B(pp_row112_9),
    .CIN(pp_row112_10),
    .COUT(\c$3362 ),
    .SUM(\s$3363 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_112_1 (.A(\c$2726 ),
    .B(\c$2728 ),
    .CIN(\c$2730 ),
    .COUT(\c$3364 ),
    .SUM(\s$3365 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_112_2 (.A(\s$2733 ),
    .B(\s$2735 ),
    .CIN(\s$2737 ),
    .COUT(\c$3366 ),
    .SUM(\s$3367 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_113_0 (.A(pp_row113_6),
    .B(pp_row113_7),
    .CIN(pp_row113_8),
    .COUT(\c$3368 ),
    .SUM(\s$3369 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_113_1 (.A(pp_row113_9),
    .B(\c$2732 ),
    .CIN(\c$2734 ),
    .COUT(\c$3370 ),
    .SUM(\s$3371 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_113_2 (.A(\c$2736 ),
    .B(\s$2739 ),
    .CIN(\s$2741 ),
    .COUT(\c$3372 ),
    .SUM(\s$3373 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_114_0 (.A(pp_row114_5),
    .B(pp_row114_6),
    .CIN(pp_row114_7),
    .COUT(\c$3374 ),
    .SUM(\s$3375 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_114_1 (.A(pp_row114_8),
    .B(pp_row114_9),
    .CIN(\c$2738 ),
    .COUT(\c$3376 ),
    .SUM(\s$3377 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_114_2 (.A(\c$2740 ),
    .B(\s$2743 ),
    .CIN(\s$2745 ),
    .COUT(\c$3378 ),
    .SUM(\s$3379 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_4_115_0 (.A(pp_row115_3),
    .B(pp_row115_4),
    .CIN(pp_row115_5),
    .COUT(\c$3380 ),
    .SUM(\s$3381 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_115_1 (.A(pp_row115_6),
    .B(pp_row115_7),
    .CIN(pp_row115_8),
    .COUT(\c$3382 ),
    .SUM(\s$3383 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_115_2 (.A(\c$2742 ),
    .B(\c$2744 ),
    .CIN(\s$2747 ),
    .COUT(\c$3384 ),
    .SUM(\s$3385 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_116_0 (.A(pp_row116_2),
    .B(pp_row116_3),
    .CIN(pp_row116_4),
    .COUT(\c$3386 ),
    .SUM(\s$3387 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_116_1 (.A(pp_row116_5),
    .B(pp_row116_6),
    .CIN(pp_row116_7),
    .COUT(\c$3388 ),
    .SUM(\s$3389 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_4_116_2 (.A(pp_row116_8),
    .B(\c$2746 ),
    .CIN(\s$2749 ),
    .COUT(\c$3390 ),
    .SUM(\s$3391 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_117_0 (.A(pp_row117_0),
    .B(pp_row117_1),
    .CIN(pp_row117_2),
    .COUT(\c$3392 ),
    .SUM(\s$3393 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_117_1 (.A(pp_row117_3),
    .B(pp_row117_4),
    .CIN(pp_row117_5),
    .COUT(\c$3394 ),
    .SUM(\s$3395 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_117_2 (.A(pp_row117_6),
    .B(pp_row117_7),
    .CIN(\c$2748 ),
    .COUT(\c$3396 ),
    .SUM(\s$3397 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_118_0 (.A(net1912),
    .B(pp_row118_1),
    .CIN(pp_row118_2),
    .COUT(\c$3398 ),
    .SUM(\s$3399 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_118_1 (.A(pp_row118_3),
    .B(pp_row118_4),
    .CIN(pp_row118_5),
    .COUT(\c$3400 ),
    .SUM(\s$3401 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_119_0 (.A(pp_row119_0),
    .B(pp_row119_1),
    .CIN(pp_row119_2),
    .COUT(\c$3404 ),
    .SUM(\s$3405 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_119_1 (.A(pp_row119_3),
    .B(pp_row119_4),
    .CIN(pp_row119_5),
    .COUT(\c$3406 ),
    .SUM(\s$3407 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_11_0 (.A(pp_row11_0),
    .B(pp_row11_1),
    .CIN(pp_row11_2),
    .COUT(\c$2758 ),
    .SUM(\s$2759 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_120_0 (.A(net1913),
    .B(pp_row120_1),
    .CIN(pp_row120_2),
    .COUT(\c$3408 ),
    .SUM(\s$3409 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_121_0 (.A(pp_row121_0),
    .B(pp_row121_1),
    .CIN(pp_row121_2),
    .COUT(\c$3412 ),
    .SUM(\s$3413 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_12_0 (.A(pp_row12_0),
    .B(pp_row12_1),
    .CIN(pp_row12_2),
    .COUT(\c$2762 ),
    .SUM(\s$2763 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_12_1 (.A(pp_row12_3),
    .B(pp_row12_4),
    .CIN(pp_row12_5),
    .COUT(\c$2764 ),
    .SUM(\s$2765 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_13_0 (.A(pp_row13_0),
    .B(pp_row13_1),
    .CIN(pp_row13_2),
    .COUT(\c$2768 ),
    .SUM(\s$2769 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_13_1 (.A(pp_row13_3),
    .B(pp_row13_4),
    .CIN(pp_row13_5),
    .COUT(\c$2770 ),
    .SUM(\s$2771 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_14_0 (.A(pp_row14_2),
    .B(pp_row14_3),
    .CIN(pp_row14_4),
    .COUT(\c$2774 ),
    .SUM(\s$2775 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_14_1 (.A(pp_row14_5),
    .B(pp_row14_6),
    .CIN(pp_row14_7),
    .COUT(\c$2776 ),
    .SUM(\s$2777 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_14_2 (.A(pp_row14_8),
    .B(pp_row14_9),
    .CIN(\s$1975 ),
    .COUT(\c$2778 ),
    .SUM(\s$2779 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_15_0 (.A(pp_row15_2),
    .B(pp_row15_3),
    .CIN(pp_row15_4),
    .COUT(\c$2780 ),
    .SUM(\s$2781 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_15_1 (.A(pp_row15_5),
    .B(pp_row15_6),
    .CIN(pp_row15_7),
    .COUT(\c$2782 ),
    .SUM(\s$2783 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_15_2 (.A(pp_row15_8),
    .B(\c$1974 ),
    .CIN(\s$1977 ),
    .COUT(\c$2784 ),
    .SUM(\s$2785 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_16_0 (.A(pp_row16_5),
    .B(pp_row16_6),
    .CIN(pp_row16_7),
    .COUT(\c$2786 ),
    .SUM(\s$2787 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_16_1 (.A(pp_row16_8),
    .B(pp_row16_9),
    .CIN(pp_row16_10),
    .COUT(\c$2788 ),
    .SUM(\s$2789 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_16_2 (.A(\c$1976 ),
    .B(\s$1979 ),
    .CIN(\s$1981 ),
    .COUT(\c$2790 ),
    .SUM(\s$2791 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_17_0 (.A(pp_row17_5),
    .B(pp_row17_6),
    .CIN(pp_row17_7),
    .COUT(\c$2792 ),
    .SUM(\s$2793 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_17_1 (.A(pp_row17_8),
    .B(pp_row17_9),
    .CIN(\c$1978 ),
    .COUT(\c$2794 ),
    .SUM(\s$2795 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_17_2 (.A(\c$1980 ),
    .B(\s$1983 ),
    .CIN(\s$1985 ),
    .COUT(\c$2796 ),
    .SUM(\s$2797 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_18_0 (.A(pp_row18_8),
    .B(pp_row18_9),
    .CIN(pp_row18_10),
    .COUT(\c$2798 ),
    .SUM(\s$2799 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_18_1 (.A(pp_row18_11),
    .B(\c$1982 ),
    .CIN(\c$1984 ),
    .COUT(\c$2800 ),
    .SUM(\s$2801 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_18_2 (.A(\s$1987 ),
    .B(\s$1989 ),
    .CIN(\s$1991 ),
    .COUT(\c$2802 ),
    .SUM(\s$2803 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_19_0 (.A(pp_row19_8),
    .B(pp_row19_9),
    .CIN(pp_row19_10),
    .COUT(\c$2804 ),
    .SUM(\s$2805 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_19_1 (.A(\c$1986 ),
    .B(\c$1988 ),
    .CIN(\c$1990 ),
    .COUT(\c$2806 ),
    .SUM(\s$2807 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_19_2 (.A(\s$1993 ),
    .B(\s$1995 ),
    .CIN(\s$1997 ),
    .COUT(\c$2808 ),
    .SUM(\s$2809 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_20_0 (.A(pp_row20_11),
    .B(pp_row20_12),
    .CIN(\c$1992 ),
    .COUT(\c$2810 ),
    .SUM(\s$2811 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_20_1 (.A(\c$1994 ),
    .B(\c$1996 ),
    .CIN(\s$1999 ),
    .COUT(\c$2812 ),
    .SUM(\s$2813 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_20_2 (.A(\s$2001 ),
    .B(\s$2003 ),
    .CIN(\s$2005 ),
    .COUT(\c$2814 ),
    .SUM(\s$2815 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_21_0 (.A(pp_row21_11),
    .B(\c$1998 ),
    .CIN(\c$2000 ),
    .COUT(\c$2816 ),
    .SUM(\s$2817 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_21_1 (.A(\c$2002 ),
    .B(\c$2004 ),
    .CIN(\s$2007 ),
    .COUT(\c$2818 ),
    .SUM(\s$2819 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_21_2 (.A(\s$2009 ),
    .B(\s$2011 ),
    .CIN(\s$2013 ),
    .COUT(\c$2820 ),
    .SUM(\s$2821 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_22_0 (.A(\s$1051 ),
    .B(\c$2006 ),
    .CIN(\c$2008 ),
    .COUT(\c$2822 ),
    .SUM(\s$2823 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_22_1 (.A(\c$2010 ),
    .B(\c$2012 ),
    .CIN(\s$2015 ),
    .COUT(\c$2824 ),
    .SUM(\s$2825 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_22_2 (.A(\s$2017 ),
    .B(\s$2019 ),
    .CIN(\s$2021 ),
    .COUT(\c$2826 ),
    .SUM(\s$2827 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_23_0 (.A(\s$1053 ),
    .B(\c$2014 ),
    .CIN(\c$2016 ),
    .COUT(\c$2828 ),
    .SUM(\s$2829 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_23_1 (.A(\c$2018 ),
    .B(\c$2020 ),
    .CIN(\s$2023 ),
    .COUT(\c$2830 ),
    .SUM(\s$2831 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_23_2 (.A(\s$2025 ),
    .B(\s$2027 ),
    .CIN(\s$2029 ),
    .COUT(\c$2832 ),
    .SUM(\s$2833 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_24_0 (.A(\s$1057 ),
    .B(\c$2022 ),
    .CIN(\c$2024 ),
    .COUT(\c$2834 ),
    .SUM(\s$2835 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_24_1 (.A(\c$2026 ),
    .B(\c$2028 ),
    .CIN(\s$2031 ),
    .COUT(\c$2836 ),
    .SUM(\s$2837 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_24_2 (.A(\s$2033 ),
    .B(\s$2035 ),
    .CIN(\s$2037 ),
    .COUT(\c$2838 ),
    .SUM(\s$2839 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_25_0 (.A(\s$1061 ),
    .B(\c$2030 ),
    .CIN(\c$2032 ),
    .COUT(\c$2840 ),
    .SUM(\s$2841 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_25_1 (.A(\c$2034 ),
    .B(\c$2036 ),
    .CIN(\s$2039 ),
    .COUT(\c$2842 ),
    .SUM(\s$2843 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_25_2 (.A(\s$2041 ),
    .B(\s$2043 ),
    .CIN(\s$2045 ),
    .COUT(\c$2844 ),
    .SUM(\s$2845 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_26_0 (.A(\s$1067 ),
    .B(\c$2038 ),
    .CIN(\c$2040 ),
    .COUT(\c$2846 ),
    .SUM(\s$2847 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_26_1 (.A(\c$2042 ),
    .B(\c$2044 ),
    .CIN(\s$2047 ),
    .COUT(\c$2848 ),
    .SUM(\s$2849 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_26_2 (.A(\s$2049 ),
    .B(\s$2051 ),
    .CIN(\s$2053 ),
    .COUT(\c$2850 ),
    .SUM(\s$2851 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_27_0 (.A(\s$1073 ),
    .B(\c$2046 ),
    .CIN(\c$2048 ),
    .COUT(\c$2852 ),
    .SUM(\s$2853 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_27_1 (.A(\c$2050 ),
    .B(\c$2052 ),
    .CIN(\s$2055 ),
    .COUT(\c$2854 ),
    .SUM(\s$2855 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_27_2 (.A(\s$2057 ),
    .B(\s$2059 ),
    .CIN(\s$2061 ),
    .COUT(\c$2856 ),
    .SUM(\s$2857 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_28_0 (.A(\s$1081 ),
    .B(\c$2054 ),
    .CIN(\c$2056 ),
    .COUT(\c$2858 ),
    .SUM(\s$2859 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_28_1 (.A(\c$2058 ),
    .B(\c$2060 ),
    .CIN(\s$2063 ),
    .COUT(\c$2860 ),
    .SUM(\s$2861 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_28_2 (.A(\s$2065 ),
    .B(\s$2067 ),
    .CIN(\s$2069 ),
    .COUT(\c$2862 ),
    .SUM(\s$2863 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_29_0 (.A(\s$1089 ),
    .B(\c$2062 ),
    .CIN(\c$2064 ),
    .COUT(\c$2864 ),
    .SUM(\s$2865 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_29_1 (.A(\c$2066 ),
    .B(\c$2068 ),
    .CIN(\s$2071 ),
    .COUT(\c$2866 ),
    .SUM(\s$2867 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_29_2 (.A(\s$2073 ),
    .B(\s$2075 ),
    .CIN(\s$2077 ),
    .COUT(\c$2868 ),
    .SUM(\s$2869 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_30_0 (.A(\s$1099 ),
    .B(\c$2070 ),
    .CIN(\c$2072 ),
    .COUT(\c$2870 ),
    .SUM(\s$2871 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_30_1 (.A(\c$2074 ),
    .B(\c$2076 ),
    .CIN(\s$2079 ),
    .COUT(\c$2872 ),
    .SUM(\s$2873 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_30_2 (.A(\s$2081 ),
    .B(\s$2083 ),
    .CIN(\s$2085 ),
    .COUT(\c$2874 ),
    .SUM(\s$2875 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_31_0 (.A(\s$1109 ),
    .B(\c$2078 ),
    .CIN(\c$2080 ),
    .COUT(\c$2876 ),
    .SUM(\s$2877 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_31_1 (.A(\c$2082 ),
    .B(\c$2084 ),
    .CIN(\s$2087 ),
    .COUT(\c$2878 ),
    .SUM(\s$2879 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_31_2 (.A(\s$2089 ),
    .B(\s$2091 ),
    .CIN(\s$2093 ),
    .COUT(\c$2880 ),
    .SUM(\s$2881 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_32_0 (.A(\s$1121 ),
    .B(\c$2086 ),
    .CIN(\c$2088 ),
    .COUT(\c$2882 ),
    .SUM(\s$2883 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_32_1 (.A(\c$2090 ),
    .B(\c$2092 ),
    .CIN(\s$2095 ),
    .COUT(\c$2884 ),
    .SUM(\s$2885 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_32_2 (.A(\s$2097 ),
    .B(\s$2099 ),
    .CIN(\s$2101 ),
    .COUT(\c$2886 ),
    .SUM(\s$2887 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_33_0 (.A(\s$1133 ),
    .B(\c$2094 ),
    .CIN(\c$2096 ),
    .COUT(\c$2888 ),
    .SUM(\s$2889 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_33_1 (.A(\c$2098 ),
    .B(\c$2100 ),
    .CIN(\s$2103 ),
    .COUT(\c$2890 ),
    .SUM(\s$2891 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_33_2 (.A(\s$2105 ),
    .B(\s$2107 ),
    .CIN(\s$2109 ),
    .COUT(\c$2892 ),
    .SUM(\s$2893 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_34_0 (.A(\s$1145 ),
    .B(\c$2102 ),
    .CIN(\c$2104 ),
    .COUT(\c$2894 ),
    .SUM(\s$2895 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_34_1 (.A(\c$2106 ),
    .B(\c$2108 ),
    .CIN(\s$2111 ),
    .COUT(\c$2896 ),
    .SUM(\s$2897 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_34_2 (.A(\s$2113 ),
    .B(\s$2115 ),
    .CIN(\s$2117 ),
    .COUT(\c$2898 ),
    .SUM(\s$2899 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_35_0 (.A(\s$1157 ),
    .B(\c$2110 ),
    .CIN(\c$2112 ),
    .COUT(\c$2900 ),
    .SUM(\s$2901 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_35_1 (.A(\c$2114 ),
    .B(\c$2116 ),
    .CIN(\s$2119 ),
    .COUT(\c$2902 ),
    .SUM(\s$2903 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_35_2 (.A(\s$2121 ),
    .B(\s$2123 ),
    .CIN(\s$2125 ),
    .COUT(\c$2904 ),
    .SUM(\s$2905 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_36_0 (.A(\s$1169 ),
    .B(\c$2118 ),
    .CIN(\c$2120 ),
    .COUT(\c$2906 ),
    .SUM(\s$2907 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_36_1 (.A(\c$2122 ),
    .B(\c$2124 ),
    .CIN(\s$2127 ),
    .COUT(\c$2908 ),
    .SUM(\s$2909 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_36_2 (.A(\s$2129 ),
    .B(\s$2131 ),
    .CIN(\s$2133 ),
    .COUT(\c$2910 ),
    .SUM(\s$2911 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_37_0 (.A(\s$1181 ),
    .B(\c$2126 ),
    .CIN(\c$2128 ),
    .COUT(\c$2912 ),
    .SUM(\s$2913 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_37_1 (.A(\c$2130 ),
    .B(\c$2132 ),
    .CIN(\s$2135 ),
    .COUT(\c$2914 ),
    .SUM(\s$2915 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_37_2 (.A(\s$2137 ),
    .B(\s$2139 ),
    .CIN(\s$2141 ),
    .COUT(\c$2916 ),
    .SUM(\s$2917 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_38_0 (.A(\s$1193 ),
    .B(\c$2134 ),
    .CIN(\c$2136 ),
    .COUT(\c$2918 ),
    .SUM(\s$2919 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_38_1 (.A(\c$2138 ),
    .B(\c$2140 ),
    .CIN(\s$2143 ),
    .COUT(\c$2920 ),
    .SUM(\s$2921 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_38_2 (.A(\s$2145 ),
    .B(\s$2147 ),
    .CIN(\s$2149 ),
    .COUT(\c$2922 ),
    .SUM(\s$2923 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_39_0 (.A(\s$1205 ),
    .B(\c$2142 ),
    .CIN(\c$2144 ),
    .COUT(\c$2924 ),
    .SUM(\s$2925 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_39_1 (.A(\c$2146 ),
    .B(\c$2148 ),
    .CIN(\s$2151 ),
    .COUT(\c$2926 ),
    .SUM(\s$2927 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_39_2 (.A(\s$2153 ),
    .B(\s$2155 ),
    .CIN(\s$2157 ),
    .COUT(\c$2928 ),
    .SUM(\s$2929 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_40_0 (.A(\s$1217 ),
    .B(\c$2150 ),
    .CIN(\c$2152 ),
    .COUT(\c$2930 ),
    .SUM(\s$2931 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_40_1 (.A(\c$2154 ),
    .B(\c$2156 ),
    .CIN(\s$2159 ),
    .COUT(\c$2932 ),
    .SUM(\s$2933 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_40_2 (.A(\s$2161 ),
    .B(\s$2163 ),
    .CIN(\s$2165 ),
    .COUT(\c$2934 ),
    .SUM(\s$2935 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_41_0 (.A(\s$1229 ),
    .B(\c$2158 ),
    .CIN(\c$2160 ),
    .COUT(\c$2936 ),
    .SUM(\s$2937 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_41_1 (.A(\c$2162 ),
    .B(\c$2164 ),
    .CIN(\s$2167 ),
    .COUT(\c$2938 ),
    .SUM(\s$2939 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_41_2 (.A(\s$2169 ),
    .B(\s$2171 ),
    .CIN(\s$2173 ),
    .COUT(\c$2940 ),
    .SUM(\s$2941 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_42_0 (.A(\s$1241 ),
    .B(\c$2166 ),
    .CIN(\c$2168 ),
    .COUT(\c$2942 ),
    .SUM(\s$2943 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_42_1 (.A(\c$2170 ),
    .B(\c$2172 ),
    .CIN(\s$2175 ),
    .COUT(\c$2944 ),
    .SUM(\s$2945 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_42_2 (.A(\s$2177 ),
    .B(\s$2179 ),
    .CIN(\s$2181 ),
    .COUT(\c$2946 ),
    .SUM(\s$2947 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_43_0 (.A(\s$1253 ),
    .B(\c$2174 ),
    .CIN(\c$2176 ),
    .COUT(\c$2948 ),
    .SUM(\s$2949 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_43_1 (.A(\c$2178 ),
    .B(\c$2180 ),
    .CIN(\s$2183 ),
    .COUT(\c$2950 ),
    .SUM(\s$2951 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_43_2 (.A(\s$2185 ),
    .B(\s$2187 ),
    .CIN(\s$2189 ),
    .COUT(\c$2952 ),
    .SUM(\s$2953 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_44_0 (.A(\s$1265 ),
    .B(\c$2182 ),
    .CIN(\c$2184 ),
    .COUT(\c$2954 ),
    .SUM(\s$2955 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_44_1 (.A(\c$2186 ),
    .B(\c$2188 ),
    .CIN(\s$2191 ),
    .COUT(\c$2956 ),
    .SUM(\s$2957 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_44_2 (.A(\s$2193 ),
    .B(\s$2195 ),
    .CIN(\s$2197 ),
    .COUT(\c$2958 ),
    .SUM(\s$2959 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_45_0 (.A(\s$1277 ),
    .B(\c$2190 ),
    .CIN(\c$2192 ),
    .COUT(\c$2960 ),
    .SUM(\s$2961 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_45_1 (.A(\c$2194 ),
    .B(\c$2196 ),
    .CIN(\s$2199 ),
    .COUT(\c$2962 ),
    .SUM(\s$2963 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_45_2 (.A(\s$2201 ),
    .B(\s$2203 ),
    .CIN(\s$2205 ),
    .COUT(\c$2964 ),
    .SUM(\s$2965 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_46_0 (.A(\s$1289 ),
    .B(\c$2198 ),
    .CIN(\c$2200 ),
    .COUT(\c$2966 ),
    .SUM(\s$2967 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_46_1 (.A(\c$2202 ),
    .B(\c$2204 ),
    .CIN(\s$2207 ),
    .COUT(\c$2968 ),
    .SUM(\s$2969 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_46_2 (.A(\s$2209 ),
    .B(\s$2211 ),
    .CIN(\s$2213 ),
    .COUT(\c$2970 ),
    .SUM(\s$2971 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_47_0 (.A(\s$1301 ),
    .B(\c$2206 ),
    .CIN(\c$2208 ),
    .COUT(\c$2972 ),
    .SUM(\s$2973 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_47_1 (.A(\c$2210 ),
    .B(\c$2212 ),
    .CIN(\s$2215 ),
    .COUT(\c$2974 ),
    .SUM(\s$2975 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_47_2 (.A(\s$2217 ),
    .B(\s$2219 ),
    .CIN(\s$2221 ),
    .COUT(\c$2976 ),
    .SUM(\s$2977 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_48_0 (.A(\s$1313 ),
    .B(\c$2214 ),
    .CIN(\c$2216 ),
    .COUT(\c$2978 ),
    .SUM(\s$2979 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_48_1 (.A(\c$2218 ),
    .B(\c$2220 ),
    .CIN(\s$2223 ),
    .COUT(\c$2980 ),
    .SUM(\s$2981 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_48_2 (.A(\s$2225 ),
    .B(\s$2227 ),
    .CIN(\s$2229 ),
    .COUT(\c$2982 ),
    .SUM(\s$2983 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_49_0 (.A(\s$1325 ),
    .B(\c$2222 ),
    .CIN(\c$2224 ),
    .COUT(\c$2984 ),
    .SUM(\s$2985 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_49_1 (.A(\c$2226 ),
    .B(\c$2228 ),
    .CIN(\s$2231 ),
    .COUT(\c$2986 ),
    .SUM(\s$2987 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_49_2 (.A(\s$2233 ),
    .B(\s$2235 ),
    .CIN(\s$2237 ),
    .COUT(\c$2988 ),
    .SUM(\s$2989 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_50_0 (.A(\s$1337 ),
    .B(\c$2230 ),
    .CIN(\c$2232 ),
    .COUT(\c$2990 ),
    .SUM(\s$2991 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_50_1 (.A(\c$2234 ),
    .B(\c$2236 ),
    .CIN(\s$2239 ),
    .COUT(\c$2992 ),
    .SUM(\s$2993 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_50_2 (.A(\s$2241 ),
    .B(\s$2243 ),
    .CIN(\s$2245 ),
    .COUT(\c$2994 ),
    .SUM(\s$2995 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_51_0 (.A(\s$1349 ),
    .B(\c$2238 ),
    .CIN(\c$2240 ),
    .COUT(\c$2996 ),
    .SUM(\s$2997 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_51_1 (.A(\c$2242 ),
    .B(\c$2244 ),
    .CIN(\s$2247 ),
    .COUT(\c$2998 ),
    .SUM(\s$2999 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_51_2 (.A(\s$2249 ),
    .B(\s$2251 ),
    .CIN(\s$2253 ),
    .COUT(\c$3000 ),
    .SUM(\s$3001 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_52_0 (.A(\s$1361 ),
    .B(\c$2246 ),
    .CIN(\c$2248 ),
    .COUT(\c$3002 ),
    .SUM(\s$3003 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_52_1 (.A(\c$2250 ),
    .B(\c$2252 ),
    .CIN(\s$2255 ),
    .COUT(\c$3004 ),
    .SUM(\s$3005 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_52_2 (.A(\s$2257 ),
    .B(\s$2259 ),
    .CIN(\s$2261 ),
    .COUT(\c$3006 ),
    .SUM(\s$3007 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_53_0 (.A(\s$1373 ),
    .B(\c$2254 ),
    .CIN(\c$2256 ),
    .COUT(\c$3008 ),
    .SUM(\s$3009 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_53_1 (.A(\c$2258 ),
    .B(\c$2260 ),
    .CIN(\s$2263 ),
    .COUT(\c$3010 ),
    .SUM(\s$3011 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_53_2 (.A(\s$2265 ),
    .B(\s$2267 ),
    .CIN(\s$2269 ),
    .COUT(\c$3012 ),
    .SUM(\s$3013 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_54_0 (.A(\s$1385 ),
    .B(\c$2262 ),
    .CIN(\c$2264 ),
    .COUT(\c$3014 ),
    .SUM(\s$3015 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_54_1 (.A(\c$2266 ),
    .B(\c$2268 ),
    .CIN(\s$2271 ),
    .COUT(\c$3016 ),
    .SUM(\s$3017 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_54_2 (.A(\s$2273 ),
    .B(\s$2275 ),
    .CIN(\s$2277 ),
    .COUT(\c$3018 ),
    .SUM(\s$3019 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_55_0 (.A(\s$1397 ),
    .B(\c$2270 ),
    .CIN(\c$2272 ),
    .COUT(\c$3020 ),
    .SUM(\s$3021 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_55_1 (.A(\c$2274 ),
    .B(\c$2276 ),
    .CIN(\s$2279 ),
    .COUT(\c$3022 ),
    .SUM(\s$3023 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_55_2 (.A(\s$2281 ),
    .B(\s$2283 ),
    .CIN(\s$2285 ),
    .COUT(\c$3024 ),
    .SUM(\s$3025 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_56_0 (.A(\s$1409 ),
    .B(\c$2278 ),
    .CIN(\c$2280 ),
    .COUT(\c$3026 ),
    .SUM(\s$3027 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_56_1 (.A(\c$2282 ),
    .B(\c$2284 ),
    .CIN(\s$2287 ),
    .COUT(\c$3028 ),
    .SUM(\s$3029 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_56_2 (.A(\s$2289 ),
    .B(\s$2291 ),
    .CIN(\s$2293 ),
    .COUT(\c$3030 ),
    .SUM(\s$3031 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_57_0 (.A(\s$1421 ),
    .B(\c$2286 ),
    .CIN(\c$2288 ),
    .COUT(\c$3032 ),
    .SUM(\s$3033 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_57_1 (.A(\c$2290 ),
    .B(\c$2292 ),
    .CIN(\s$2295 ),
    .COUT(\c$3034 ),
    .SUM(\s$3035 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_57_2 (.A(\s$2297 ),
    .B(\s$2299 ),
    .CIN(\s$2301 ),
    .COUT(\c$3036 ),
    .SUM(\s$3037 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_58_0 (.A(\s$1433 ),
    .B(\c$2294 ),
    .CIN(\c$2296 ),
    .COUT(\c$3038 ),
    .SUM(\s$3039 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_58_1 (.A(\c$2298 ),
    .B(\c$2300 ),
    .CIN(\s$2303 ),
    .COUT(\c$3040 ),
    .SUM(\s$3041 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_58_2 (.A(\s$2305 ),
    .B(\s$2307 ),
    .CIN(\s$2309 ),
    .COUT(\c$3042 ),
    .SUM(\s$3043 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_59_0 (.A(\s$1445 ),
    .B(\c$2302 ),
    .CIN(\c$2304 ),
    .COUT(\c$3044 ),
    .SUM(\s$3045 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_59_1 (.A(\c$2306 ),
    .B(\c$2308 ),
    .CIN(\s$2311 ),
    .COUT(\c$3046 ),
    .SUM(\s$3047 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_59_2 (.A(\s$2313 ),
    .B(\s$2315 ),
    .CIN(\s$2317 ),
    .COUT(\c$3048 ),
    .SUM(\s$3049 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_60_0 (.A(\s$1457 ),
    .B(\c$2310 ),
    .CIN(\c$2312 ),
    .COUT(\c$3050 ),
    .SUM(\s$3051 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_60_1 (.A(\c$2314 ),
    .B(\c$2316 ),
    .CIN(\s$2319 ),
    .COUT(\c$3052 ),
    .SUM(\s$3053 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_60_2 (.A(\s$2321 ),
    .B(\s$2323 ),
    .CIN(\s$2325 ),
    .COUT(\c$3054 ),
    .SUM(\s$3055 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_61_0 (.A(\s$1469 ),
    .B(\c$2318 ),
    .CIN(\c$2320 ),
    .COUT(\c$3056 ),
    .SUM(\s$3057 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_61_1 (.A(\c$2322 ),
    .B(\c$2324 ),
    .CIN(\s$2327 ),
    .COUT(\c$3058 ),
    .SUM(\s$3059 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_61_2 (.A(\s$2329 ),
    .B(\s$2331 ),
    .CIN(\s$2333 ),
    .COUT(\c$3060 ),
    .SUM(\s$3061 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_62_0 (.A(\s$1481 ),
    .B(\c$2326 ),
    .CIN(\c$2328 ),
    .COUT(\c$3062 ),
    .SUM(\s$3063 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_62_1 (.A(\c$2330 ),
    .B(\c$2332 ),
    .CIN(\s$2335 ),
    .COUT(\c$3064 ),
    .SUM(\s$3065 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_62_2 (.A(\s$2337 ),
    .B(\s$2339 ),
    .CIN(\s$2341 ),
    .COUT(\c$3066 ),
    .SUM(\s$3067 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_63_0 (.A(\s$1493 ),
    .B(\c$2334 ),
    .CIN(\c$2336 ),
    .COUT(\c$3068 ),
    .SUM(\s$3069 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_63_1 (.A(\c$2338 ),
    .B(\c$2340 ),
    .CIN(\s$2343 ),
    .COUT(\c$3070 ),
    .SUM(\s$3071 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_63_2 (.A(\s$2345 ),
    .B(\s$2347 ),
    .CIN(\s$2349 ),
    .COUT(\c$3072 ),
    .SUM(\s$3073 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_64_0 (.A(\s$1505 ),
    .B(\c$2342 ),
    .CIN(\c$2344 ),
    .COUT(\c$3074 ),
    .SUM(\s$3075 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_64_1 (.A(\c$2346 ),
    .B(\c$2348 ),
    .CIN(\s$2351 ),
    .COUT(\c$3076 ),
    .SUM(\s$3077 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_64_2 (.A(\s$2353 ),
    .B(\s$2355 ),
    .CIN(\s$2357 ),
    .COUT(\c$3078 ),
    .SUM(\s$3079 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_65_0 (.A(\s$1517 ),
    .B(\c$2350 ),
    .CIN(\c$2352 ),
    .COUT(\c$3080 ),
    .SUM(\s$3081 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_65_1 (.A(\c$2354 ),
    .B(\c$2356 ),
    .CIN(\s$2359 ),
    .COUT(\c$3082 ),
    .SUM(\s$3083 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_65_2 (.A(\s$2361 ),
    .B(\s$2363 ),
    .CIN(\s$2365 ),
    .COUT(\c$3084 ),
    .SUM(\s$3085 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_66_0 (.A(\s$1529 ),
    .B(\c$2358 ),
    .CIN(\c$2360 ),
    .COUT(\c$3086 ),
    .SUM(\s$3087 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_66_1 (.A(\c$2362 ),
    .B(\c$2364 ),
    .CIN(\s$2367 ),
    .COUT(\c$3088 ),
    .SUM(\s$3089 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_66_2 (.A(\s$2369 ),
    .B(\s$2371 ),
    .CIN(\s$2373 ),
    .COUT(\c$3090 ),
    .SUM(\s$3091 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_67_0 (.A(\s$1541 ),
    .B(\c$2366 ),
    .CIN(\c$2368 ),
    .COUT(\c$3092 ),
    .SUM(\s$3093 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_67_1 (.A(\c$2370 ),
    .B(\c$2372 ),
    .CIN(\s$2375 ),
    .COUT(\c$3094 ),
    .SUM(\s$3095 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_67_2 (.A(\s$2377 ),
    .B(\s$2379 ),
    .CIN(\s$2381 ),
    .COUT(\c$3096 ),
    .SUM(\s$3097 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_68_0 (.A(\s$1553 ),
    .B(\c$2374 ),
    .CIN(\c$2376 ),
    .COUT(\c$3098 ),
    .SUM(\s$3099 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_68_1 (.A(\c$2378 ),
    .B(\c$2380 ),
    .CIN(\s$2383 ),
    .COUT(\c$3100 ),
    .SUM(\s$3101 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_68_2 (.A(\s$2385 ),
    .B(\s$2387 ),
    .CIN(\s$2389 ),
    .COUT(\c$3102 ),
    .SUM(\s$3103 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_69_0 (.A(\s$1565 ),
    .B(\c$2382 ),
    .CIN(\c$2384 ),
    .COUT(\c$3104 ),
    .SUM(\s$3105 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_69_1 (.A(\c$2386 ),
    .B(\c$2388 ),
    .CIN(\s$2391 ),
    .COUT(\c$3106 ),
    .SUM(\s$3107 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_69_2 (.A(\s$2393 ),
    .B(\s$2395 ),
    .CIN(\s$2397 ),
    .COUT(\c$3108 ),
    .SUM(\s$3109 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_70_0 (.A(\s$1577 ),
    .B(\c$2390 ),
    .CIN(\c$2392 ),
    .COUT(\c$3110 ),
    .SUM(\s$3111 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_70_1 (.A(\c$2394 ),
    .B(\c$2396 ),
    .CIN(\s$2399 ),
    .COUT(\c$3112 ),
    .SUM(\s$3113 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_70_2 (.A(\s$2401 ),
    .B(\s$2403 ),
    .CIN(\s$2405 ),
    .COUT(\c$3114 ),
    .SUM(\s$3115 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_71_0 (.A(\s$1589 ),
    .B(\c$2398 ),
    .CIN(\c$2400 ),
    .COUT(\c$3116 ),
    .SUM(\s$3117 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_71_1 (.A(\c$2402 ),
    .B(\c$2404 ),
    .CIN(\s$2407 ),
    .COUT(\c$3118 ),
    .SUM(\s$3119 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_71_2 (.A(\s$2409 ),
    .B(\s$2411 ),
    .CIN(\s$2413 ),
    .COUT(\c$3120 ),
    .SUM(\s$3121 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_72_0 (.A(\s$1601 ),
    .B(\c$2406 ),
    .CIN(\c$2408 ),
    .COUT(\c$3122 ),
    .SUM(\s$3123 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_72_1 (.A(\c$2410 ),
    .B(\c$2412 ),
    .CIN(\s$2415 ),
    .COUT(\c$3124 ),
    .SUM(\s$3125 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_72_2 (.A(\s$2417 ),
    .B(\s$2419 ),
    .CIN(\s$2421 ),
    .COUT(\c$3126 ),
    .SUM(\s$3127 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_73_0 (.A(\s$1613 ),
    .B(\c$2414 ),
    .CIN(\c$2416 ),
    .COUT(\c$3128 ),
    .SUM(\s$3129 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_73_1 (.A(\c$2418 ),
    .B(\c$2420 ),
    .CIN(\s$2423 ),
    .COUT(\c$3130 ),
    .SUM(\s$3131 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_73_2 (.A(\s$2425 ),
    .B(\s$2427 ),
    .CIN(\s$2429 ),
    .COUT(\c$3132 ),
    .SUM(\s$3133 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_74_0 (.A(\s$1625 ),
    .B(\c$2422 ),
    .CIN(\c$2424 ),
    .COUT(\c$3134 ),
    .SUM(\s$3135 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_74_1 (.A(\c$2426 ),
    .B(\c$2428 ),
    .CIN(\s$2431 ),
    .COUT(\c$3136 ),
    .SUM(\s$3137 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_74_2 (.A(\s$2433 ),
    .B(\s$2435 ),
    .CIN(\s$2437 ),
    .COUT(\c$3138 ),
    .SUM(\s$3139 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_75_0 (.A(\s$1637 ),
    .B(\c$2430 ),
    .CIN(\c$2432 ),
    .COUT(\c$3140 ),
    .SUM(\s$3141 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_75_1 (.A(\c$2434 ),
    .B(\c$2436 ),
    .CIN(\s$2439 ),
    .COUT(\c$3142 ),
    .SUM(\s$3143 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_75_2 (.A(\s$2441 ),
    .B(\s$2443 ),
    .CIN(\s$2445 ),
    .COUT(\c$3144 ),
    .SUM(\s$3145 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_76_0 (.A(\s$1649 ),
    .B(\c$2438 ),
    .CIN(\c$2440 ),
    .COUT(\c$3146 ),
    .SUM(\s$3147 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_76_1 (.A(\c$2442 ),
    .B(\c$2444 ),
    .CIN(\s$2447 ),
    .COUT(\c$3148 ),
    .SUM(\s$3149 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_76_2 (.A(\s$2449 ),
    .B(\s$2451 ),
    .CIN(\s$2453 ),
    .COUT(\c$3150 ),
    .SUM(\s$3151 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_77_0 (.A(\s$1661 ),
    .B(\c$2446 ),
    .CIN(\c$2448 ),
    .COUT(\c$3152 ),
    .SUM(\s$3153 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_77_1 (.A(\c$2450 ),
    .B(\c$2452 ),
    .CIN(\s$2455 ),
    .COUT(\c$3154 ),
    .SUM(\s$3155 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_77_2 (.A(\s$2457 ),
    .B(\s$2459 ),
    .CIN(\s$2461 ),
    .COUT(\c$3156 ),
    .SUM(\s$3157 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_78_0 (.A(\s$1673 ),
    .B(\c$2454 ),
    .CIN(\c$2456 ),
    .COUT(\c$3158 ),
    .SUM(\s$3159 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_78_1 (.A(\c$2458 ),
    .B(\c$2460 ),
    .CIN(\s$2463 ),
    .COUT(\c$3160 ),
    .SUM(\s$3161 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_78_2 (.A(\s$2465 ),
    .B(\s$2467 ),
    .CIN(\s$2469 ),
    .COUT(\c$3162 ),
    .SUM(\s$3163 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_79_0 (.A(\s$1685 ),
    .B(\c$2462 ),
    .CIN(\c$2464 ),
    .COUT(\c$3164 ),
    .SUM(\s$3165 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_79_1 (.A(\c$2466 ),
    .B(\c$2468 ),
    .CIN(\s$2471 ),
    .COUT(\c$3166 ),
    .SUM(\s$3167 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_79_2 (.A(\s$2473 ),
    .B(\s$2475 ),
    .CIN(\s$2477 ),
    .COUT(\c$3168 ),
    .SUM(\s$3169 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_80_0 (.A(\s$1697 ),
    .B(\c$2470 ),
    .CIN(\c$2472 ),
    .COUT(\c$3170 ),
    .SUM(\s$3171 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_80_1 (.A(\c$2474 ),
    .B(\c$2476 ),
    .CIN(\s$2479 ),
    .COUT(\c$3172 ),
    .SUM(\s$3173 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_80_2 (.A(\s$2481 ),
    .B(\s$2483 ),
    .CIN(\s$2485 ),
    .COUT(\c$3174 ),
    .SUM(\s$3175 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_81_0 (.A(\s$1709 ),
    .B(\c$2478 ),
    .CIN(\c$2480 ),
    .COUT(\c$3176 ),
    .SUM(\s$3177 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_81_1 (.A(\c$2482 ),
    .B(\c$2484 ),
    .CIN(\s$2487 ),
    .COUT(\c$3178 ),
    .SUM(\s$3179 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_81_2 (.A(\s$2489 ),
    .B(\s$2491 ),
    .CIN(\s$2493 ),
    .COUT(\c$3180 ),
    .SUM(\s$3181 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_82_0 (.A(\s$1721 ),
    .B(\c$2486 ),
    .CIN(\c$2488 ),
    .COUT(\c$3182 ),
    .SUM(\s$3183 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_82_1 (.A(\c$2490 ),
    .B(\c$2492 ),
    .CIN(\s$2495 ),
    .COUT(\c$3184 ),
    .SUM(\s$3185 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_82_2 (.A(\s$2497 ),
    .B(\s$2499 ),
    .CIN(\s$2501 ),
    .COUT(\c$3186 ),
    .SUM(\s$3187 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_83_0 (.A(\s$1733 ),
    .B(\c$2494 ),
    .CIN(\c$2496 ),
    .COUT(\c$3188 ),
    .SUM(\s$3189 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_83_1 (.A(\c$2498 ),
    .B(\c$2500 ),
    .CIN(\s$2503 ),
    .COUT(\c$3190 ),
    .SUM(\s$3191 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_83_2 (.A(\s$2505 ),
    .B(\s$2507 ),
    .CIN(\s$2509 ),
    .COUT(\c$3192 ),
    .SUM(\s$3193 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_84_0 (.A(\s$1745 ),
    .B(\c$2502 ),
    .CIN(\c$2504 ),
    .COUT(\c$3194 ),
    .SUM(\s$3195 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_84_1 (.A(\c$2506 ),
    .B(\c$2508 ),
    .CIN(\s$2511 ),
    .COUT(\c$3196 ),
    .SUM(\s$3197 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_84_2 (.A(\s$2513 ),
    .B(\s$2515 ),
    .CIN(\s$2517 ),
    .COUT(\c$3198 ),
    .SUM(\s$3199 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_85_0 (.A(\s$1757 ),
    .B(\c$2510 ),
    .CIN(\c$2512 ),
    .COUT(\c$3200 ),
    .SUM(\s$3201 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_85_1 (.A(\c$2514 ),
    .B(\c$2516 ),
    .CIN(\s$2519 ),
    .COUT(\c$3202 ),
    .SUM(\s$3203 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_85_2 (.A(\s$2521 ),
    .B(\s$2523 ),
    .CIN(\s$2525 ),
    .COUT(\c$3204 ),
    .SUM(\s$3205 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_86_0 (.A(\s$1769 ),
    .B(\c$2518 ),
    .CIN(\c$2520 ),
    .COUT(\c$3206 ),
    .SUM(\s$3207 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_86_1 (.A(\c$2522 ),
    .B(\c$2524 ),
    .CIN(\s$2527 ),
    .COUT(\c$3208 ),
    .SUM(\s$3209 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_86_2 (.A(\s$2529 ),
    .B(\s$2531 ),
    .CIN(\s$2533 ),
    .COUT(\c$3210 ),
    .SUM(\s$3211 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_87_0 (.A(\s$1781 ),
    .B(\c$2526 ),
    .CIN(\c$2528 ),
    .COUT(\c$3212 ),
    .SUM(\s$3213 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_87_1 (.A(\c$2530 ),
    .B(\c$2532 ),
    .CIN(\s$2535 ),
    .COUT(\c$3214 ),
    .SUM(\s$3215 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_87_2 (.A(\s$2537 ),
    .B(\s$2539 ),
    .CIN(\s$2541 ),
    .COUT(\c$3216 ),
    .SUM(\s$3217 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_88_0 (.A(\s$1793 ),
    .B(\c$2534 ),
    .CIN(\c$2536 ),
    .COUT(\c$3218 ),
    .SUM(\s$3219 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_88_1 (.A(\c$2538 ),
    .B(\c$2540 ),
    .CIN(\s$2543 ),
    .COUT(\c$3220 ),
    .SUM(\s$3221 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_88_2 (.A(\s$2545 ),
    .B(\s$2547 ),
    .CIN(\s$2549 ),
    .COUT(\c$3222 ),
    .SUM(\s$3223 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_89_0 (.A(\s$1805 ),
    .B(\c$2542 ),
    .CIN(\c$2544 ),
    .COUT(\c$3224 ),
    .SUM(\s$3225 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_89_1 (.A(\c$2546 ),
    .B(\c$2548 ),
    .CIN(\s$2551 ),
    .COUT(\c$3226 ),
    .SUM(\s$3227 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_89_2 (.A(\s$2553 ),
    .B(\s$2555 ),
    .CIN(\s$2557 ),
    .COUT(\c$3228 ),
    .SUM(\s$3229 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_90_0 (.A(\s$1817 ),
    .B(\c$2550 ),
    .CIN(\c$2552 ),
    .COUT(\c$3230 ),
    .SUM(\s$3231 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_90_1 (.A(\c$2554 ),
    .B(\c$2556 ),
    .CIN(\s$2559 ),
    .COUT(\c$3232 ),
    .SUM(\s$3233 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_90_2 (.A(\s$2561 ),
    .B(\s$2563 ),
    .CIN(\s$2565 ),
    .COUT(\c$3234 ),
    .SUM(\s$3235 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_91_0 (.A(\s$1829 ),
    .B(\c$2558 ),
    .CIN(\c$2560 ),
    .COUT(\c$3236 ),
    .SUM(\s$3237 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_91_1 (.A(\c$2562 ),
    .B(\c$2564 ),
    .CIN(\s$2567 ),
    .COUT(\c$3238 ),
    .SUM(\s$3239 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_91_2 (.A(\s$2569 ),
    .B(\s$2571 ),
    .CIN(\s$2573 ),
    .COUT(\c$3240 ),
    .SUM(\s$3241 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_92_0 (.A(\s$1841 ),
    .B(\c$2566 ),
    .CIN(\c$2568 ),
    .COUT(\c$3242 ),
    .SUM(\s$3243 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_92_1 (.A(\c$2570 ),
    .B(\c$2572 ),
    .CIN(\s$2575 ),
    .COUT(\c$3244 ),
    .SUM(\s$3245 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_92_2 (.A(\s$2577 ),
    .B(\s$2579 ),
    .CIN(\s$2581 ),
    .COUT(\c$3246 ),
    .SUM(\s$3247 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_93_0 (.A(\s$1853 ),
    .B(\c$2574 ),
    .CIN(\c$2576 ),
    .COUT(\c$3248 ),
    .SUM(\s$3249 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_93_1 (.A(\c$2578 ),
    .B(\c$2580 ),
    .CIN(\s$2583 ),
    .COUT(\c$3250 ),
    .SUM(\s$3251 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_93_2 (.A(\s$2585 ),
    .B(\s$2587 ),
    .CIN(\s$2589 ),
    .COUT(\c$3252 ),
    .SUM(\s$3253 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_94_0 (.A(\s$1865 ),
    .B(\c$2582 ),
    .CIN(\c$2584 ),
    .COUT(\c$3254 ),
    .SUM(\s$3255 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_94_1 (.A(\c$2586 ),
    .B(\c$2588 ),
    .CIN(\s$2591 ),
    .COUT(\c$3256 ),
    .SUM(\s$3257 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_94_2 (.A(\s$2593 ),
    .B(\s$2595 ),
    .CIN(\s$2597 ),
    .COUT(\c$3258 ),
    .SUM(\s$3259 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_95_0 (.A(\s$1877 ),
    .B(\c$2590 ),
    .CIN(\c$2592 ),
    .COUT(\c$3260 ),
    .SUM(\s$3261 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_95_1 (.A(\c$2594 ),
    .B(\c$2596 ),
    .CIN(\s$2599 ),
    .COUT(\c$3262 ),
    .SUM(\s$3263 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_95_2 (.A(\s$2601 ),
    .B(\s$2603 ),
    .CIN(\s$2605 ),
    .COUT(\c$3264 ),
    .SUM(\s$3265 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_96_0 (.A(\s$1889 ),
    .B(\c$2598 ),
    .CIN(\c$2600 ),
    .COUT(\c$3266 ),
    .SUM(\s$3267 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_96_1 (.A(\c$2602 ),
    .B(\c$2604 ),
    .CIN(\s$2607 ),
    .COUT(\c$3268 ),
    .SUM(\s$3269 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_96_2 (.A(\s$2609 ),
    .B(\s$2611 ),
    .CIN(\s$2613 ),
    .COUT(\c$3270 ),
    .SUM(\s$3271 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_97_0 (.A(\s$1901 ),
    .B(\c$2606 ),
    .CIN(\c$2608 ),
    .COUT(\c$3272 ),
    .SUM(\s$3273 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_97_1 (.A(\c$2610 ),
    .B(\c$2612 ),
    .CIN(\s$2615 ),
    .COUT(\c$3274 ),
    .SUM(\s$3275 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_97_2 (.A(\s$2617 ),
    .B(\s$2619 ),
    .CIN(\s$2621 ),
    .COUT(\c$3276 ),
    .SUM(\s$3277 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_98_0 (.A(\s$1913 ),
    .B(\c$2614 ),
    .CIN(\c$2616 ),
    .COUT(\c$3278 ),
    .SUM(\s$3279 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_98_1 (.A(\c$2618 ),
    .B(\c$2620 ),
    .CIN(\s$2623 ),
    .COUT(\c$3280 ),
    .SUM(\s$3281 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_98_2 (.A(\s$2625 ),
    .B(\s$2627 ),
    .CIN(\s$2629 ),
    .COUT(\c$3282 ),
    .SUM(\s$3283 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_99_0 (.A(\s$1923 ),
    .B(\c$2622 ),
    .CIN(\c$2624 ),
    .COUT(\c$3284 ),
    .SUM(\s$3285 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_99_1 (.A(\c$2626 ),
    .B(\c$2628 ),
    .CIN(\s$2631 ),
    .COUT(\c$3286 ),
    .SUM(\s$3287 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_4_99_2 (.A(\s$2633 ),
    .B(\s$2635 ),
    .CIN(\s$2637 ),
    .COUT(\c$3288 ),
    .SUM(\s$3289 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_100_0 (.A(\c$3284 ),
    .B(\c$3286 ),
    .CIN(\c$3288 ),
    .COUT(\c$3796 ),
    .SUM(\s$3797 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_100_1 (.A(\s$3291 ),
    .B(\s$3293 ),
    .CIN(\s$3295 ),
    .COUT(\c$3798 ),
    .SUM(\s$3799 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_101_0 (.A(\c$3290 ),
    .B(\c$3292 ),
    .CIN(\c$3294 ),
    .COUT(\c$3800 ),
    .SUM(\s$3801 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_101_1 (.A(\s$3297 ),
    .B(\s$3299 ),
    .CIN(\s$3301 ),
    .COUT(\c$3802 ),
    .SUM(\s$3803 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_102_0 (.A(\c$3296 ),
    .B(\c$3298 ),
    .CIN(\c$3300 ),
    .COUT(\c$3804 ),
    .SUM(\s$3805 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_102_1 (.A(\s$3303 ),
    .B(\s$3305 ),
    .CIN(\s$3307 ),
    .COUT(\c$3806 ),
    .SUM(\s$3807 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_103_0 (.A(\c$3302 ),
    .B(\c$3304 ),
    .CIN(\c$3306 ),
    .COUT(\c$3808 ),
    .SUM(\s$3809 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_103_1 (.A(\s$3309 ),
    .B(\s$3311 ),
    .CIN(\s$3313 ),
    .COUT(\c$3810 ),
    .SUM(\s$3811 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_104_0 (.A(\c$3308 ),
    .B(\c$3310 ),
    .CIN(\c$3312 ),
    .COUT(\c$3812 ),
    .SUM(\s$3813 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_104_1 (.A(\s$3315 ),
    .B(\s$3317 ),
    .CIN(\s$3319 ),
    .COUT(\c$3814 ),
    .SUM(\s$3815 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_105_0 (.A(\c$3314 ),
    .B(\c$3316 ),
    .CIN(\c$3318 ),
    .COUT(\c$3816 ),
    .SUM(\s$3817 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_105_1 (.A(\s$3321 ),
    .B(\s$3323 ),
    .CIN(\s$3325 ),
    .COUT(\c$3818 ),
    .SUM(\s$3819 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_106_0 (.A(\c$3320 ),
    .B(\c$3322 ),
    .CIN(\c$3324 ),
    .COUT(\c$3820 ),
    .SUM(\s$3821 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_106_1 (.A(\s$3327 ),
    .B(\s$3329 ),
    .CIN(\s$3331 ),
    .COUT(\c$3822 ),
    .SUM(\s$3823 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_107_0 (.A(\c$3326 ),
    .B(\c$3328 ),
    .CIN(\c$3330 ),
    .COUT(\c$3824 ),
    .SUM(\s$3825 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_107_1 (.A(\s$3333 ),
    .B(\s$3335 ),
    .CIN(\s$3337 ),
    .COUT(\c$3826 ),
    .SUM(\s$3827 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_108_0 (.A(\c$3332 ),
    .B(\c$3334 ),
    .CIN(\c$3336 ),
    .COUT(\c$3828 ),
    .SUM(\s$3829 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_108_1 (.A(\s$3339 ),
    .B(\s$3341 ),
    .CIN(\s$3343 ),
    .COUT(\c$3830 ),
    .SUM(\s$3831 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_109_0 (.A(\c$3338 ),
    .B(\c$3340 ),
    .CIN(\c$3342 ),
    .COUT(\c$3832 ),
    .SUM(\s$3833 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_109_1 (.A(\s$3345 ),
    .B(\s$3347 ),
    .CIN(\s$3349 ),
    .COUT(\c$3834 ),
    .SUM(\s$3835 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_10_0 (.A(pp_row10_5),
    .B(pp_row10_6),
    .CIN(pp_row10_7),
    .COUT(\c$3436 ),
    .SUM(\s$3437 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_10_1 (.A(\c$2752 ),
    .B(\s$2755 ),
    .CIN(\s$2757 ),
    .COUT(\c$3438 ),
    .SUM(\s$3439 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_110_0 (.A(\c$3344 ),
    .B(\c$3346 ),
    .CIN(\c$3348 ),
    .COUT(\c$3836 ),
    .SUM(\s$3837 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_110_1 (.A(\s$3351 ),
    .B(\s$3353 ),
    .CIN(\s$3355 ),
    .COUT(\c$3838 ),
    .SUM(\s$3839 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_111_0 (.A(\c$3350 ),
    .B(\c$3352 ),
    .CIN(\c$3354 ),
    .COUT(\c$3840 ),
    .SUM(\s$3841 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_111_1 (.A(\s$3357 ),
    .B(\s$3359 ),
    .CIN(\s$3361 ),
    .COUT(\c$3842 ),
    .SUM(\s$3843 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_112_0 (.A(\c$3356 ),
    .B(\c$3358 ),
    .CIN(\c$3360 ),
    .COUT(\c$3844 ),
    .SUM(\s$3845 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_112_1 (.A(\s$3363 ),
    .B(\s$3365 ),
    .CIN(\s$3367 ),
    .COUT(\c$3846 ),
    .SUM(\s$3847 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_113_0 (.A(\c$3362 ),
    .B(\c$3364 ),
    .CIN(\c$3366 ),
    .COUT(\c$3848 ),
    .SUM(\s$3849 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_113_1 (.A(\s$3369 ),
    .B(\s$3371 ),
    .CIN(\s$3373 ),
    .COUT(\c$3850 ),
    .SUM(\s$3851 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_114_0 (.A(\c$3368 ),
    .B(\c$3370 ),
    .CIN(\c$3372 ),
    .COUT(\c$3852 ),
    .SUM(\s$3853 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_114_1 (.A(\s$3375 ),
    .B(\s$3377 ),
    .CIN(\s$3379 ),
    .COUT(\c$3854 ),
    .SUM(\s$3855 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_115_0 (.A(\c$3374 ),
    .B(\c$3376 ),
    .CIN(\c$3378 ),
    .COUT(\c$3856 ),
    .SUM(\s$3857 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_115_1 (.A(\s$3381 ),
    .B(\s$3383 ),
    .CIN(\s$3385 ),
    .COUT(\c$3858 ),
    .SUM(\s$3859 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_116_0 (.A(\c$3380 ),
    .B(\c$3382 ),
    .CIN(\c$3384 ),
    .COUT(\c$3860 ),
    .SUM(\s$3861 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_116_1 (.A(\s$3387 ),
    .B(\s$3389 ),
    .CIN(\s$3391 ),
    .COUT(\c$3862 ),
    .SUM(\s$3863 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_117_0 (.A(\c$3386 ),
    .B(\c$3388 ),
    .CIN(\c$3390 ),
    .COUT(\c$3864 ),
    .SUM(\s$3865 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_117_1 (.A(\s$3393 ),
    .B(\s$3395 ),
    .CIN(\s$3397 ),
    .COUT(\c$3866 ),
    .SUM(\s$3867 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_118_0 (.A(\c$3392 ),
    .B(\c$3394 ),
    .CIN(\c$3396 ),
    .COUT(\c$3868 ),
    .SUM(\s$3869 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_118_1 (.A(\s$3399 ),
    .B(\s$3401 ),
    .CIN(\s$3403 ),
    .COUT(\c$3870 ),
    .SUM(\s$3871 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_119_0 (.A(pp_row119_6),
    .B(\c$3398 ),
    .CIN(\c$3400 ),
    .COUT(\c$3872 ),
    .SUM(\s$3873 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_119_1 (.A(\c$3402 ),
    .B(\s$3405 ),
    .CIN(\s$3407 ),
    .COUT(\c$3874 ),
    .SUM(\s$3875 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_11_0 (.A(pp_row11_5),
    .B(pp_row11_6),
    .CIN(\c$2754 ),
    .COUT(\c$3440 ),
    .SUM(\s$3441 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_11_1 (.A(\c$2756 ),
    .B(\s$2759 ),
    .CIN(\s$2761 ),
    .COUT(\c$3442 ),
    .SUM(\s$3443 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_120_0 (.A(pp_row120_5),
    .B(pp_row120_6),
    .CIN(\c$3404 ),
    .COUT(\c$3876 ),
    .SUM(\s$3877 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_120_1 (.A(\c$3406 ),
    .B(\s$3409 ),
    .CIN(\s$3411 ),
    .COUT(\c$3878 ),
    .SUM(\s$3879 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_121_0 (.A(pp_row121_3),
    .B(pp_row121_4),
    .CIN(pp_row121_5),
    .COUT(\c$3880 ),
    .SUM(\s$3881 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_121_1 (.A(\c$3408 ),
    .B(\c$3410 ),
    .CIN(\s$3413 ),
    .COUT(\c$3882 ),
    .SUM(\s$3883 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_122_0 (.A(pp_row122_2),
    .B(pp_row122_3),
    .CIN(pp_row122_4),
    .COUT(\c$3884 ),
    .SUM(\s$3885 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_122_1 (.A(pp_row122_5),
    .B(\c$3412 ),
    .CIN(\s$3415 ),
    .COUT(\c$3886 ),
    .SUM(\s$3887 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_123_0 (.A(pp_row123_0),
    .B(pp_row123_1),
    .CIN(pp_row123_2),
    .COUT(\c$3888 ),
    .SUM(\s$3889 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_123_1 (.A(pp_row123_3),
    .B(pp_row123_4),
    .CIN(\c$3414 ),
    .COUT(\c$3890 ),
    .SUM(\s$3891 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_124_0 (.A(net1914),
    .B(pp_row124_1),
    .CIN(pp_row124_2),
    .COUT(\c$3892 ),
    .SUM(\s$3893 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_125_0 (.A(pp_row125_0),
    .B(pp_row125_1),
    .CIN(pp_row125_2),
    .COUT(\c$3896 ),
    .SUM(\s$3897 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_12_0 (.A(pp_row12_8),
    .B(\c$2758 ),
    .CIN(\c$2760 ),
    .COUT(\c$3444 ),
    .SUM(\s$3445 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_12_1 (.A(\s$2763 ),
    .B(\s$2765 ),
    .CIN(\s$2767 ),
    .COUT(\c$3446 ),
    .SUM(\s$3447 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_13_0 (.A(\c$2762 ),
    .B(\c$2764 ),
    .CIN(\c$2766 ),
    .COUT(\c$3448 ),
    .SUM(\s$3449 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_13_1 (.A(\s$2769 ),
    .B(\s$2771 ),
    .CIN(\s$2773 ),
    .COUT(\c$3450 ),
    .SUM(\s$3451 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_14_0 (.A(\c$2768 ),
    .B(\c$2770 ),
    .CIN(\c$2772 ),
    .COUT(\c$3452 ),
    .SUM(\s$3453 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_14_1 (.A(\s$2775 ),
    .B(\s$2777 ),
    .CIN(\s$2779 ),
    .COUT(\c$3454 ),
    .SUM(\s$3455 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_15_0 (.A(\c$2774 ),
    .B(\c$2776 ),
    .CIN(\c$2778 ),
    .COUT(\c$3456 ),
    .SUM(\s$3457 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_15_1 (.A(\s$2781 ),
    .B(\s$2783 ),
    .CIN(\s$2785 ),
    .COUT(\c$3458 ),
    .SUM(\s$3459 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_16_0 (.A(\c$2780 ),
    .B(\c$2782 ),
    .CIN(\c$2784 ),
    .COUT(\c$3460 ),
    .SUM(\s$3461 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_16_1 (.A(\s$2787 ),
    .B(\s$2789 ),
    .CIN(\s$2791 ),
    .COUT(\c$3462 ),
    .SUM(\s$3463 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_17_0 (.A(\c$2786 ),
    .B(\c$2788 ),
    .CIN(\c$2790 ),
    .COUT(\c$3464 ),
    .SUM(\s$3465 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_17_1 (.A(\s$2793 ),
    .B(\s$2795 ),
    .CIN(\s$2797 ),
    .COUT(\c$3466 ),
    .SUM(\s$3467 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_18_0 (.A(\c$2792 ),
    .B(\c$2794 ),
    .CIN(\c$2796 ),
    .COUT(\c$3468 ),
    .SUM(\s$3469 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_18_1 (.A(\s$2799 ),
    .B(\s$2801 ),
    .CIN(\s$2803 ),
    .COUT(\c$3470 ),
    .SUM(\s$3471 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_19_0 (.A(\c$2798 ),
    .B(\c$2800 ),
    .CIN(\c$2802 ),
    .COUT(\c$3472 ),
    .SUM(\s$3473 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_19_1 (.A(\s$2805 ),
    .B(\s$2807 ),
    .CIN(\s$2809 ),
    .COUT(\c$3474 ),
    .SUM(\s$3475 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_20_0 (.A(\c$2804 ),
    .B(\c$2806 ),
    .CIN(\c$2808 ),
    .COUT(\c$3476 ),
    .SUM(\s$3477 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_20_1 (.A(\s$2811 ),
    .B(\s$2813 ),
    .CIN(\s$2815 ),
    .COUT(\c$3478 ),
    .SUM(\s$3479 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_21_0 (.A(\c$2810 ),
    .B(\c$2812 ),
    .CIN(\c$2814 ),
    .COUT(\c$3480 ),
    .SUM(\s$3481 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_21_1 (.A(\s$2817 ),
    .B(\s$2819 ),
    .CIN(\s$2821 ),
    .COUT(\c$3482 ),
    .SUM(\s$3483 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_22_0 (.A(\c$2816 ),
    .B(\c$2818 ),
    .CIN(\c$2820 ),
    .COUT(\c$3484 ),
    .SUM(\s$3485 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_22_1 (.A(\s$2823 ),
    .B(\s$2825 ),
    .CIN(\s$2827 ),
    .COUT(\c$3486 ),
    .SUM(\s$3487 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_23_0 (.A(\c$2822 ),
    .B(\c$2824 ),
    .CIN(\c$2826 ),
    .COUT(\c$3488 ),
    .SUM(\s$3489 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_23_1 (.A(\s$2829 ),
    .B(\s$2831 ),
    .CIN(\s$2833 ),
    .COUT(\c$3490 ),
    .SUM(\s$3491 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_24_0 (.A(\c$2828 ),
    .B(\c$2830 ),
    .CIN(\c$2832 ),
    .COUT(\c$3492 ),
    .SUM(\s$3493 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_24_1 (.A(\s$2835 ),
    .B(\s$2837 ),
    .CIN(\s$2839 ),
    .COUT(\c$3494 ),
    .SUM(\s$3495 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_25_0 (.A(\c$2834 ),
    .B(\c$2836 ),
    .CIN(\c$2838 ),
    .COUT(\c$3496 ),
    .SUM(\s$3497 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_25_1 (.A(\s$2841 ),
    .B(\s$2843 ),
    .CIN(\s$2845 ),
    .COUT(\c$3498 ),
    .SUM(\s$3499 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_26_0 (.A(\c$2840 ),
    .B(\c$2842 ),
    .CIN(\c$2844 ),
    .COUT(\c$3500 ),
    .SUM(\s$3501 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_26_1 (.A(\s$2847 ),
    .B(\s$2849 ),
    .CIN(\s$2851 ),
    .COUT(\c$3502 ),
    .SUM(\s$3503 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_27_0 (.A(\c$2846 ),
    .B(\c$2848 ),
    .CIN(\c$2850 ),
    .COUT(\c$3504 ),
    .SUM(\s$3505 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_27_1 (.A(\s$2853 ),
    .B(\s$2855 ),
    .CIN(\s$2857 ),
    .COUT(\c$3506 ),
    .SUM(\s$3507 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_28_0 (.A(\c$2852 ),
    .B(\c$2854 ),
    .CIN(\c$2856 ),
    .COUT(\c$3508 ),
    .SUM(\s$3509 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_28_1 (.A(\s$2859 ),
    .B(\s$2861 ),
    .CIN(\s$2863 ),
    .COUT(\c$3510 ),
    .SUM(\s$3511 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_29_0 (.A(\c$2858 ),
    .B(\c$2860 ),
    .CIN(\c$2862 ),
    .COUT(\c$3512 ),
    .SUM(\s$3513 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_29_1 (.A(\s$2865 ),
    .B(\s$2867 ),
    .CIN(\s$2869 ),
    .COUT(\c$3514 ),
    .SUM(\s$3515 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_30_0 (.A(\c$2864 ),
    .B(\c$2866 ),
    .CIN(\c$2868 ),
    .COUT(\c$3516 ),
    .SUM(\s$3517 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_30_1 (.A(\s$2871 ),
    .B(\s$2873 ),
    .CIN(\s$2875 ),
    .COUT(\c$3518 ),
    .SUM(\s$3519 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_31_0 (.A(\c$2870 ),
    .B(\c$2872 ),
    .CIN(\c$2874 ),
    .COUT(\c$3520 ),
    .SUM(\s$3521 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_31_1 (.A(\s$2877 ),
    .B(\s$2879 ),
    .CIN(\s$2881 ),
    .COUT(\c$3522 ),
    .SUM(\s$3523 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_32_0 (.A(\c$2876 ),
    .B(\c$2878 ),
    .CIN(\c$2880 ),
    .COUT(\c$3524 ),
    .SUM(\s$3525 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_32_1 (.A(\s$2883 ),
    .B(\s$2885 ),
    .CIN(\s$2887 ),
    .COUT(\c$3526 ),
    .SUM(\s$3527 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_33_0 (.A(\c$2882 ),
    .B(\c$2884 ),
    .CIN(\c$2886 ),
    .COUT(\c$3528 ),
    .SUM(\s$3529 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_33_1 (.A(\s$2889 ),
    .B(\s$2891 ),
    .CIN(\s$2893 ),
    .COUT(\c$3530 ),
    .SUM(\s$3531 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_34_0 (.A(\c$2888 ),
    .B(\c$2890 ),
    .CIN(\c$2892 ),
    .COUT(\c$3532 ),
    .SUM(\s$3533 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_34_1 (.A(\s$2895 ),
    .B(\s$2897 ),
    .CIN(\s$2899 ),
    .COUT(\c$3534 ),
    .SUM(\s$3535 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_35_0 (.A(\c$2894 ),
    .B(\c$2896 ),
    .CIN(\c$2898 ),
    .COUT(\c$3536 ),
    .SUM(\s$3537 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_35_1 (.A(\s$2901 ),
    .B(\s$2903 ),
    .CIN(\s$2905 ),
    .COUT(\c$3538 ),
    .SUM(\s$3539 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_36_0 (.A(\c$2900 ),
    .B(\c$2902 ),
    .CIN(\c$2904 ),
    .COUT(\c$3540 ),
    .SUM(\s$3541 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_36_1 (.A(\s$2907 ),
    .B(\s$2909 ),
    .CIN(\s$2911 ),
    .COUT(\c$3542 ),
    .SUM(\s$3543 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_37_0 (.A(\c$2906 ),
    .B(\c$2908 ),
    .CIN(\c$2910 ),
    .COUT(\c$3544 ),
    .SUM(\s$3545 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_37_1 (.A(\s$2913 ),
    .B(\s$2915 ),
    .CIN(\s$2917 ),
    .COUT(\c$3546 ),
    .SUM(\s$3547 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_38_0 (.A(\c$2912 ),
    .B(\c$2914 ),
    .CIN(\c$2916 ),
    .COUT(\c$3548 ),
    .SUM(\s$3549 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_38_1 (.A(\s$2919 ),
    .B(\s$2921 ),
    .CIN(\s$2923 ),
    .COUT(\c$3550 ),
    .SUM(\s$3551 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_39_0 (.A(\c$2918 ),
    .B(\c$2920 ),
    .CIN(\c$2922 ),
    .COUT(\c$3552 ),
    .SUM(\s$3553 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_39_1 (.A(\s$2925 ),
    .B(\s$2927 ),
    .CIN(\s$2929 ),
    .COUT(\c$3554 ),
    .SUM(\s$3555 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_40_0 (.A(\c$2924 ),
    .B(\c$2926 ),
    .CIN(\c$2928 ),
    .COUT(\c$3556 ),
    .SUM(\s$3557 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_40_1 (.A(\s$2931 ),
    .B(\s$2933 ),
    .CIN(\s$2935 ),
    .COUT(\c$3558 ),
    .SUM(\s$3559 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_41_0 (.A(\c$2930 ),
    .B(\c$2932 ),
    .CIN(\c$2934 ),
    .COUT(\c$3560 ),
    .SUM(\s$3561 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_41_1 (.A(\s$2937 ),
    .B(\s$2939 ),
    .CIN(\s$2941 ),
    .COUT(\c$3562 ),
    .SUM(\s$3563 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_42_0 (.A(\c$2936 ),
    .B(\c$2938 ),
    .CIN(\c$2940 ),
    .COUT(\c$3564 ),
    .SUM(\s$3565 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_42_1 (.A(\s$2943 ),
    .B(\s$2945 ),
    .CIN(\s$2947 ),
    .COUT(\c$3566 ),
    .SUM(\s$3567 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_43_0 (.A(\c$2942 ),
    .B(\c$2944 ),
    .CIN(\c$2946 ),
    .COUT(\c$3568 ),
    .SUM(\s$3569 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_43_1 (.A(\s$2949 ),
    .B(\s$2951 ),
    .CIN(\s$2953 ),
    .COUT(\c$3570 ),
    .SUM(\s$3571 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_44_0 (.A(\c$2948 ),
    .B(\c$2950 ),
    .CIN(\c$2952 ),
    .COUT(\c$3572 ),
    .SUM(\s$3573 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_44_1 (.A(\s$2955 ),
    .B(\s$2957 ),
    .CIN(\s$2959 ),
    .COUT(\c$3574 ),
    .SUM(\s$3575 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_45_0 (.A(\c$2954 ),
    .B(\c$2956 ),
    .CIN(\c$2958 ),
    .COUT(\c$3576 ),
    .SUM(\s$3577 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_45_1 (.A(\s$2961 ),
    .B(\s$2963 ),
    .CIN(\s$2965 ),
    .COUT(\c$3578 ),
    .SUM(\s$3579 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_46_0 (.A(\c$2960 ),
    .B(\c$2962 ),
    .CIN(\c$2964 ),
    .COUT(\c$3580 ),
    .SUM(\s$3581 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_46_1 (.A(\s$2967 ),
    .B(\s$2969 ),
    .CIN(\s$2971 ),
    .COUT(\c$3582 ),
    .SUM(\s$3583 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_47_0 (.A(\c$2966 ),
    .B(\c$2968 ),
    .CIN(\c$2970 ),
    .COUT(\c$3584 ),
    .SUM(\s$3585 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_47_1 (.A(\s$2973 ),
    .B(\s$2975 ),
    .CIN(\s$2977 ),
    .COUT(\c$3586 ),
    .SUM(\s$3587 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_48_0 (.A(\c$2972 ),
    .B(\c$2974 ),
    .CIN(\c$2976 ),
    .COUT(\c$3588 ),
    .SUM(\s$3589 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_48_1 (.A(\s$2979 ),
    .B(\s$2981 ),
    .CIN(\s$2983 ),
    .COUT(\c$3590 ),
    .SUM(\s$3591 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_49_0 (.A(\c$2978 ),
    .B(\c$2980 ),
    .CIN(\c$2982 ),
    .COUT(\c$3592 ),
    .SUM(\s$3593 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_49_1 (.A(\s$2985 ),
    .B(\s$2987 ),
    .CIN(\s$2989 ),
    .COUT(\c$3594 ),
    .SUM(\s$3595 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_50_0 (.A(\c$2984 ),
    .B(\c$2986 ),
    .CIN(\c$2988 ),
    .COUT(\c$3596 ),
    .SUM(\s$3597 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_50_1 (.A(\s$2991 ),
    .B(\s$2993 ),
    .CIN(\s$2995 ),
    .COUT(\c$3598 ),
    .SUM(\s$3599 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_51_0 (.A(\c$2990 ),
    .B(\c$2992 ),
    .CIN(\c$2994 ),
    .COUT(\c$3600 ),
    .SUM(\s$3601 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_51_1 (.A(\s$2997 ),
    .B(\s$2999 ),
    .CIN(\s$3001 ),
    .COUT(\c$3602 ),
    .SUM(\s$3603 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_52_0 (.A(\c$2996 ),
    .B(\c$2998 ),
    .CIN(\c$3000 ),
    .COUT(\c$3604 ),
    .SUM(\s$3605 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_52_1 (.A(\s$3003 ),
    .B(\s$3005 ),
    .CIN(\s$3007 ),
    .COUT(\c$3606 ),
    .SUM(\s$3607 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_53_0 (.A(\c$3002 ),
    .B(\c$3004 ),
    .CIN(\c$3006 ),
    .COUT(\c$3608 ),
    .SUM(\s$3609 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_53_1 (.A(\s$3009 ),
    .B(\s$3011 ),
    .CIN(\s$3013 ),
    .COUT(\c$3610 ),
    .SUM(\s$3611 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_54_0 (.A(\c$3008 ),
    .B(\c$3010 ),
    .CIN(\c$3012 ),
    .COUT(\c$3612 ),
    .SUM(\s$3613 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_54_1 (.A(\s$3015 ),
    .B(\s$3017 ),
    .CIN(\s$3019 ),
    .COUT(\c$3614 ),
    .SUM(\s$3615 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_55_0 (.A(\c$3014 ),
    .B(\c$3016 ),
    .CIN(\c$3018 ),
    .COUT(\c$3616 ),
    .SUM(\s$3617 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_55_1 (.A(\s$3021 ),
    .B(\s$3023 ),
    .CIN(\s$3025 ),
    .COUT(\c$3618 ),
    .SUM(\s$3619 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_56_0 (.A(\c$3020 ),
    .B(\c$3022 ),
    .CIN(\c$3024 ),
    .COUT(\c$3620 ),
    .SUM(\s$3621 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_56_1 (.A(\s$3027 ),
    .B(\s$3029 ),
    .CIN(\s$3031 ),
    .COUT(\c$3622 ),
    .SUM(\s$3623 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_57_0 (.A(\c$3026 ),
    .B(\c$3028 ),
    .CIN(\c$3030 ),
    .COUT(\c$3624 ),
    .SUM(\s$3625 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_57_1 (.A(\s$3033 ),
    .B(\s$3035 ),
    .CIN(\s$3037 ),
    .COUT(\c$3626 ),
    .SUM(\s$3627 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_58_0 (.A(\c$3032 ),
    .B(\c$3034 ),
    .CIN(\c$3036 ),
    .COUT(\c$3628 ),
    .SUM(\s$3629 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_58_1 (.A(\s$3039 ),
    .B(\s$3041 ),
    .CIN(\s$3043 ),
    .COUT(\c$3630 ),
    .SUM(\s$3631 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_59_0 (.A(\c$3038 ),
    .B(\c$3040 ),
    .CIN(\c$3042 ),
    .COUT(\c$3632 ),
    .SUM(\s$3633 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_59_1 (.A(\s$3045 ),
    .B(\s$3047 ),
    .CIN(\s$3049 ),
    .COUT(\c$3634 ),
    .SUM(\s$3635 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_60_0 (.A(\c$3044 ),
    .B(\c$3046 ),
    .CIN(\c$3048 ),
    .COUT(\c$3636 ),
    .SUM(\s$3637 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_60_1 (.A(\s$3051 ),
    .B(\s$3053 ),
    .CIN(\s$3055 ),
    .COUT(\c$3638 ),
    .SUM(\s$3639 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_61_0 (.A(\c$3050 ),
    .B(\c$3052 ),
    .CIN(\c$3054 ),
    .COUT(\c$3640 ),
    .SUM(\s$3641 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_61_1 (.A(\s$3057 ),
    .B(\s$3059 ),
    .CIN(\s$3061 ),
    .COUT(\c$3642 ),
    .SUM(\s$3643 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_62_0 (.A(\c$3056 ),
    .B(\c$3058 ),
    .CIN(\c$3060 ),
    .COUT(\c$3644 ),
    .SUM(\s$3645 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_62_1 (.A(\s$3063 ),
    .B(\s$3065 ),
    .CIN(\s$3067 ),
    .COUT(\c$3646 ),
    .SUM(\s$3647 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_63_0 (.A(\c$3062 ),
    .B(\c$3064 ),
    .CIN(\c$3066 ),
    .COUT(\c$3648 ),
    .SUM(\s$3649 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_63_1 (.A(\s$3069 ),
    .B(\s$3071 ),
    .CIN(\s$3073 ),
    .COUT(\c$3650 ),
    .SUM(\s$3651 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_64_0 (.A(\c$3068 ),
    .B(\c$3070 ),
    .CIN(\c$3072 ),
    .COUT(\c$3652 ),
    .SUM(\s$3653 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_64_1 (.A(\s$3075 ),
    .B(\s$3077 ),
    .CIN(\s$3079 ),
    .COUT(\c$3654 ),
    .SUM(\s$3655 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_65_0 (.A(\c$3074 ),
    .B(\c$3076 ),
    .CIN(\c$3078 ),
    .COUT(\c$3656 ),
    .SUM(\s$3657 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_65_1 (.A(\s$3081 ),
    .B(\s$3083 ),
    .CIN(\s$3085 ),
    .COUT(\c$3658 ),
    .SUM(\s$3659 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_66_0 (.A(\c$3080 ),
    .B(\c$3082 ),
    .CIN(\c$3084 ),
    .COUT(\c$3660 ),
    .SUM(\s$3661 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_66_1 (.A(\s$3087 ),
    .B(\s$3089 ),
    .CIN(\s$3091 ),
    .COUT(\c$3662 ),
    .SUM(\s$3663 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_67_0 (.A(\c$3086 ),
    .B(\c$3088 ),
    .CIN(\c$3090 ),
    .COUT(\c$3664 ),
    .SUM(\s$3665 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_67_1 (.A(\s$3093 ),
    .B(\s$3095 ),
    .CIN(\s$3097 ),
    .COUT(\c$3666 ),
    .SUM(\s$3667 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_68_0 (.A(\c$3092 ),
    .B(\c$3094 ),
    .CIN(\c$3096 ),
    .COUT(\c$3668 ),
    .SUM(\s$3669 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_68_1 (.A(\s$3099 ),
    .B(\s$3101 ),
    .CIN(\s$3103 ),
    .COUT(\c$3670 ),
    .SUM(\s$3671 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_69_0 (.A(\c$3098 ),
    .B(\c$3100 ),
    .CIN(\c$3102 ),
    .COUT(\c$3672 ),
    .SUM(\s$3673 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_69_1 (.A(\s$3105 ),
    .B(\s$3107 ),
    .CIN(\s$3109 ),
    .COUT(\c$3674 ),
    .SUM(\s$3675 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_6_0 (.A(pp_row6_0),
    .B(pp_row6_1),
    .CIN(pp_row6_2),
    .COUT(\c$3420 ),
    .SUM(\s$3421 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_70_0 (.A(\c$3104 ),
    .B(\c$3106 ),
    .CIN(\c$3108 ),
    .COUT(\c$3676 ),
    .SUM(\s$3677 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_70_1 (.A(\s$3111 ),
    .B(\s$3113 ),
    .CIN(\s$3115 ),
    .COUT(\c$3678 ),
    .SUM(\s$3679 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_71_0 (.A(\c$3110 ),
    .B(\c$3112 ),
    .CIN(\c$3114 ),
    .COUT(\c$3680 ),
    .SUM(\s$3681 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_71_1 (.A(\s$3117 ),
    .B(\s$3119 ),
    .CIN(\s$3121 ),
    .COUT(\c$3682 ),
    .SUM(\s$3683 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_72_0 (.A(\c$3116 ),
    .B(\c$3118 ),
    .CIN(\c$3120 ),
    .COUT(\c$3684 ),
    .SUM(\s$3685 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_72_1 (.A(\s$3123 ),
    .B(\s$3125 ),
    .CIN(\s$3127 ),
    .COUT(\c$3686 ),
    .SUM(\s$3687 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_73_0 (.A(\c$3122 ),
    .B(\c$3124 ),
    .CIN(\c$3126 ),
    .COUT(\c$3688 ),
    .SUM(\s$3689 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_73_1 (.A(\s$3129 ),
    .B(\s$3131 ),
    .CIN(\s$3133 ),
    .COUT(\c$3690 ),
    .SUM(\s$3691 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_74_0 (.A(\c$3128 ),
    .B(\c$3130 ),
    .CIN(\c$3132 ),
    .COUT(\c$3692 ),
    .SUM(\s$3693 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_74_1 (.A(\s$3135 ),
    .B(\s$3137 ),
    .CIN(\s$3139 ),
    .COUT(\c$3694 ),
    .SUM(\s$3695 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_75_0 (.A(\c$3134 ),
    .B(\c$3136 ),
    .CIN(\c$3138 ),
    .COUT(\c$3696 ),
    .SUM(\s$3697 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_75_1 (.A(\s$3141 ),
    .B(\s$3143 ),
    .CIN(\s$3145 ),
    .COUT(\c$3698 ),
    .SUM(\s$3699 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_76_0 (.A(\c$3140 ),
    .B(\c$3142 ),
    .CIN(\c$3144 ),
    .COUT(\c$3700 ),
    .SUM(\s$3701 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_76_1 (.A(\s$3147 ),
    .B(\s$3149 ),
    .CIN(\s$3151 ),
    .COUT(\c$3702 ),
    .SUM(\s$3703 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_77_0 (.A(\c$3146 ),
    .B(\c$3148 ),
    .CIN(\c$3150 ),
    .COUT(\c$3704 ),
    .SUM(\s$3705 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_77_1 (.A(\s$3153 ),
    .B(\s$3155 ),
    .CIN(\s$3157 ),
    .COUT(\c$3706 ),
    .SUM(\s$3707 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_78_0 (.A(\c$3152 ),
    .B(\c$3154 ),
    .CIN(\c$3156 ),
    .COUT(\c$3708 ),
    .SUM(\s$3709 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_78_1 (.A(\s$3159 ),
    .B(\s$3161 ),
    .CIN(\s$3163 ),
    .COUT(\c$3710 ),
    .SUM(\s$3711 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_79_0 (.A(\c$3158 ),
    .B(\c$3160 ),
    .CIN(\c$3162 ),
    .COUT(\c$3712 ),
    .SUM(\s$3713 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_79_1 (.A(\s$3165 ),
    .B(\s$3167 ),
    .CIN(\s$3169 ),
    .COUT(\c$3714 ),
    .SUM(\s$3715 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_7_0 (.A(pp_row7_0),
    .B(pp_row7_1),
    .CIN(pp_row7_2),
    .COUT(\c$3424 ),
    .SUM(\s$3425 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_80_0 (.A(\c$3164 ),
    .B(\c$3166 ),
    .CIN(\c$3168 ),
    .COUT(\c$3716 ),
    .SUM(\s$3717 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_80_1 (.A(\s$3171 ),
    .B(\s$3173 ),
    .CIN(\s$3175 ),
    .COUT(\c$3718 ),
    .SUM(\s$3719 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_81_0 (.A(\c$3170 ),
    .B(\c$3172 ),
    .CIN(\c$3174 ),
    .COUT(\c$3720 ),
    .SUM(\s$3721 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_81_1 (.A(\s$3177 ),
    .B(\s$3179 ),
    .CIN(\s$3181 ),
    .COUT(\c$3722 ),
    .SUM(\s$3723 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_82_0 (.A(\c$3176 ),
    .B(\c$3178 ),
    .CIN(\c$3180 ),
    .COUT(\c$3724 ),
    .SUM(\s$3725 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_82_1 (.A(\s$3183 ),
    .B(\s$3185 ),
    .CIN(\s$3187 ),
    .COUT(\c$3726 ),
    .SUM(\s$3727 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_83_0 (.A(\c$3182 ),
    .B(\c$3184 ),
    .CIN(\c$3186 ),
    .COUT(\c$3728 ),
    .SUM(\s$3729 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_83_1 (.A(\s$3189 ),
    .B(\s$3191 ),
    .CIN(\s$3193 ),
    .COUT(\c$3730 ),
    .SUM(\s$3731 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_84_0 (.A(\c$3188 ),
    .B(\c$3190 ),
    .CIN(\c$3192 ),
    .COUT(\c$3732 ),
    .SUM(\s$3733 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_84_1 (.A(\s$3195 ),
    .B(\s$3197 ),
    .CIN(\s$3199 ),
    .COUT(\c$3734 ),
    .SUM(\s$3735 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_85_0 (.A(\c$3194 ),
    .B(\c$3196 ),
    .CIN(\c$3198 ),
    .COUT(\c$3736 ),
    .SUM(\s$3737 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_85_1 (.A(\s$3201 ),
    .B(\s$3203 ),
    .CIN(\s$3205 ),
    .COUT(\c$3738 ),
    .SUM(\s$3739 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_86_0 (.A(\c$3200 ),
    .B(\c$3202 ),
    .CIN(\c$3204 ),
    .COUT(\c$3740 ),
    .SUM(\s$3741 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_86_1 (.A(\s$3207 ),
    .B(\s$3209 ),
    .CIN(\s$3211 ),
    .COUT(\c$3742 ),
    .SUM(\s$3743 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_87_0 (.A(\c$3206 ),
    .B(\c$3208 ),
    .CIN(\c$3210 ),
    .COUT(\c$3744 ),
    .SUM(\s$3745 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_87_1 (.A(\s$3213 ),
    .B(\s$3215 ),
    .CIN(\s$3217 ),
    .COUT(\c$3746 ),
    .SUM(\s$3747 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_88_0 (.A(\c$3212 ),
    .B(\c$3214 ),
    .CIN(\c$3216 ),
    .COUT(\c$3748 ),
    .SUM(\s$3749 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_88_1 (.A(\s$3219 ),
    .B(\s$3221 ),
    .CIN(\s$3223 ),
    .COUT(\c$3750 ),
    .SUM(\s$3751 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_89_0 (.A(\c$3218 ),
    .B(\c$3220 ),
    .CIN(\c$3222 ),
    .COUT(\c$3752 ),
    .SUM(\s$3753 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_89_1 (.A(\s$3225 ),
    .B(\s$3227 ),
    .CIN(\s$3229 ),
    .COUT(\c$3754 ),
    .SUM(\s$3755 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_8_0 (.A(pp_row8_2),
    .B(pp_row8_3),
    .CIN(pp_row8_4),
    .COUT(\c$3428 ),
    .SUM(\s$3429 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_8_1 (.A(pp_row8_5),
    .B(pp_row8_6),
    .CIN(\s$2751 ),
    .COUT(\c$3430 ),
    .SUM(\s$3431 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_5_90_0 (.A(\c$3224 ),
    .B(\c$3226 ),
    .CIN(\c$3228 ),
    .COUT(\c$3756 ),
    .SUM(\s$3757 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_90_1 (.A(\s$3231 ),
    .B(\s$3233 ),
    .CIN(\s$3235 ),
    .COUT(\c$3758 ),
    .SUM(\s$3759 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_91_0 (.A(\c$3230 ),
    .B(\c$3232 ),
    .CIN(\c$3234 ),
    .COUT(\c$3760 ),
    .SUM(\s$3761 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_91_1 (.A(\s$3237 ),
    .B(\s$3239 ),
    .CIN(\s$3241 ),
    .COUT(\c$3762 ),
    .SUM(\s$3763 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_92_0 (.A(\c$3236 ),
    .B(\c$3238 ),
    .CIN(\c$3240 ),
    .COUT(\c$3764 ),
    .SUM(\s$3765 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_92_1 (.A(\s$3243 ),
    .B(\s$3245 ),
    .CIN(\s$3247 ),
    .COUT(\c$3766 ),
    .SUM(\s$3767 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_93_0 (.A(\c$3242 ),
    .B(\c$3244 ),
    .CIN(\c$3246 ),
    .COUT(\c$3768 ),
    .SUM(\s$3769 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_93_1 (.A(\s$3249 ),
    .B(\s$3251 ),
    .CIN(\s$3253 ),
    .COUT(\c$3770 ),
    .SUM(\s$3771 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_94_0 (.A(\c$3248 ),
    .B(\c$3250 ),
    .CIN(\c$3252 ),
    .COUT(\c$3772 ),
    .SUM(\s$3773 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_94_1 (.A(\s$3255 ),
    .B(\s$3257 ),
    .CIN(\s$3259 ),
    .COUT(\c$3774 ),
    .SUM(\s$3775 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_95_0 (.A(\c$3254 ),
    .B(\c$3256 ),
    .CIN(\c$3258 ),
    .COUT(\c$3776 ),
    .SUM(\s$3777 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_95_1 (.A(\s$3261 ),
    .B(\s$3263 ),
    .CIN(\s$3265 ),
    .COUT(\c$3778 ),
    .SUM(\s$3779 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_96_0 (.A(\c$3260 ),
    .B(\c$3262 ),
    .CIN(\c$3264 ),
    .COUT(\c$3780 ),
    .SUM(\s$3781 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_96_1 (.A(\s$3267 ),
    .B(\s$3269 ),
    .CIN(\s$3271 ),
    .COUT(\c$3782 ),
    .SUM(\s$3783 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_97_0 (.A(\c$3266 ),
    .B(\c$3268 ),
    .CIN(\c$3270 ),
    .COUT(\c$3784 ),
    .SUM(\s$3785 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_97_1 (.A(\s$3273 ),
    .B(\s$3275 ),
    .CIN(\s$3277 ),
    .COUT(\c$3786 ),
    .SUM(\s$3787 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_98_0 (.A(\c$3272 ),
    .B(\c$3274 ),
    .CIN(\c$3276 ),
    .COUT(\c$3788 ),
    .SUM(\s$3789 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_98_1 (.A(\s$3279 ),
    .B(\s$3281 ),
    .CIN(\s$3283 ),
    .COUT(\c$3790 ),
    .SUM(\s$3791 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_99_0 (.A(\c$3278 ),
    .B(\c$3280 ),
    .CIN(\c$3282 ),
    .COUT(\c$3792 ),
    .SUM(\s$3793 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_99_1 (.A(\s$3285 ),
    .B(\s$3287 ),
    .CIN(\s$3289 ),
    .COUT(\c$3794 ),
    .SUM(\s$3795 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_9_0 (.A(pp_row9_2),
    .B(pp_row9_3),
    .CIN(pp_row9_4),
    .COUT(\c$3432 ),
    .SUM(\s$3433 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_5_9_1 (.A(pp_row9_5),
    .B(\c$2750 ),
    .CIN(\s$2753 ),
    .COUT(\c$3434 ),
    .SUM(\s$3435 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_100_0 (.A(\c$3792 ),
    .B(\c$3794 ),
    .CIN(\s$3797 ),
    .COUT(\c$4096 ),
    .SUM(\s$4097 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_101_0 (.A(\c$3796 ),
    .B(\c$3798 ),
    .CIN(\s$3801 ),
    .COUT(\c$4098 ),
    .SUM(\s$4099 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_102_0 (.A(\c$3800 ),
    .B(\c$3802 ),
    .CIN(\s$3805 ),
    .COUT(\c$4100 ),
    .SUM(\s$4101 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_103_0 (.A(\c$3804 ),
    .B(\c$3806 ),
    .CIN(\s$3809 ),
    .COUT(\c$4102 ),
    .SUM(\s$4103 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_104_0 (.A(\c$3808 ),
    .B(\c$3810 ),
    .CIN(\s$3813 ),
    .COUT(\c$4104 ),
    .SUM(\s$4105 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_105_0 (.A(\c$3812 ),
    .B(\c$3814 ),
    .CIN(\s$3817 ),
    .COUT(\c$4106 ),
    .SUM(\s$4107 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_106_0 (.A(\c$3816 ),
    .B(\c$3818 ),
    .CIN(\s$3821 ),
    .COUT(\c$4108 ),
    .SUM(\s$4109 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_107_0 (.A(\c$3820 ),
    .B(\c$3822 ),
    .CIN(\s$3825 ),
    .COUT(\c$4110 ),
    .SUM(\s$4111 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_108_0 (.A(\c$3824 ),
    .B(\c$3826 ),
    .CIN(\s$3829 ),
    .COUT(\c$4112 ),
    .SUM(\s$4113 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_109_0 (.A(\c$3828 ),
    .B(\c$3830 ),
    .CIN(\s$3833 ),
    .COUT(\c$4114 ),
    .SUM(\s$4115 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_10_0 (.A(\c$3432 ),
    .B(\c$3434 ),
    .CIN(\s$3437 ),
    .COUT(\c$3916 ),
    .SUM(\s$3917 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_110_0 (.A(\c$3832 ),
    .B(\c$3834 ),
    .CIN(\s$3837 ),
    .COUT(\c$4116 ),
    .SUM(\s$4117 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_111_0 (.A(\c$3836 ),
    .B(\c$3838 ),
    .CIN(\s$3841 ),
    .COUT(\c$4118 ),
    .SUM(\s$4119 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_112_0 (.A(\c$3840 ),
    .B(\c$3842 ),
    .CIN(\s$3845 ),
    .COUT(\c$4120 ),
    .SUM(\s$4121 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_113_0 (.A(\c$3844 ),
    .B(\c$3846 ),
    .CIN(\s$3849 ),
    .COUT(\c$4122 ),
    .SUM(\s$4123 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_114_0 (.A(\c$3848 ),
    .B(\c$3850 ),
    .CIN(\s$3853 ),
    .COUT(\c$4124 ),
    .SUM(\s$4125 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_115_0 (.A(\c$3852 ),
    .B(\c$3854 ),
    .CIN(\s$3857 ),
    .COUT(\c$4126 ),
    .SUM(\s$4127 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_116_0 (.A(\c$3856 ),
    .B(\c$3858 ),
    .CIN(\s$3861 ),
    .COUT(\c$4128 ),
    .SUM(\s$4129 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_117_0 (.A(\c$3860 ),
    .B(\c$3862 ),
    .CIN(\s$3865 ),
    .COUT(\c$4130 ),
    .SUM(\s$4131 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_118_0 (.A(\c$3864 ),
    .B(\c$3866 ),
    .CIN(\s$3869 ),
    .COUT(\c$4132 ),
    .SUM(\s$4133 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_119_0 (.A(\c$3868 ),
    .B(\c$3870 ),
    .CIN(\s$3873 ),
    .COUT(\c$4134 ),
    .SUM(\s$4135 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_11_0 (.A(\c$3436 ),
    .B(\c$3438 ),
    .CIN(\s$3441 ),
    .COUT(\c$3918 ),
    .SUM(\s$3919 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_120_0 (.A(\c$3872 ),
    .B(\c$3874 ),
    .CIN(\s$3877 ),
    .COUT(\c$4136 ),
    .SUM(\s$4137 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_121_0 (.A(\c$3876 ),
    .B(\c$3878 ),
    .CIN(\s$3881 ),
    .COUT(\c$4138 ),
    .SUM(\s$4139 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_122_0 (.A(\c$3880 ),
    .B(\c$3882 ),
    .CIN(\s$3885 ),
    .COUT(\c$4140 ),
    .SUM(\s$4141 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_123_0 (.A(\c$3884 ),
    .B(\c$3886 ),
    .CIN(\s$3889 ),
    .COUT(\c$4142 ),
    .SUM(\s$4143 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_124_0 (.A(\c$3888 ),
    .B(\c$3890 ),
    .CIN(\s$3893 ),
    .COUT(\c$4144 ),
    .SUM(\s$4145 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_6_125_0 (.A(pp_row125_3),
    .B(\c$3892 ),
    .CIN(\c$3894 ),
    .COUT(\c$4146 ),
    .SUM(\s$4147 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_126_0 (.A(pp_row126_2),
    .B(pp_row126_3),
    .CIN(\c$3896 ),
    .COUT(\c$4148 ),
    .SUM(\s$4149 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_127_0 (.A(pp_row127_0),
    .B(pp_row127_1),
    .CIN(pp_row127_2),
    .COUT(\c$4150 ),
    .SUM(\s$4151 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_12_0 (.A(\c$3440 ),
    .B(\c$3442 ),
    .CIN(\s$3445 ),
    .COUT(\c$3920 ),
    .SUM(\s$3921 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_13_0 (.A(\c$3444 ),
    .B(\c$3446 ),
    .CIN(\s$3449 ),
    .COUT(\c$3922 ),
    .SUM(\s$3923 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_14_0 (.A(\c$3448 ),
    .B(\c$3450 ),
    .CIN(\s$3453 ),
    .COUT(\c$3924 ),
    .SUM(\s$3925 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_6_15_0 (.A(\c$3452 ),
    .B(\c$3454 ),
    .CIN(\s$3457 ),
    .COUT(\c$3926 ),
    .SUM(\s$3927 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_16_0 (.A(\c$3456 ),
    .B(\c$3458 ),
    .CIN(\s$3461 ),
    .COUT(\c$3928 ),
    .SUM(\s$3929 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_17_0 (.A(\c$3460 ),
    .B(\c$3462 ),
    .CIN(\s$3465 ),
    .COUT(\c$3930 ),
    .SUM(\s$3931 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_6_18_0 (.A(\c$3464 ),
    .B(\c$3466 ),
    .CIN(\s$3469 ),
    .COUT(\c$3932 ),
    .SUM(\s$3933 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_19_0 (.A(\c$3468 ),
    .B(\c$3470 ),
    .CIN(\s$3473 ),
    .COUT(\c$3934 ),
    .SUM(\s$3935 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_20_0 (.A(\c$3472 ),
    .B(\c$3474 ),
    .CIN(\s$3477 ),
    .COUT(\c$3936 ),
    .SUM(\s$3937 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_21_0 (.A(\c$3476 ),
    .B(\c$3478 ),
    .CIN(\s$3481 ),
    .COUT(\c$3938 ),
    .SUM(\s$3939 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_22_0 (.A(\c$3480 ),
    .B(\c$3482 ),
    .CIN(\s$3485 ),
    .COUT(\c$3940 ),
    .SUM(\s$3941 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_23_0 (.A(\c$3484 ),
    .B(\c$3486 ),
    .CIN(\s$3489 ),
    .COUT(\c$3942 ),
    .SUM(\s$3943 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_24_0 (.A(\c$3488 ),
    .B(\c$3490 ),
    .CIN(\s$3493 ),
    .COUT(\c$3944 ),
    .SUM(\s$3945 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_25_0 (.A(\c$3492 ),
    .B(\c$3494 ),
    .CIN(\s$3497 ),
    .COUT(\c$3946 ),
    .SUM(\s$3947 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_26_0 (.A(\c$3496 ),
    .B(\c$3498 ),
    .CIN(\s$3501 ),
    .COUT(\c$3948 ),
    .SUM(\s$3949 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_6_27_0 (.A(\c$3500 ),
    .B(\c$3502 ),
    .CIN(\s$3505 ),
    .COUT(\c$3950 ),
    .SUM(\s$3951 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_28_0 (.A(\c$3504 ),
    .B(\c$3506 ),
    .CIN(\s$3509 ),
    .COUT(\c$3952 ),
    .SUM(\s$3953 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_29_0 (.A(\c$3508 ),
    .B(\c$3510 ),
    .CIN(\s$3513 ),
    .COUT(\c$3954 ),
    .SUM(\s$3955 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_30_0 (.A(\c$3512 ),
    .B(\c$3514 ),
    .CIN(\s$3517 ),
    .COUT(\c$3956 ),
    .SUM(\s$3957 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_31_0 (.A(\c$3516 ),
    .B(\c$3518 ),
    .CIN(\s$3521 ),
    .COUT(\c$3958 ),
    .SUM(\s$3959 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_6_32_0 (.A(\c$3520 ),
    .B(\c$3522 ),
    .CIN(\s$3525 ),
    .COUT(\c$3960 ),
    .SUM(\s$3961 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_6_33_0 (.A(\c$3524 ),
    .B(\c$3526 ),
    .CIN(\s$3529 ),
    .COUT(\c$3962 ),
    .SUM(\s$3963 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_34_0 (.A(\c$3528 ),
    .B(\c$3530 ),
    .CIN(\s$3533 ),
    .COUT(\c$3964 ),
    .SUM(\s$3965 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_35_0 (.A(\c$3532 ),
    .B(\c$3534 ),
    .CIN(\s$3537 ),
    .COUT(\c$3966 ),
    .SUM(\s$3967 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_36_0 (.A(\c$3536 ),
    .B(\c$3538 ),
    .CIN(\s$3541 ),
    .COUT(\c$3968 ),
    .SUM(\s$3969 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_37_0 (.A(\c$3540 ),
    .B(\c$3542 ),
    .CIN(\s$3545 ),
    .COUT(\c$3970 ),
    .SUM(\s$3971 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_38_0 (.A(\c$3544 ),
    .B(\c$3546 ),
    .CIN(\s$3549 ),
    .COUT(\c$3972 ),
    .SUM(\s$3973 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_39_0 (.A(\c$3548 ),
    .B(\c$3550 ),
    .CIN(\s$3553 ),
    .COUT(\c$3974 ),
    .SUM(\s$3975 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_40_0 (.A(\c$3552 ),
    .B(\c$3554 ),
    .CIN(\s$3557 ),
    .COUT(\c$3976 ),
    .SUM(\s$3977 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_41_0 (.A(\c$3556 ),
    .B(\c$3558 ),
    .CIN(\s$3561 ),
    .COUT(\c$3978 ),
    .SUM(\s$3979 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_42_0 (.A(\c$3560 ),
    .B(\c$3562 ),
    .CIN(\s$3565 ),
    .COUT(\c$3980 ),
    .SUM(\s$3981 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_43_0 (.A(\c$3564 ),
    .B(\c$3566 ),
    .CIN(\s$3569 ),
    .COUT(\c$3982 ),
    .SUM(\s$3983 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_44_0 (.A(\c$3568 ),
    .B(\c$3570 ),
    .CIN(\s$3573 ),
    .COUT(\c$3984 ),
    .SUM(\s$3985 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_6_45_0 (.A(\c$3572 ),
    .B(\c$3574 ),
    .CIN(\s$3577 ),
    .COUT(\c$3986 ),
    .SUM(\s$3987 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_46_0 (.A(\c$3576 ),
    .B(\c$3578 ),
    .CIN(\s$3581 ),
    .COUT(\c$3988 ),
    .SUM(\s$3989 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_47_0 (.A(\c$3580 ),
    .B(\c$3582 ),
    .CIN(\s$3585 ),
    .COUT(\c$3990 ),
    .SUM(\s$3991 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_48_0 (.A(\c$3584 ),
    .B(\c$3586 ),
    .CIN(\s$3589 ),
    .COUT(\c$3992 ),
    .SUM(\s$3993 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_49_0 (.A(\c$3588 ),
    .B(\c$3590 ),
    .CIN(\s$3593 ),
    .COUT(\c$3994 ),
    .SUM(\s$3995 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_4_0 (.A(pp_row4_2),
    .B(pp_row4_3),
    .CIN(pp_row4_4),
    .COUT(\c$3904 ),
    .SUM(\s$3905 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_6_50_0 (.A(\c$3592 ),
    .B(\c$3594 ),
    .CIN(\s$3597 ),
    .COUT(\c$3996 ),
    .SUM(\s$3997 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_6_51_0 (.A(\c$3596 ),
    .B(\c$3598 ),
    .CIN(\s$3601 ),
    .COUT(\c$3998 ),
    .SUM(\s$3999 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_6_52_0 (.A(\c$3600 ),
    .B(\c$3602 ),
    .CIN(\s$3605 ),
    .COUT(\c$4000 ),
    .SUM(\s$4001 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_53_0 (.A(\c$3604 ),
    .B(\c$3606 ),
    .CIN(\s$3609 ),
    .COUT(\c$4002 ),
    .SUM(\s$4003 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_54_0 (.A(\c$3608 ),
    .B(\c$3610 ),
    .CIN(\s$3613 ),
    .COUT(\c$4004 ),
    .SUM(\s$4005 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_55_0 (.A(\c$3612 ),
    .B(\c$3614 ),
    .CIN(\s$3617 ),
    .COUT(\c$4006 ),
    .SUM(\s$4007 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_56_0 (.A(\c$3616 ),
    .B(\c$3618 ),
    .CIN(\s$3621 ),
    .COUT(\c$4008 ),
    .SUM(\s$4009 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_57_0 (.A(\c$3620 ),
    .B(\c$3622 ),
    .CIN(\s$3625 ),
    .COUT(\c$4010 ),
    .SUM(\s$4011 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_58_0 (.A(\c$3624 ),
    .B(\c$3626 ),
    .CIN(\s$3629 ),
    .COUT(\c$4012 ),
    .SUM(\s$4013 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_59_0 (.A(\c$3628 ),
    .B(\c$3630 ),
    .CIN(\s$3633 ),
    .COUT(\c$4014 ),
    .SUM(\s$4015 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_5_0 (.A(pp_row5_2),
    .B(pp_row5_3),
    .CIN(\c$3416 ),
    .COUT(\c$3906 ),
    .SUM(\s$3907 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_60_0 (.A(\c$3632 ),
    .B(\c$3634 ),
    .CIN(\s$3637 ),
    .COUT(\c$4016 ),
    .SUM(\s$4017 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_61_0 (.A(\c$3636 ),
    .B(\c$3638 ),
    .CIN(\s$3641 ),
    .COUT(\c$4018 ),
    .SUM(\s$4019 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_62_0 (.A(\c$3640 ),
    .B(\c$3642 ),
    .CIN(\s$3645 ),
    .COUT(\c$4020 ),
    .SUM(\s$4021 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_63_0 (.A(\c$3644 ),
    .B(\c$3646 ),
    .CIN(\s$3649 ),
    .COUT(\c$4022 ),
    .SUM(\s$4023 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_64_0 (.A(\c$3648 ),
    .B(\c$3650 ),
    .CIN(\s$3653 ),
    .COUT(\c$4024 ),
    .SUM(\s$4025 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_6_65_0 (.A(\c$3652 ),
    .B(\c$3654 ),
    .CIN(\s$3657 ),
    .COUT(\c$4026 ),
    .SUM(\s$4027 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_66_0 (.A(\c$3656 ),
    .B(\c$3658 ),
    .CIN(\s$3661 ),
    .COUT(\c$4028 ),
    .SUM(\s$4029 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_67_0 (.A(\c$3660 ),
    .B(\c$3662 ),
    .CIN(\s$3665 ),
    .COUT(\c$4030 ),
    .SUM(\s$4031 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_68_0 (.A(\c$3664 ),
    .B(\c$3666 ),
    .CIN(\s$3669 ),
    .COUT(\c$4032 ),
    .SUM(\s$4033 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_69_0 (.A(\c$3668 ),
    .B(\c$3670 ),
    .CIN(\s$3673 ),
    .COUT(\c$4034 ),
    .SUM(\s$4035 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_6_0 (.A(pp_row6_5),
    .B(\c$3418 ),
    .CIN(\s$3421 ),
    .COUT(\c$3908 ),
    .SUM(\s$3909 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_70_0 (.A(\c$3672 ),
    .B(\c$3674 ),
    .CIN(\s$3677 ),
    .COUT(\c$4036 ),
    .SUM(\s$4037 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_71_0 (.A(\c$3676 ),
    .B(\c$3678 ),
    .CIN(\s$3681 ),
    .COUT(\c$4038 ),
    .SUM(\s$4039 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_72_0 (.A(\c$3680 ),
    .B(\c$3682 ),
    .CIN(\s$3685 ),
    .COUT(\c$4040 ),
    .SUM(\s$4041 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_73_0 (.A(\c$3684 ),
    .B(\c$3686 ),
    .CIN(\s$3689 ),
    .COUT(\c$4042 ),
    .SUM(\s$4043 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_74_0 (.A(\c$3688 ),
    .B(\c$3690 ),
    .CIN(\s$3693 ),
    .COUT(\c$4044 ),
    .SUM(\s$4045 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_75_0 (.A(\c$3692 ),
    .B(\c$3694 ),
    .CIN(\s$3697 ),
    .COUT(\c$4046 ),
    .SUM(\s$4047 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_76_0 (.A(\c$3696 ),
    .B(\c$3698 ),
    .CIN(\s$3701 ),
    .COUT(\c$4048 ),
    .SUM(\s$4049 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_77_0 (.A(\c$3700 ),
    .B(\c$3702 ),
    .CIN(\s$3705 ),
    .COUT(\c$4050 ),
    .SUM(\s$4051 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_78_0 (.A(\c$3704 ),
    .B(\c$3706 ),
    .CIN(\s$3709 ),
    .COUT(\c$4052 ),
    .SUM(\s$4053 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_79_0 (.A(\c$3708 ),
    .B(\c$3710 ),
    .CIN(\s$3713 ),
    .COUT(\c$4054 ),
    .SUM(\s$4055 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_7_0 (.A(\c$3420 ),
    .B(\c$3422 ),
    .CIN(\s$3425 ),
    .COUT(\c$3910 ),
    .SUM(\s$3911 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_80_0 (.A(\c$3712 ),
    .B(\c$3714 ),
    .CIN(\s$3717 ),
    .COUT(\c$4056 ),
    .SUM(\s$4057 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_81_0 (.A(\c$3716 ),
    .B(\c$3718 ),
    .CIN(\s$3721 ),
    .COUT(\c$4058 ),
    .SUM(\s$4059 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_82_0 (.A(\c$3720 ),
    .B(\c$3722 ),
    .CIN(\s$3725 ),
    .COUT(\c$4060 ),
    .SUM(\s$4061 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_83_0 (.A(\c$3724 ),
    .B(\c$3726 ),
    .CIN(\s$3729 ),
    .COUT(\c$4062 ),
    .SUM(\s$4063 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_84_0 (.A(\c$3728 ),
    .B(\c$3730 ),
    .CIN(\s$3733 ),
    .COUT(\c$4064 ),
    .SUM(\s$4065 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_85_0 (.A(\c$3732 ),
    .B(\c$3734 ),
    .CIN(\s$3737 ),
    .COUT(\c$4066 ),
    .SUM(\s$4067 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_86_0 (.A(\c$3736 ),
    .B(\c$3738 ),
    .CIN(\s$3741 ),
    .COUT(\c$4068 ),
    .SUM(\s$4069 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_6_87_0 (.A(\c$3740 ),
    .B(\c$3742 ),
    .CIN(\s$3745 ),
    .COUT(\c$4070 ),
    .SUM(\s$4071 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_6_88_0 (.A(\c$3744 ),
    .B(\c$3746 ),
    .CIN(\s$3749 ),
    .COUT(\c$4072 ),
    .SUM(\s$4073 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_6_89_0 (.A(\c$3748 ),
    .B(\c$3750 ),
    .CIN(\s$3753 ),
    .COUT(\c$4074 ),
    .SUM(\s$4075 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_8_0 (.A(\c$3424 ),
    .B(\c$3426 ),
    .CIN(\s$3429 ),
    .COUT(\c$3912 ),
    .SUM(\s$3913 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_6_90_0 (.A(\c$3752 ),
    .B(\c$3754 ),
    .CIN(\s$3757 ),
    .COUT(\c$4076 ),
    .SUM(\s$4077 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_91_0 (.A(\c$3756 ),
    .B(\c$3758 ),
    .CIN(\s$3761 ),
    .COUT(\c$4078 ),
    .SUM(\s$4079 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_92_0 (.A(\c$3760 ),
    .B(\c$3762 ),
    .CIN(\s$3765 ),
    .COUT(\c$4080 ),
    .SUM(\s$4081 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_93_0 (.A(\c$3764 ),
    .B(\c$3766 ),
    .CIN(\s$3769 ),
    .COUT(\c$4082 ),
    .SUM(\s$4083 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_94_0 (.A(\c$3768 ),
    .B(\c$3770 ),
    .CIN(\s$3773 ),
    .COUT(\c$4084 ),
    .SUM(\s$4085 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_95_0 (.A(\c$3772 ),
    .B(\c$3774 ),
    .CIN(\s$3777 ),
    .COUT(\c$4086 ),
    .SUM(\s$4087 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_96_0 (.A(\c$3776 ),
    .B(\c$3778 ),
    .CIN(\s$3781 ),
    .COUT(\c$4088 ),
    .SUM(\s$4089 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_97_0 (.A(\c$3780 ),
    .B(\c$3782 ),
    .CIN(\s$3785 ),
    .COUT(\c$4090 ),
    .SUM(\s$4091 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_98_0 (.A(\c$3784 ),
    .B(\c$3786 ),
    .CIN(\s$3789 ),
    .COUT(\c$4092 ),
    .SUM(\s$4093 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_99_0 (.A(\c$3788 ),
    .B(\c$3790 ),
    .CIN(\s$3793 ),
    .COUT(\c$4094 ),
    .SUM(\s$4095 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_6_9_0 (.A(\c$3428 ),
    .B(\c$3430 ),
    .CIN(\s$3433 ),
    .COUT(\c$3914 ),
    .SUM(\s$3915 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_100_0 (.A(\s$3799 ),
    .B(\c$4094 ),
    .CIN(\s$4097 ),
    .COUT(\c$4352 ),
    .SUM(\s$4353 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_101_0 (.A(\s$3803 ),
    .B(\c$4096 ),
    .CIN(\s$4099 ),
    .COUT(\c$4354 ),
    .SUM(\s$4355 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_102_0 (.A(\s$3807 ),
    .B(\c$4098 ),
    .CIN(\s$4101 ),
    .COUT(\c$4356 ),
    .SUM(\s$4357 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_103_0 (.A(\s$3811 ),
    .B(\c$4100 ),
    .CIN(\s$4103 ),
    .COUT(\c$4358 ),
    .SUM(\s$4359 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_104_0 (.A(\s$3815 ),
    .B(\c$4102 ),
    .CIN(\s$4105 ),
    .COUT(\c$4360 ),
    .SUM(\s$4361 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_105_0 (.A(\s$3819 ),
    .B(\c$4104 ),
    .CIN(\s$4107 ),
    .COUT(\c$4362 ),
    .SUM(\s$4363 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_106_0 (.A(\s$3823 ),
    .B(\c$4106 ),
    .CIN(\s$4109 ),
    .COUT(\c$4364 ),
    .SUM(\s$4365 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_107_0 (.A(\s$3827 ),
    .B(\c$4108 ),
    .CIN(\s$4111 ),
    .COUT(\c$4366 ),
    .SUM(\s$4367 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_108_0 (.A(\s$3831 ),
    .B(\c$4110 ),
    .CIN(\s$4113 ),
    .COUT(\c$4368 ),
    .SUM(\s$4369 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_109_0 (.A(\s$3835 ),
    .B(\c$4112 ),
    .CIN(\s$4115 ),
    .COUT(\c$4370 ),
    .SUM(\s$4371 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_10_0 (.A(\s$3439 ),
    .B(\c$3914 ),
    .CIN(\s$3917 ),
    .COUT(\c$4172 ),
    .SUM(\s$4173 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_110_0 (.A(\s$3839 ),
    .B(\c$4114 ),
    .CIN(\s$4117 ),
    .COUT(\c$4372 ),
    .SUM(\s$4373 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_111_0 (.A(\s$3843 ),
    .B(\c$4116 ),
    .CIN(\s$4119 ),
    .COUT(\c$4374 ),
    .SUM(\s$4375 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_112_0 (.A(\s$3847 ),
    .B(\c$4118 ),
    .CIN(\s$4121 ),
    .COUT(\c$4376 ),
    .SUM(\s$4377 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_113_0 (.A(\s$3851 ),
    .B(\c$4120 ),
    .CIN(\s$4123 ),
    .COUT(\c$4378 ),
    .SUM(\s$4379 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_114_0 (.A(\s$3855 ),
    .B(\c$4122 ),
    .CIN(\s$4125 ),
    .COUT(\c$4380 ),
    .SUM(\s$4381 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_115_0 (.A(\s$3859 ),
    .B(\c$4124 ),
    .CIN(\s$4127 ),
    .COUT(\c$4382 ),
    .SUM(\s$4383 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_116_0 (.A(\s$3863 ),
    .B(\c$4126 ),
    .CIN(\s$4129 ),
    .COUT(\c$4384 ),
    .SUM(\s$4385 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_117_0 (.A(\s$3867 ),
    .B(\c$4128 ),
    .CIN(\s$4131 ),
    .COUT(\c$4386 ),
    .SUM(\s$4387 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_118_0 (.A(\s$3871 ),
    .B(\c$4130 ),
    .CIN(\s$4133 ),
    .COUT(\c$4388 ),
    .SUM(\s$4389 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_119_0 (.A(\s$3875 ),
    .B(\c$4132 ),
    .CIN(\s$4135 ),
    .COUT(\c$4390 ),
    .SUM(\s$4391 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_11_0 (.A(\s$3443 ),
    .B(\c$3916 ),
    .CIN(\s$3919 ),
    .COUT(\c$4174 ),
    .SUM(\s$4175 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_120_0 (.A(\s$3879 ),
    .B(\c$4134 ),
    .CIN(\s$4137 ),
    .COUT(\c$4392 ),
    .SUM(\s$4393 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_121_0 (.A(\s$3883 ),
    .B(\c$4136 ),
    .CIN(\s$4139 ),
    .COUT(\c$4394 ),
    .SUM(\s$4395 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_122_0 (.A(\s$3887 ),
    .B(\c$4138 ),
    .CIN(\s$4141 ),
    .COUT(\c$4396 ),
    .SUM(\s$4397 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_123_0 (.A(\s$3891 ),
    .B(\c$4140 ),
    .CIN(\s$4143 ),
    .COUT(\c$4398 ),
    .SUM(\s$4399 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_124_0 (.A(\s$3895 ),
    .B(\c$4142 ),
    .CIN(\s$4145 ),
    .COUT(\c$4400 ),
    .SUM(\s$4401 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_125_0 (.A(\s$3897 ),
    .B(\c$4144 ),
    .CIN(\s$4147 ),
    .COUT(\c$4402 ),
    .SUM(\s$4403 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_126_0 (.A(\s$3899 ),
    .B(\c$4146 ),
    .CIN(\s$4149 ),
    .COUT(\c$4404 ),
    .SUM(\s$4405 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_127_0 (.A(\c$3898 ),
    .B(\c$4148 ),
    .CIN(\s$4151 ),
    .COUT(\c$4406 ),
    .SUM(\s$4407 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_12_0 (.A(\s$3447 ),
    .B(\c$3918 ),
    .CIN(\s$3921 ),
    .COUT(\c$4176 ),
    .SUM(\s$4177 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_13_0 (.A(\s$3451 ),
    .B(\c$3920 ),
    .CIN(\s$3923 ),
    .COUT(\c$4178 ),
    .SUM(\s$4179 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_14_0 (.A(\s$3455 ),
    .B(\c$3922 ),
    .CIN(\s$3925 ),
    .COUT(\c$4180 ),
    .SUM(\s$4181 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_15_0 (.A(\s$3459 ),
    .B(\c$3924 ),
    .CIN(\s$3927 ),
    .COUT(\c$4182 ),
    .SUM(\s$4183 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_16_0 (.A(\s$3463 ),
    .B(\c$3926 ),
    .CIN(\s$3929 ),
    .COUT(\c$4184 ),
    .SUM(\s$4185 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_17_0 (.A(\s$3467 ),
    .B(\c$3928 ),
    .CIN(\s$3931 ),
    .COUT(\c$4186 ),
    .SUM(\s$4187 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_18_0 (.A(\s$3471 ),
    .B(\c$3930 ),
    .CIN(\s$3933 ),
    .COUT(\c$4188 ),
    .SUM(\s$4189 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_19_0 (.A(\s$3475 ),
    .B(\c$3932 ),
    .CIN(\s$3935 ),
    .COUT(\c$4190 ),
    .SUM(\s$4191 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_20_0 (.A(\s$3479 ),
    .B(\c$3934 ),
    .CIN(\s$3937 ),
    .COUT(\c$4192 ),
    .SUM(\s$4193 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_21_0 (.A(\s$3483 ),
    .B(\c$3936 ),
    .CIN(\s$3939 ),
    .COUT(\c$4194 ),
    .SUM(\s$4195 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_22_0 (.A(\s$3487 ),
    .B(\c$3938 ),
    .CIN(\s$3941 ),
    .COUT(\c$4196 ),
    .SUM(\s$4197 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_23_0 (.A(\s$3491 ),
    .B(\c$3940 ),
    .CIN(\s$3943 ),
    .COUT(\c$4198 ),
    .SUM(\s$4199 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_24_0 (.A(\s$3495 ),
    .B(\c$3942 ),
    .CIN(\s$3945 ),
    .COUT(\c$4200 ),
    .SUM(\s$4201 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_25_0 (.A(\s$3499 ),
    .B(\c$3944 ),
    .CIN(\s$3947 ),
    .COUT(\c$4202 ),
    .SUM(\s$4203 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_26_0 (.A(\s$3503 ),
    .B(\c$3946 ),
    .CIN(\s$3949 ),
    .COUT(\c$4204 ),
    .SUM(\s$4205 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_27_0 (.A(\s$3507 ),
    .B(\c$3948 ),
    .CIN(\s$3951 ),
    .COUT(\c$4206 ),
    .SUM(\s$4207 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_28_0 (.A(\s$3511 ),
    .B(\c$3950 ),
    .CIN(\s$3953 ),
    .COUT(\c$4208 ),
    .SUM(\s$4209 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_29_0 (.A(\s$3515 ),
    .B(\c$3952 ),
    .CIN(\s$3955 ),
    .COUT(\c$4210 ),
    .SUM(\s$4211 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_2_0 (.A(pp_row2_2),
    .B(pp_row2_3),
    .CIN(\s$3901 ),
    .COUT(\c$4156 ),
    .SUM(\s$4157 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_30_0 (.A(\s$3519 ),
    .B(\c$3954 ),
    .CIN(\s$3957 ),
    .COUT(\c$4212 ),
    .SUM(\s$4213 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_31_0 (.A(\s$3523 ),
    .B(\c$3956 ),
    .CIN(\s$3959 ),
    .COUT(\c$4214 ),
    .SUM(\s$4215 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_32_0 (.A(\s$3527 ),
    .B(\c$3958 ),
    .CIN(\s$3961 ),
    .COUT(\c$4216 ),
    .SUM(\s$4217 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_33_0 (.A(\s$3531 ),
    .B(\c$3960 ),
    .CIN(\s$3963 ),
    .COUT(\c$4218 ),
    .SUM(\s$4219 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_34_0 (.A(\s$3535 ),
    .B(\c$3962 ),
    .CIN(\s$3965 ),
    .COUT(\c$4220 ),
    .SUM(\s$4221 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_35_0 (.A(\s$3539 ),
    .B(\c$3964 ),
    .CIN(\s$3967 ),
    .COUT(\c$4222 ),
    .SUM(\s$4223 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_36_0 (.A(\s$3543 ),
    .B(\c$3966 ),
    .CIN(\s$3969 ),
    .COUT(\c$4224 ),
    .SUM(\s$4225 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_37_0 (.A(\s$3547 ),
    .B(\c$3968 ),
    .CIN(\s$3971 ),
    .COUT(\c$4226 ),
    .SUM(\s$4227 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_38_0 (.A(\s$3551 ),
    .B(\c$3970 ),
    .CIN(\s$3973 ),
    .COUT(\c$4228 ),
    .SUM(\s$4229 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_39_0 (.A(\s$3555 ),
    .B(\c$3972 ),
    .CIN(\s$3975 ),
    .COUT(\c$4230 ),
    .SUM(\s$4231 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_3_0 (.A(pp_row3_2),
    .B(\c$3900 ),
    .CIN(\s$3903 ),
    .COUT(\c$4158 ),
    .SUM(\s$4159 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_40_0 (.A(\s$3559 ),
    .B(\c$3974 ),
    .CIN(\s$3977 ),
    .COUT(\c$4232 ),
    .SUM(\s$4233 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_41_0 (.A(\s$3563 ),
    .B(\c$3976 ),
    .CIN(\s$3979 ),
    .COUT(\c$4234 ),
    .SUM(\s$4235 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_42_0 (.A(\s$3567 ),
    .B(\c$3978 ),
    .CIN(\s$3981 ),
    .COUT(\c$4236 ),
    .SUM(\s$4237 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_43_0 (.A(\s$3571 ),
    .B(\c$3980 ),
    .CIN(\s$3983 ),
    .COUT(\c$4238 ),
    .SUM(\s$4239 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_44_0 (.A(\s$3575 ),
    .B(\c$3982 ),
    .CIN(\s$3985 ),
    .COUT(\c$4240 ),
    .SUM(\s$4241 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_45_0 (.A(\s$3579 ),
    .B(\c$3984 ),
    .CIN(\s$3987 ),
    .COUT(\c$4242 ),
    .SUM(\s$4243 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_46_0 (.A(\s$3583 ),
    .B(\c$3986 ),
    .CIN(\s$3989 ),
    .COUT(\c$4244 ),
    .SUM(\s$4245 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_47_0 (.A(\s$3587 ),
    .B(\c$3988 ),
    .CIN(\s$3991 ),
    .COUT(\c$4246 ),
    .SUM(\s$4247 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_48_0 (.A(\s$3591 ),
    .B(\c$3990 ),
    .CIN(\s$3993 ),
    .COUT(\c$4248 ),
    .SUM(\s$4249 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_49_0 (.A(\s$3595 ),
    .B(\c$3992 ),
    .CIN(\s$3995 ),
    .COUT(\c$4250 ),
    .SUM(\s$4251 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_4_0 (.A(\s$3417 ),
    .B(\c$3902 ),
    .CIN(\s$3905 ),
    .COUT(\c$4160 ),
    .SUM(\s$4161 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_50_0 (.A(\s$3599 ),
    .B(\c$3994 ),
    .CIN(\s$3997 ),
    .COUT(\c$4252 ),
    .SUM(\s$4253 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_51_0 (.A(\s$3603 ),
    .B(\c$3996 ),
    .CIN(\s$3999 ),
    .COUT(\c$4254 ),
    .SUM(\s$4255 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_52_0 (.A(\s$3607 ),
    .B(\c$3998 ),
    .CIN(\s$4001 ),
    .COUT(\c$4256 ),
    .SUM(\s$4257 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_53_0 (.A(\s$3611 ),
    .B(\c$4000 ),
    .CIN(\s$4003 ),
    .COUT(\c$4258 ),
    .SUM(\s$4259 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_54_0 (.A(\s$3615 ),
    .B(\c$4002 ),
    .CIN(\s$4005 ),
    .COUT(\c$4260 ),
    .SUM(\s$4261 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_55_0 (.A(\s$3619 ),
    .B(\c$4004 ),
    .CIN(\s$4007 ),
    .COUT(\c$4262 ),
    .SUM(\s$4263 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_56_0 (.A(\s$3623 ),
    .B(\c$4006 ),
    .CIN(\s$4009 ),
    .COUT(\c$4264 ),
    .SUM(\s$4265 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_57_0 (.A(\s$3627 ),
    .B(\c$4008 ),
    .CIN(\s$4011 ),
    .COUT(\c$4266 ),
    .SUM(\s$4267 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_58_0 (.A(\s$3631 ),
    .B(\c$4010 ),
    .CIN(\s$4013 ),
    .COUT(\c$4268 ),
    .SUM(\s$4269 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_59_0 (.A(\s$3635 ),
    .B(\c$4012 ),
    .CIN(\s$4015 ),
    .COUT(\c$4270 ),
    .SUM(\s$4271 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_5_0 (.A(\s$3419 ),
    .B(\c$3904 ),
    .CIN(\s$3907 ),
    .COUT(\c$4162 ),
    .SUM(\s$4163 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_60_0 (.A(\s$3639 ),
    .B(\c$4014 ),
    .CIN(\s$4017 ),
    .COUT(\c$4272 ),
    .SUM(\s$4273 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_61_0 (.A(\s$3643 ),
    .B(\c$4016 ),
    .CIN(\s$4019 ),
    .COUT(\c$4274 ),
    .SUM(\s$4275 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_62_0 (.A(\s$3647 ),
    .B(\c$4018 ),
    .CIN(\s$4021 ),
    .COUT(\c$4276 ),
    .SUM(\s$4277 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_63_0 (.A(\s$3651 ),
    .B(\c$4020 ),
    .CIN(\s$4023 ),
    .COUT(\c$4278 ),
    .SUM(\s$4279 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_64_0 (.A(\s$3655 ),
    .B(\c$4022 ),
    .CIN(\s$4025 ),
    .COUT(\c$4280 ),
    .SUM(\s$4281 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_65_0 (.A(\s$3659 ),
    .B(\c$4024 ),
    .CIN(\s$4027 ),
    .COUT(\c$4282 ),
    .SUM(\s$4283 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_66_0 (.A(\s$3663 ),
    .B(\c$4026 ),
    .CIN(\s$4029 ),
    .COUT(\c$4284 ),
    .SUM(\s$4285 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_67_0 (.A(\s$3667 ),
    .B(\c$4028 ),
    .CIN(\s$4031 ),
    .COUT(\c$4286 ),
    .SUM(\s$4287 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_68_0 (.A(\s$3671 ),
    .B(\c$4030 ),
    .CIN(\s$4033 ),
    .COUT(\c$4288 ),
    .SUM(\s$4289 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_69_0 (.A(\s$3675 ),
    .B(\c$4032 ),
    .CIN(\s$4035 ),
    .COUT(\c$4290 ),
    .SUM(\s$4291 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_6_0 (.A(\s$3423 ),
    .B(\c$3906 ),
    .CIN(\s$3909 ),
    .COUT(\c$4164 ),
    .SUM(\s$4165 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_70_0 (.A(\s$3679 ),
    .B(\c$4034 ),
    .CIN(\s$4037 ),
    .COUT(\c$4292 ),
    .SUM(\s$4293 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_71_0 (.A(\s$3683 ),
    .B(\c$4036 ),
    .CIN(\s$4039 ),
    .COUT(\c$4294 ),
    .SUM(\s$4295 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_72_0 (.A(\s$3687 ),
    .B(\c$4038 ),
    .CIN(\s$4041 ),
    .COUT(\c$4296 ),
    .SUM(\s$4297 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_73_0 (.A(\s$3691 ),
    .B(\c$4040 ),
    .CIN(\s$4043 ),
    .COUT(\c$4298 ),
    .SUM(\s$4299 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_74_0 (.A(\s$3695 ),
    .B(\c$4042 ),
    .CIN(\s$4045 ),
    .COUT(\c$4300 ),
    .SUM(\s$4301 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_75_0 (.A(\s$3699 ),
    .B(\c$4044 ),
    .CIN(\s$4047 ),
    .COUT(\c$4302 ),
    .SUM(\s$4303 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_76_0 (.A(\s$3703 ),
    .B(\c$4046 ),
    .CIN(\s$4049 ),
    .COUT(\c$4304 ),
    .SUM(\s$4305 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_77_0 (.A(\s$3707 ),
    .B(\c$4048 ),
    .CIN(\s$4051 ),
    .COUT(\c$4306 ),
    .SUM(\s$4307 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_78_0 (.A(\s$3711 ),
    .B(\c$4050 ),
    .CIN(\s$4053 ),
    .COUT(\c$4308 ),
    .SUM(\s$4309 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_79_0 (.A(\s$3715 ),
    .B(\c$4052 ),
    .CIN(\s$4055 ),
    .COUT(\c$4310 ),
    .SUM(\s$4311 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_7_0 (.A(\s$3427 ),
    .B(\c$3908 ),
    .CIN(\s$3911 ),
    .COUT(\c$4166 ),
    .SUM(\s$4167 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_80_0 (.A(\s$3719 ),
    .B(\c$4054 ),
    .CIN(\s$4057 ),
    .COUT(\c$4312 ),
    .SUM(\s$4313 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_81_0 (.A(\s$3723 ),
    .B(\c$4056 ),
    .CIN(\s$4059 ),
    .COUT(\c$4314 ),
    .SUM(\s$4315 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_82_0 (.A(\s$3727 ),
    .B(\c$4058 ),
    .CIN(\s$4061 ),
    .COUT(\c$4316 ),
    .SUM(\s$4317 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_83_0 (.A(\s$3731 ),
    .B(\c$4060 ),
    .CIN(\s$4063 ),
    .COUT(\c$4318 ),
    .SUM(\s$4319 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_84_0 (.A(\s$3735 ),
    .B(\c$4062 ),
    .CIN(\s$4065 ),
    .COUT(\c$4320 ),
    .SUM(\s$4321 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_85_0 (.A(\s$3739 ),
    .B(\c$4064 ),
    .CIN(\s$4067 ),
    .COUT(\c$4322 ),
    .SUM(\s$4323 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_86_0 (.A(\s$3743 ),
    .B(\c$4066 ),
    .CIN(\s$4069 ),
    .COUT(\c$4324 ),
    .SUM(\s$4325 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_87_0 (.A(\s$3747 ),
    .B(\c$4068 ),
    .CIN(\s$4071 ),
    .COUT(\c$4326 ),
    .SUM(\s$4327 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_88_0 (.A(\s$3751 ),
    .B(\c$4070 ),
    .CIN(\s$4073 ),
    .COUT(\c$4328 ),
    .SUM(\s$4329 ));
 sky130_fd_sc_hd__fa_2 dadda_fa_7_89_0 (.A(\s$3755 ),
    .B(\c$4072 ),
    .CIN(\s$4075 ),
    .COUT(\c$4330 ),
    .SUM(\s$4331 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_8_0 (.A(\s$3431 ),
    .B(\c$3910 ),
    .CIN(\s$3913 ),
    .COUT(\c$4168 ),
    .SUM(\s$4169 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_90_0 (.A(\s$3759 ),
    .B(\c$4074 ),
    .CIN(\s$4077 ),
    .COUT(\c$4332 ),
    .SUM(\s$4333 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_91_0 (.A(\s$3763 ),
    .B(\c$4076 ),
    .CIN(\s$4079 ),
    .COUT(\c$4334 ),
    .SUM(\s$4335 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_92_0 (.A(\s$3767 ),
    .B(\c$4078 ),
    .CIN(\s$4081 ),
    .COUT(\c$4336 ),
    .SUM(\s$4337 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_93_0 (.A(\s$3771 ),
    .B(\c$4080 ),
    .CIN(\s$4083 ),
    .COUT(\c$4338 ),
    .SUM(\s$4339 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_94_0 (.A(\s$3775 ),
    .B(\c$4082 ),
    .CIN(\s$4085 ),
    .COUT(\c$4340 ),
    .SUM(\s$4341 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_95_0 (.A(\s$3779 ),
    .B(\c$4084 ),
    .CIN(\s$4087 ),
    .COUT(\c$4342 ),
    .SUM(\s$4343 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_96_0 (.A(\s$3783 ),
    .B(\c$4086 ),
    .CIN(\s$4089 ),
    .COUT(\c$4344 ),
    .SUM(\s$4345 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_97_0 (.A(\s$3787 ),
    .B(\c$4088 ),
    .CIN(\s$4091 ),
    .COUT(\c$4346 ),
    .SUM(\s$4347 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_98_0 (.A(\s$3791 ),
    .B(\c$4090 ),
    .CIN(\s$4093 ),
    .COUT(\c$4348 ),
    .SUM(\s$4349 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_99_0 (.A(\s$3795 ),
    .B(\c$4092 ),
    .CIN(\s$4095 ),
    .COUT(\c$4350 ),
    .SUM(\s$4351 ));
 sky130_fd_sc_hd__fa_1 dadda_fa_7_9_0 (.A(\s$3435 ),
    .B(\c$3912 ),
    .CIN(\s$3915 ),
    .COUT(\c$4170 ),
    .SUM(\s$4171 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_52_0 (.A(pp_row52_0),
    .B(pp_row52_1),
    .COUT(\c$1 ),
    .SUM(s));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_53_0 (.A(pp_row53_0),
    .B(pp_row53_1),
    .COUT(\c$2 ),
    .SUM(\s$3 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_54_1 (.A(pp_row54_3),
    .B(pp_row54_4),
    .COUT(\c$6 ),
    .SUM(\s$7 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_55_1 (.A(pp_row55_3),
    .B(pp_row55_4),
    .COUT(\c$10 ),
    .SUM(\s$11 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_56_2 (.A(pp_row56_6),
    .B(pp_row56_7),
    .COUT(\c$16 ),
    .SUM(\s$17 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_57_2 (.A(pp_row57_6),
    .B(pp_row57_7),
    .COUT(\c$22 ),
    .SUM(\s$23 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_58_3 (.A(pp_row58_9),
    .B(pp_row58_10),
    .COUT(\c$30 ),
    .SUM(\s$31 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_59_3 (.A(pp_row59_9),
    .B(pp_row59_10),
    .COUT(\c$38 ),
    .SUM(\s$39 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_60_4 (.A(pp_row60_12),
    .B(pp_row60_13),
    .COUT(\c$48 ),
    .SUM(\s$49 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_61_4 (.A(pp_row61_12),
    .B(pp_row61_13),
    .COUT(\c$58 ),
    .SUM(\s$59 ));
 sky130_fd_sc_hd__ha_2 dadda_ha_0_62_5 (.A(pp_row62_15),
    .B(pp_row62_16),
    .COUT(\c$70 ),
    .SUM(\s$71 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_63_5 (.A(pp_row63_15),
    .B(pp_row63_16),
    .COUT(\c$82 ),
    .SUM(\s$83 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_68_5 (.A(pp_row68_15),
    .B(pp_row68_16),
    .COUT(\c$142 ),
    .SUM(\s$143 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_70_4 (.A(pp_row70_12),
    .B(pp_row70_13),
    .COUT(\c$162 ),
    .SUM(\s$163 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_72_3 (.A(pp_row72_9),
    .B(pp_row72_10),
    .COUT(\c$178 ),
    .SUM(\s$179 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_74_2 (.A(pp_row74_6),
    .B(pp_row74_7),
    .COUT(\c$190 ),
    .SUM(\s$191 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_76_1 (.A(pp_row76_3),
    .B(pp_row76_4),
    .COUT(\c$198 ),
    .SUM(\s$199 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_0_78_0 (.A(net1915),
    .B(pp_row78_1),
    .COUT(\c$202 ),
    .SUM(\s$203 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_34_0 (.A(pp_row34_0),
    .B(pp_row34_1),
    .COUT(\c$204 ),
    .SUM(\s$205 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_35_0 (.A(pp_row35_0),
    .B(pp_row35_1),
    .COUT(\c$206 ),
    .SUM(\s$207 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_36_1 (.A(pp_row36_3),
    .B(pp_row36_4),
    .COUT(\c$210 ),
    .SUM(\s$211 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_37_1 (.A(pp_row37_3),
    .B(pp_row37_4),
    .COUT(\c$214 ),
    .SUM(\s$215 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_38_2 (.A(pp_row38_6),
    .B(pp_row38_7),
    .COUT(\c$220 ),
    .SUM(\s$221 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_39_2 (.A(pp_row39_6),
    .B(pp_row39_7),
    .COUT(\c$226 ),
    .SUM(\s$227 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_40_3 (.A(pp_row40_9),
    .B(pp_row40_10),
    .COUT(\c$234 ),
    .SUM(\s$235 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_41_3 (.A(pp_row41_9),
    .B(pp_row41_10),
    .COUT(\c$242 ),
    .SUM(\s$243 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_42_4 (.A(pp_row42_12),
    .B(pp_row42_13),
    .COUT(\c$252 ),
    .SUM(\s$253 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_43_4 (.A(pp_row43_12),
    .B(pp_row43_13),
    .COUT(\c$262 ),
    .SUM(\s$263 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_44_5 (.A(pp_row44_15),
    .B(pp_row44_16),
    .COUT(\c$274 ),
    .SUM(\s$275 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_45_5 (.A(pp_row45_15),
    .B(pp_row45_16),
    .COUT(\c$286 ),
    .SUM(\s$287 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_46_6 (.A(pp_row46_18),
    .B(pp_row46_19),
    .COUT(\c$300 ),
    .SUM(\s$301 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_47_6 (.A(pp_row47_18),
    .B(pp_row47_19),
    .COUT(\c$314 ),
    .SUM(\s$315 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_48_7 (.A(pp_row48_21),
    .B(pp_row48_22),
    .COUT(\c$330 ),
    .SUM(\s$331 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_49_7 (.A(pp_row49_21),
    .B(pp_row49_22),
    .COUT(\c$346 ),
    .SUM(\s$347 ));
 sky130_fd_sc_hd__ha_2 dadda_ha_1_50_8 (.A(pp_row50_24),
    .B(pp_row50_25),
    .COUT(\c$364 ),
    .SUM(\s$365 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_51_8 (.A(pp_row51_24),
    .B(pp_row51_25),
    .COUT(\c$382 ),
    .SUM(\s$383 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_80_8 (.A(pp_row80_24),
    .B(pp_row80_25),
    .COUT(\c$904 ),
    .SUM(\s$905 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_82_7 (.A(pp_row82_21),
    .B(pp_row82_22),
    .COUT(\c$936 ),
    .SUM(\s$937 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_84_6 (.A(pp_row84_18),
    .B(pp_row84_19),
    .COUT(\c$964 ),
    .SUM(\s$965 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_86_5 (.A(pp_row86_15),
    .B(pp_row86_16),
    .COUT(\c$988 ),
    .SUM(\s$989 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_88_4 (.A(pp_row88_12),
    .B(pp_row88_13),
    .COUT(\c$1008 ),
    .SUM(\s$1009 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_90_3 (.A(pp_row90_9),
    .B(pp_row90_10),
    .COUT(\c$1024 ),
    .SUM(\s$1025 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_92_2 (.A(pp_row92_6),
    .B(pp_row92_7),
    .COUT(\c$1036 ),
    .SUM(\s$1037 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_94_1 (.A(pp_row94_3),
    .B(pp_row94_4),
    .COUT(\c$1044 ),
    .SUM(\s$1045 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_1_96_0 (.A(net1916),
    .B(pp_row96_1),
    .COUT(\c$1048 ),
    .SUM(\s$1049 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_100_4 (.A(pp_row100_12),
    .B(pp_row100_13),
    .COUT(\c$1932 ),
    .SUM(\s$1933 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_102_3 (.A(pp_row102_9),
    .B(pp_row102_10),
    .COUT(\c$1948 ),
    .SUM(\s$1949 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_104_2 (.A(pp_row104_6),
    .B(pp_row104_7),
    .COUT(\c$1960 ),
    .SUM(\s$1961 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_106_1 (.A(pp_row106_3),
    .B(pp_row106_4),
    .COUT(\c$1968 ),
    .SUM(\s$1969 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_108_0 (.A(net1917),
    .B(pp_row108_1),
    .COUT(\c$1972 ),
    .SUM(\s$1973 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_22_0 (.A(pp_row22_0),
    .B(pp_row22_1),
    .COUT(\c$1050 ),
    .SUM(\s$1051 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_23_0 (.A(pp_row23_0),
    .B(pp_row23_1),
    .COUT(\c$1052 ),
    .SUM(\s$1053 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_24_1 (.A(pp_row24_3),
    .B(pp_row24_4),
    .COUT(\c$1056 ),
    .SUM(\s$1057 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_25_1 (.A(pp_row25_3),
    .B(pp_row25_4),
    .COUT(\c$1060 ),
    .SUM(\s$1061 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_26_2 (.A(pp_row26_6),
    .B(pp_row26_7),
    .COUT(\c$1066 ),
    .SUM(\s$1067 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_27_2 (.A(pp_row27_6),
    .B(pp_row27_7),
    .COUT(\c$1072 ),
    .SUM(\s$1073 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_28_3 (.A(pp_row28_9),
    .B(pp_row28_10),
    .COUT(\c$1080 ),
    .SUM(\s$1081 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_29_3 (.A(pp_row29_9),
    .B(pp_row29_10),
    .COUT(\c$1088 ),
    .SUM(\s$1089 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_30_4 (.A(pp_row30_12),
    .B(pp_row30_13),
    .COUT(\c$1098 ),
    .SUM(\s$1099 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_31_4 (.A(pp_row31_12),
    .B(pp_row31_13),
    .COUT(\c$1108 ),
    .SUM(\s$1109 ));
 sky130_fd_sc_hd__ha_2 dadda_ha_2_32_5 (.A(pp_row32_15),
    .B(pp_row32_16),
    .COUT(\c$1120 ),
    .SUM(\s$1121 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_33_5 (.A(pp_row33_15),
    .B(pp_row33_16),
    .COUT(\c$1132 ),
    .SUM(\s$1133 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_2_98_5 (.A(pp_row98_15),
    .B(pp_row98_16),
    .COUT(\c$1912 ),
    .SUM(\s$1913 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_3_110_3 (.A(pp_row110_9),
    .B(pp_row110_10),
    .COUT(\c$2724 ),
    .SUM(\s$2725 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_3_112_2 (.A(pp_row112_6),
    .B(pp_row112_7),
    .COUT(\c$2736 ),
    .SUM(\s$2737 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_3_114_1 (.A(pp_row114_3),
    .B(pp_row114_4),
    .COUT(\c$2744 ),
    .SUM(\s$2745 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_3_116_0 (.A(net1918),
    .B(pp_row116_1),
    .COUT(\c$2748 ),
    .SUM(\s$2749 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_3_14_0 (.A(pp_row14_0),
    .B(pp_row14_1),
    .COUT(\c$1974 ),
    .SUM(\s$1975 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_3_15_0 (.A(pp_row15_0),
    .B(pp_row15_1),
    .COUT(\c$1976 ),
    .SUM(\s$1977 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_3_16_1 (.A(pp_row16_3),
    .B(pp_row16_4),
    .COUT(\c$1980 ),
    .SUM(\s$1981 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_3_17_1 (.A(pp_row17_3),
    .B(pp_row17_4),
    .COUT(\c$1984 ),
    .SUM(\s$1985 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_3_18_2 (.A(pp_row18_6),
    .B(pp_row18_7),
    .COUT(\c$1990 ),
    .SUM(\s$1991 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_3_19_2 (.A(pp_row19_6),
    .B(pp_row19_7),
    .COUT(\c$1996 ),
    .SUM(\s$1997 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_3_20_3 (.A(pp_row20_9),
    .B(pp_row20_10),
    .COUT(\c$2004 ),
    .SUM(\s$2005 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_3_21_3 (.A(pp_row21_9),
    .B(pp_row21_10),
    .COUT(\c$2012 ),
    .SUM(\s$2013 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_4_10_1 (.A(pp_row10_3),
    .B(pp_row10_4),
    .COUT(\c$2756 ),
    .SUM(\s$2757 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_4_118_2 (.A(pp_row118_6),
    .B(pp_row118_7),
    .COUT(\c$3402 ),
    .SUM(\s$3403 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_4_11_1 (.A(pp_row11_3),
    .B(pp_row11_4),
    .COUT(\c$2760 ),
    .SUM(\s$2761 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_4_120_1 (.A(pp_row120_3),
    .B(pp_row120_4),
    .COUT(\c$3410 ),
    .SUM(\s$3411 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_4_122_0 (.A(net1919),
    .B(pp_row122_1),
    .COUT(\c$3414 ),
    .SUM(\s$3415 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_4_12_2 (.A(pp_row12_6),
    .B(pp_row12_7),
    .COUT(\c$2766 ),
    .SUM(\s$2767 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_4_13_2 (.A(pp_row13_6),
    .B(pp_row13_7),
    .COUT(\c$2772 ),
    .SUM(\s$2773 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_4_8_0 (.A(pp_row8_0),
    .B(pp_row8_1),
    .COUT(\c$2750 ),
    .SUM(\s$2751 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_4_9_0 (.A(pp_row9_0),
    .B(pp_row9_1),
    .COUT(\c$2752 ),
    .SUM(\s$2753 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_5_124_1 (.A(pp_row124_3),
    .B(pp_row124_4),
    .COUT(\c$3894 ),
    .SUM(\s$3895 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_5_126_0 (.A(net1920),
    .B(pp_row126_1),
    .COUT(\c$3898 ),
    .SUM(\s$3899 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_5_4_0 (.A(pp_row4_0),
    .B(pp_row4_1),
    .COUT(\c$3416 ),
    .SUM(\s$3417 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_5_5_0 (.A(pp_row5_0),
    .B(pp_row5_1),
    .COUT(\c$3418 ),
    .SUM(\s$3419 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_5_6_1 (.A(pp_row6_3),
    .B(pp_row6_4),
    .COUT(\c$3422 ),
    .SUM(\s$3423 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_5_7_1 (.A(pp_row7_3),
    .B(pp_row7_4),
    .COUT(\c$3426 ),
    .SUM(\s$3427 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_6_2_0 (.A(pp_row2_0),
    .B(pp_row2_1),
    .COUT(\c$3900 ),
    .SUM(\s$3901 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_6_3_0 (.A(pp_row3_0),
    .B(pp_row3_1),
    .COUT(\c$3902 ),
    .SUM(\s$3903 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_7_0_0 (.A(pp_row0_0),
    .B(pp_row0_1),
    .COUT(\c$4152 ),
    .SUM(\s$4153 ));
 sky130_fd_sc_hd__ha_1 dadda_ha_7_1_0 (.A(pp_row1_0),
    .B(pp_row1_1),
    .COUT(\c$4154 ),
    .SUM(\s$4155 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$0  (.A(pp_row0_2),
    .B(\s$4153 ),
    .COUT(\final_adder.$signal ),
    .SUM(\final_adder.$signal$1 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$1  (.A(\c$4152 ),
    .B(\s$4155 ),
    .COUT(\final_adder.$signal$4 ),
    .SUM(\final_adder.$signal$1091 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$10  (.A(\c$4170 ),
    .B(\s$4173 ),
    .COUT(\final_adder.$signal$22 ),
    .SUM(\final_adder.$signal$1100 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$100  (.A(\c$4350 ),
    .B(\s$4353 ),
    .COUT(\final_adder.$signal$202 ),
    .SUM(\final_adder.$signal$1190 ));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1000  (.A(\final_adder.$signal$1129 ),
    .B(\final_adder.g_new$1070 ),
    .X(net317));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1001  (.A(\final_adder.$signal$1130 ),
    .B(\final_adder.g_new$955 ),
    .X(net319));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1002  (.A(\final_adder.$signal$1131 ),
    .B(\final_adder.g_new$1069 ),
    .X(net320));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1003  (.A(\final_adder.$signal$1132 ),
    .B(\final_adder.g_new$953 ),
    .X(net321));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1004  (.A(\final_adder.$signal$1133 ),
    .B(\final_adder.g_new$1068 ),
    .X(net322));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1005  (.A(\final_adder.$signal$1134 ),
    .B(\final_adder.g_new$951 ),
    .X(net323));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1006  (.A(\final_adder.$signal$1135 ),
    .B(\final_adder.g_new$1067 ),
    .X(net324));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1007  (.A(\final_adder.$signal$1136 ),
    .B(\final_adder.g_new$949 ),
    .X(net325));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1008  (.A(\final_adder.$signal$1137 ),
    .B(\final_adder.g_new$1066 ),
    .X(net326));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1009  (.A(\final_adder.$signal$1138 ),
    .B(\final_adder.g_new$947 ),
    .X(net327));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$101  (.A(\c$4352 ),
    .B(\s$4355 ),
    .COUT(\final_adder.$signal$204 ),
    .SUM(\final_adder.$signal$1191 ));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1010  (.A(\final_adder.$signal$101 ),
    .B(\final_adder.g_new$1065 ),
    .X(net328));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1011  (.A(\final_adder.$signal$103 ),
    .B(\final_adder.g_new$945 ),
    .X(net330));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1012  (.A(\final_adder.$signal$105 ),
    .B(\final_adder.g_new$1064 ),
    .X(net331));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1013  (.A(\final_adder.$signal$107 ),
    .B(\final_adder.g_new$943 ),
    .X(net332));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1014  (.A(\final_adder.$signal$109 ),
    .B(\final_adder.g_new$1063 ),
    .X(net333));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1015  (.A(\final_adder.$signal$111 ),
    .B(\final_adder.g_new$941 ),
    .X(net334));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1016  (.A(\final_adder.$signal$113 ),
    .B(\final_adder.g_new$1062 ),
    .X(net335));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$1017  (.A(\final_adder.$signal$1146 ),
    .B(\final_adder.g_new$939 ),
    .X(net336));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$1018  (.A(\final_adder.$signal$1147 ),
    .B(\final_adder.g_new$1061 ),
    .X(net337));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1019  (.A(\final_adder.$signal$1148 ),
    .B(\final_adder.g_new$937 ),
    .X(net338));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$102  (.A(\c$4354 ),
    .B(\s$4357 ),
    .COUT(\final_adder.$signal$206 ),
    .SUM(\final_adder.$signal$1192 ));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1020  (.A(\final_adder.$signal$1149 ),
    .B(\final_adder.g_new$1060 ),
    .X(net339));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1021  (.A(\final_adder.$signal$1150 ),
    .B(\final_adder.g_new$935 ),
    .X(net341));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1022  (.A(\final_adder.$signal$1151 ),
    .B(\final_adder.g_new$1059 ),
    .X(net342));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1023  (.A(\final_adder.$signal$1152 ),
    .B(\final_adder.g_new$933 ),
    .X(net343));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1024  (.A(\final_adder.$signal$1153 ),
    .B(\final_adder.g_new$1058 ),
    .X(net344));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1025  (.A(\final_adder.$signal$1154 ),
    .B(\final_adder.g_new$931 ),
    .X(net345));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1026  (.A(\final_adder.$signal$1155 ),
    .B(\final_adder.g_new$1057 ),
    .X(net346));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1027  (.A(\final_adder.$signal$1156 ),
    .B(\final_adder.g_new$1025 ),
    .X(net347));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1028  (.A(\final_adder.$signal$1157 ),
    .B(\final_adder.g_new$1056 ),
    .X(net348));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1029  (.A(\final_adder.$signal$1158 ),
    .B(\final_adder.g_new$1023 ),
    .X(net349));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$103  (.A(\c$4356 ),
    .B(\s$4359 ),
    .COUT(\final_adder.$signal$208 ),
    .SUM(\final_adder.$signal$1193 ));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1030  (.A(\final_adder.$signal$1159 ),
    .B(\final_adder.g_new$1055 ),
    .X(net350));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1031  (.A(\final_adder.$signal$1160 ),
    .B(\final_adder.g_new$1021 ),
    .X(net352));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1032  (.A(\final_adder.$signal$1161 ),
    .B(\final_adder.g_new$1054 ),
    .X(net353));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1033  (.A(\final_adder.$signal$1162 ),
    .B(\final_adder.g_new$1019 ),
    .X(net354));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1034  (.A(\final_adder.$signal$1163 ),
    .B(\final_adder.g_new$1053 ),
    .X(net355));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1035  (.A(\final_adder.$signal$1164 ),
    .B(\final_adder.g_new$1017 ),
    .X(net356));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1036  (.A(\final_adder.$signal$1165 ),
    .B(\final_adder.g_new$1052 ),
    .X(net357));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1037  (.A(\final_adder.$signal$1166 ),
    .B(\final_adder.g_new$1015 ),
    .X(net358));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1038  (.A(\final_adder.$signal$1167 ),
    .B(\final_adder.g_new$1051 ),
    .X(net359));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1039  (.A(\final_adder.$signal$1168 ),
    .B(\final_adder.g_new$1013 ),
    .X(net360));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$104  (.A(\c$4358 ),
    .B(\s$4361 ),
    .COUT(\final_adder.$signal$210 ),
    .SUM(\final_adder.$signal$1194 ));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1040  (.A(\final_adder.$signal$1169 ),
    .B(\final_adder.g_new$1050 ),
    .X(net361));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1041  (.A(\final_adder.$signal$1170 ),
    .B(\final_adder.g_new$1011 ),
    .X(net363));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1042  (.A(\final_adder.$signal$1171 ),
    .B(\final_adder.g_new$1049 ),
    .X(net364));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1043  (.A(\final_adder.$signal$1172 ),
    .B(\final_adder.g_new$1009 ),
    .X(net365));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1044  (.A(\final_adder.$signal$1173 ),
    .B(\final_adder.g_new$1048 ),
    .X(net366));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1045  (.A(\final_adder.$signal$1174 ),
    .B(\final_adder.g_new$1007 ),
    .X(net367));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1046  (.A(\final_adder.$signal$1175 ),
    .B(\final_adder.g_new$1047 ),
    .X(net368));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1047  (.A(\final_adder.$signal$1176 ),
    .B(\final_adder.g_new$1005 ),
    .X(net369));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1048  (.A(\final_adder.$signal$1177 ),
    .B(\final_adder.g_new$1046 ),
    .X(net370));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1049  (.A(\final_adder.$signal$1178 ),
    .B(\final_adder.g_new$1003 ),
    .X(net371));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$105  (.A(\c$4360 ),
    .B(\s$4363 ),
    .COUT(\final_adder.$signal$212 ),
    .SUM(\final_adder.$signal$1195 ));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1050  (.A(\final_adder.$signal$1179 ),
    .B(\final_adder.g_new$1045 ),
    .X(net372));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1051  (.A(\final_adder.$signal$1180 ),
    .B(\final_adder.g_new$1001 ),
    .X(net374));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1052  (.A(\final_adder.$signal$1181 ),
    .B(\final_adder.g_new$1044 ),
    .X(net375));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1053  (.A(\final_adder.$signal$1182 ),
    .B(\final_adder.g_new$999 ),
    .X(net376));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1054  (.A(\final_adder.$signal$1183 ),
    .B(\final_adder.g_new$1043 ),
    .X(net377));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1055  (.A(\final_adder.$signal$1184 ),
    .B(\final_adder.g_new$997 ),
    .X(net378));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$1056  (.A(\final_adder.$signal$1185 ),
    .B(\final_adder.g_new$1042 ),
    .X(net379));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1057  (.A(\final_adder.$signal$1186 ),
    .B(\final_adder.g_new$995 ),
    .X(net380));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1058  (.A(\final_adder.$signal$1187 ),
    .B(\final_adder.g_new$1041 ),
    .X(net381));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$1059  (.A(\final_adder.$signal$1188 ),
    .B(\final_adder.g_new$993 ),
    .X(net382));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$106  (.A(\c$4362 ),
    .B(\s$4365 ),
    .COUT(\final_adder.$signal$214 ),
    .SUM(\final_adder.$signal$1196 ));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$1060  (.A(\final_adder.$signal$1189 ),
    .B(\final_adder.g_new$1040 ),
    .X(net383));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$1061  (.A(\final_adder.$signal$1190 ),
    .B(\final_adder.g_new$991 ),
    .X(net258));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$1062  (.A(\final_adder.$signal$1191 ),
    .B(\final_adder.g_new$1039 ),
    .X(net259));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$1063  (.A(\final_adder.$signal$1192 ),
    .B(\final_adder.g_new$989 ),
    .X(net260));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$1064  (.A(\final_adder.$signal$1193 ),
    .B(\final_adder.g_new$1038 ),
    .X(net261));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$1065  (.A(\final_adder.$signal$1194 ),
    .B(\final_adder.g_new$987 ),
    .X(net262));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$1066  (.A(\final_adder.$signal$1195 ),
    .B(\final_adder.g_new$1037 ),
    .X(net263));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1067  (.A(\final_adder.$signal$1196 ),
    .B(\final_adder.g_new$985 ),
    .X(net264));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1068  (.A(\final_adder.$signal$1197 ),
    .B(\final_adder.g_new$1036 ),
    .X(net265));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1069  (.A(\final_adder.$signal$1198 ),
    .B(\final_adder.g_new$983 ),
    .X(net266));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$107  (.A(\c$4364 ),
    .B(\s$4367 ),
    .COUT(\final_adder.$signal$216 ),
    .SUM(\final_adder.$signal$1197 ));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1070  (.A(\final_adder.$signal$1199 ),
    .B(\final_adder.g_new$1035 ),
    .X(net267));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1071  (.A(\final_adder.$signal$1200 ),
    .B(\final_adder.g_new$981 ),
    .X(net269));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1072  (.A(\final_adder.$signal$1201 ),
    .B(\final_adder.g_new$1034 ),
    .X(net270));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1073  (.A(\final_adder.$signal$1202 ),
    .B(\final_adder.g_new$979 ),
    .X(net271));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1074  (.A(\final_adder.$signal$1203 ),
    .B(\final_adder.g_new$1033 ),
    .X(net272));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1075  (.A(\final_adder.$signal$1204 ),
    .B(\final_adder.g_new$977 ),
    .X(net273));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1076  (.A(\final_adder.$signal$1205 ),
    .B(\final_adder.g_new$1032 ),
    .X(net274));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1077  (.A(\final_adder.$signal$1206 ),
    .B(\final_adder.g_new$975 ),
    .X(net275));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1078  (.A(\final_adder.$signal$1207 ),
    .B(\final_adder.g_new$1031 ),
    .X(net276));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1079  (.A(\final_adder.$signal$1208 ),
    .B(\final_adder.g_new$973 ),
    .X(net277));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$108  (.A(\c$4366 ),
    .B(\s$4369 ),
    .COUT(\final_adder.$signal$218 ),
    .SUM(\final_adder.$signal$1198 ));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1080  (.A(\final_adder.$signal$1209 ),
    .B(\final_adder.g_new$1030 ),
    .X(net278));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1081  (.A(\final_adder.$signal$1210 ),
    .B(\final_adder.g_new$971 ),
    .X(net280));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1082  (.A(\final_adder.$signal$1211 ),
    .B(\final_adder.g_new$1029 ),
    .X(net281));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1083  (.A(\final_adder.$signal$1212 ),
    .B(\final_adder.g_new$969 ),
    .X(net282));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1084  (.A(\final_adder.$signal$1213 ),
    .B(\final_adder.g_new$1028 ),
    .X(net283));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1085  (.A(\final_adder.$signal$1214 ),
    .B(\final_adder.g_new$967 ),
    .X(net284));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1086  (.A(\final_adder.$signal$1215 ),
    .B(\final_adder.g_new$1027 ),
    .X(net285));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1087  (.A(\final_adder.$signal$1216 ),
    .B(\final_adder.g_new$965 ),
    .X(net286));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$1088  (.A(\final_adder.$signal$1217 ),
    .B(\final_adder.g_new$1026 ),
    .X(net287));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$109  (.A(\c$4368 ),
    .B(\s$4371 ),
    .COUT(\final_adder.$signal$220 ),
    .SUM(\final_adder.$signal$1199 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$11  (.A(\c$4172 ),
    .B(\s$4175 ),
    .COUT(\final_adder.$signal$24 ),
    .SUM(\final_adder.$signal$1101 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$110  (.A(\c$4370 ),
    .B(\s$4373 ),
    .COUT(\final_adder.$signal$222 ),
    .SUM(\final_adder.$signal$1200 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$111  (.A(\c$4372 ),
    .B(\s$4375 ),
    .COUT(\final_adder.$signal$224 ),
    .SUM(\final_adder.$signal$1201 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$112  (.A(\c$4374 ),
    .B(\s$4377 ),
    .COUT(\final_adder.$signal$226 ),
    .SUM(\final_adder.$signal$1202 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$113  (.A(\c$4376 ),
    .B(\s$4379 ),
    .COUT(\final_adder.$signal$228 ),
    .SUM(\final_adder.$signal$1203 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$114  (.A(\c$4378 ),
    .B(\s$4381 ),
    .COUT(\final_adder.$signal$230 ),
    .SUM(\final_adder.$signal$1204 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$115  (.A(\c$4380 ),
    .B(\s$4383 ),
    .COUT(\final_adder.$signal$232 ),
    .SUM(\final_adder.$signal$1205 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$116  (.A(\c$4382 ),
    .B(\s$4385 ),
    .COUT(\final_adder.$signal$234 ),
    .SUM(\final_adder.$signal$1206 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$117  (.A(\c$4384 ),
    .B(\s$4387 ),
    .COUT(\final_adder.$signal$236 ),
    .SUM(\final_adder.$signal$1207 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$118  (.A(\c$4386 ),
    .B(\s$4389 ),
    .COUT(\final_adder.$signal$238 ),
    .SUM(\final_adder.$signal$1208 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$119  (.A(\c$4388 ),
    .B(\s$4391 ),
    .COUT(\final_adder.$signal$240 ),
    .SUM(\final_adder.$signal$1209 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$12  (.A(\c$4174 ),
    .B(\s$4177 ),
    .COUT(\final_adder.$signal$26 ),
    .SUM(\final_adder.$signal$1102 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$120  (.A(\c$4390 ),
    .B(\s$4393 ),
    .COUT(\final_adder.$signal$242 ),
    .SUM(\final_adder.$signal$1210 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$121  (.A(\c$4392 ),
    .B(\s$4395 ),
    .COUT(\final_adder.$signal$244 ),
    .SUM(\final_adder.$signal$1211 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$122  (.A(\c$4394 ),
    .B(\s$4397 ),
    .COUT(\final_adder.$signal$246 ),
    .SUM(\final_adder.$signal$1212 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$123  (.A(\c$4396 ),
    .B(\s$4399 ),
    .COUT(\final_adder.$signal$248 ),
    .SUM(\final_adder.$signal$1213 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$124  (.A(\c$4398 ),
    .B(\s$4401 ),
    .COUT(\final_adder.$signal$250 ),
    .SUM(\final_adder.$signal$1214 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$125  (.A(\c$4400 ),
    .B(\s$4403 ),
    .COUT(\final_adder.$signal$252 ),
    .SUM(\final_adder.$signal$1215 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$126  (.A(\c$4402 ),
    .B(\s$4405 ),
    .COUT(\final_adder.$signal$254 ),
    .SUM(\final_adder.$signal$1216 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$127  (.A(\c$4404 ),
    .B(\s$4407 ),
    .COUT(\final_adder.$signal$256 ),
    .SUM(\final_adder.$signal$1217 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$13  (.A(\c$4176 ),
    .B(\s$4179 ),
    .COUT(\final_adder.$signal$28 ),
    .SUM(\final_adder.$signal$1103 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$130  (.A(\final_adder.$signal$1214 ),
    .B(\final_adder.$signal$1215 ),
    .X(\final_adder.p_new$258 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$131  (.A1(\final_adder.$signal$1215 ),
    .A2(\final_adder.$signal$250 ),
    .B1(\final_adder.$signal$252 ),
    .X(\final_adder.g_new$259 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$132  (.A(\final_adder.$signal$1212 ),
    .B(\final_adder.$signal$1213 ),
    .X(\final_adder.p_new$260 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$133  (.A1(\final_adder.$signal$1213 ),
    .A2(\final_adder.$signal$246 ),
    .B1(\final_adder.$signal$248 ),
    .X(\final_adder.g_new$261 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$134  (.A(\final_adder.$signal$1210 ),
    .B(\final_adder.$signal$1211 ),
    .X(\final_adder.p_new$262 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$135  (.A1(\final_adder.$signal$1211 ),
    .A2(\final_adder.$signal$242 ),
    .B1(\final_adder.$signal$244 ),
    .X(\final_adder.g_new$263 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$136  (.A(\final_adder.$signal$1208 ),
    .B(\final_adder.$signal$1209 ),
    .X(\final_adder.p_new$264 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$137  (.A1(\final_adder.$signal$1209 ),
    .A2(\final_adder.$signal$238 ),
    .B1(\final_adder.$signal$240 ),
    .X(\final_adder.g_new$265 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$138  (.A(\final_adder.$signal$1206 ),
    .B(\final_adder.$signal$1207 ),
    .X(\final_adder.p_new$266 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$139  (.A1(\final_adder.$signal$1207 ),
    .A2(\final_adder.$signal$234 ),
    .B1(\final_adder.$signal$236 ),
    .X(\final_adder.g_new$267 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$14  (.A(\c$4178 ),
    .B(\s$4181 ),
    .COUT(\final_adder.$signal$30 ),
    .SUM(\final_adder.$signal$1104 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$140  (.A(\final_adder.$signal$1204 ),
    .B(\final_adder.$signal$1205 ),
    .X(\final_adder.p_new$268 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$141  (.A1(\final_adder.$signal$1205 ),
    .A2(\final_adder.$signal$230 ),
    .B1(\final_adder.$signal$232 ),
    .X(\final_adder.g_new$269 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$142  (.A(\final_adder.$signal$1202 ),
    .B(\final_adder.$signal$1203 ),
    .X(\final_adder.p_new$270 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$143  (.A1(\final_adder.$signal$1203 ),
    .A2(\final_adder.$signal$226 ),
    .B1(\final_adder.$signal$228 ),
    .X(\final_adder.g_new$271 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$144  (.A(\final_adder.$signal$1200 ),
    .B(\final_adder.$signal$1201 ),
    .X(\final_adder.p_new$272 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$145  (.A1(\final_adder.$signal$1201 ),
    .A2(\final_adder.$signal$222 ),
    .B1(\final_adder.$signal$224 ),
    .X(\final_adder.g_new$273 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$146  (.A(\final_adder.$signal$1198 ),
    .B(\final_adder.$signal$1199 ),
    .X(\final_adder.p_new$274 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$147  (.A1(\final_adder.$signal$1199 ),
    .A2(\final_adder.$signal$218 ),
    .B1(\final_adder.$signal$220 ),
    .X(\final_adder.g_new$275 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$148  (.A(\final_adder.$signal$1196 ),
    .B(\final_adder.$signal$1197 ),
    .X(\final_adder.p_new$276 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$149  (.A1(\final_adder.$signal$1197 ),
    .A2(\final_adder.$signal$214 ),
    .B1(\final_adder.$signal$216 ),
    .X(\final_adder.g_new$277 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$15  (.A(\c$4180 ),
    .B(\s$4183 ),
    .COUT(\final_adder.$signal$32 ),
    .SUM(\final_adder.$signal$1105 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$150  (.A(\final_adder.$signal$1194 ),
    .B(\final_adder.$signal$1195 ),
    .X(\final_adder.p_new$278 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$151  (.A1(\final_adder.$signal$1195 ),
    .A2(\final_adder.$signal$210 ),
    .B1(\final_adder.$signal$212 ),
    .X(\final_adder.g_new$279 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$152  (.A(\final_adder.$signal$1192 ),
    .B(\final_adder.$signal$1193 ),
    .X(\final_adder.p_new$280 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$153  (.A1(\final_adder.$signal$1193 ),
    .A2(\final_adder.$signal$206 ),
    .B1(\final_adder.$signal$208 ),
    .X(\final_adder.g_new$281 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$154  (.A(\final_adder.$signal$1190 ),
    .B(\final_adder.$signal$1191 ),
    .X(\final_adder.p_new$282 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$155  (.A1(\final_adder.$signal$1191 ),
    .A2(\final_adder.$signal$202 ),
    .B1(\final_adder.$signal$204 ),
    .X(\final_adder.g_new$283 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$156  (.A(\final_adder.$signal$1188 ),
    .B(\final_adder.$signal$1189 ),
    .X(\final_adder.p_new$284 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$157  (.A1(\final_adder.$signal$1189 ),
    .A2(\final_adder.$signal$198 ),
    .B1(\final_adder.$signal$200 ),
    .X(\final_adder.g_new$285 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$158  (.A(\final_adder.$signal$1186 ),
    .B(\final_adder.$signal$1187 ),
    .X(\final_adder.p_new$286 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$159  (.A1(\final_adder.$signal$1187 ),
    .A2(\final_adder.$signal$194 ),
    .B1(\final_adder.$signal$196 ),
    .X(\final_adder.g_new$287 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$16  (.A(\c$4182 ),
    .B(\s$4185 ),
    .COUT(\final_adder.$signal$34 ),
    .SUM(\final_adder.$signal$1106 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$160  (.A(\final_adder.$signal$1184 ),
    .B(\final_adder.$signal$1185 ),
    .X(\final_adder.p_new$288 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$161  (.A1(\final_adder.$signal$1185 ),
    .A2(\final_adder.$signal$190 ),
    .B1(\final_adder.$signal$192 ),
    .X(\final_adder.g_new$289 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$162  (.A(\final_adder.$signal$1182 ),
    .B(\final_adder.$signal$1183 ),
    .X(\final_adder.p_new$290 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$163  (.A1(\final_adder.$signal$1183 ),
    .A2(\final_adder.$signal$186 ),
    .B1(\final_adder.$signal$188 ),
    .X(\final_adder.g_new$291 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$164  (.A(\final_adder.$signal$1180 ),
    .B(\final_adder.$signal$1181 ),
    .X(\final_adder.p_new$292 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$165  (.A1(\final_adder.$signal$1181 ),
    .A2(\final_adder.$signal$182 ),
    .B1(\final_adder.$signal$184 ),
    .X(\final_adder.g_new$293 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$166  (.A(\final_adder.$signal$1178 ),
    .B(\final_adder.$signal$1179 ),
    .X(\final_adder.p_new$294 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$167  (.A1(\final_adder.$signal$1179 ),
    .A2(\final_adder.$signal$178 ),
    .B1(\final_adder.$signal$180 ),
    .X(\final_adder.g_new$295 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$168  (.A(\final_adder.$signal$1176 ),
    .B(\final_adder.$signal$1177 ),
    .X(\final_adder.p_new$296 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$169  (.A1(\final_adder.$signal$1177 ),
    .A2(\final_adder.$signal$174 ),
    .B1(\final_adder.$signal$176 ),
    .X(\final_adder.g_new$297 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$17  (.A(\c$4184 ),
    .B(\s$4187 ),
    .COUT(\final_adder.$signal$36 ),
    .SUM(\final_adder.$signal$1107 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$170  (.A(\final_adder.$signal$1174 ),
    .B(\final_adder.$signal$1175 ),
    .X(\final_adder.p_new$298 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$171  (.A1(\final_adder.$signal$1175 ),
    .A2(\final_adder.$signal$170 ),
    .B1(\final_adder.$signal$172 ),
    .X(\final_adder.g_new$299 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$172  (.A(\final_adder.$signal$1172 ),
    .B(\final_adder.$signal$1173 ),
    .X(\final_adder.p_new$300 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$173  (.A1(\final_adder.$signal$1173 ),
    .A2(\final_adder.$signal$166 ),
    .B1(\final_adder.$signal$168 ),
    .X(\final_adder.g_new$301 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$174  (.A(\final_adder.$signal$1170 ),
    .B(\final_adder.$signal$1171 ),
    .X(\final_adder.p_new$302 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$175  (.A1(\final_adder.$signal$1171 ),
    .A2(\final_adder.$signal$162 ),
    .B1(\final_adder.$signal$164 ),
    .X(\final_adder.g_new$303 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$176  (.A(\final_adder.$signal$1168 ),
    .B(\final_adder.$signal$1169 ),
    .X(\final_adder.p_new$304 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$177  (.A1(\final_adder.$signal$1169 ),
    .A2(\final_adder.$signal$158 ),
    .B1(\final_adder.$signal$160 ),
    .X(\final_adder.g_new$305 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$178  (.A(\final_adder.$signal$1166 ),
    .B(\final_adder.$signal$1167 ),
    .X(\final_adder.p_new$306 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$179  (.A1(\final_adder.$signal$1167 ),
    .A2(\final_adder.$signal$154 ),
    .B1(\final_adder.$signal$156 ),
    .X(\final_adder.g_new$307 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$18  (.A(\c$4186 ),
    .B(\s$4189 ),
    .COUT(\final_adder.$signal$38 ),
    .SUM(\final_adder.$signal$1108 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$180  (.A(\final_adder.$signal$1164 ),
    .B(\final_adder.$signal$1165 ),
    .X(\final_adder.p_new$308 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$181  (.A1(\final_adder.$signal$1165 ),
    .A2(\final_adder.$signal$150 ),
    .B1(\final_adder.$signal$152 ),
    .X(\final_adder.g_new$309 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$182  (.A(\final_adder.$signal$1162 ),
    .B(\final_adder.$signal$1163 ),
    .X(\final_adder.p_new$310 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$183  (.A1(\final_adder.$signal$1163 ),
    .A2(\final_adder.$signal$146 ),
    .B1(\final_adder.$signal$148 ),
    .X(\final_adder.g_new$311 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$184  (.A(\final_adder.$signal$1160 ),
    .B(\final_adder.$signal$1161 ),
    .X(\final_adder.p_new$312 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$185  (.A1(\final_adder.$signal$1161 ),
    .A2(\final_adder.$signal$142 ),
    .B1(\final_adder.$signal$144 ),
    .X(\final_adder.g_new$313 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$186  (.A(\final_adder.$signal$1158 ),
    .B(\final_adder.$signal$1159 ),
    .X(\final_adder.p_new$314 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$187  (.A1(\final_adder.$signal$1159 ),
    .A2(\final_adder.$signal$138 ),
    .B1(\final_adder.$signal$140 ),
    .X(\final_adder.g_new$315 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$188  (.A(\final_adder.$signal$1156 ),
    .B(\final_adder.$signal$1157 ),
    .X(\final_adder.p_new$316 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$189  (.A1(\final_adder.$signal$1157 ),
    .A2(\final_adder.$signal$134 ),
    .B1(\final_adder.$signal$136 ),
    .X(\final_adder.g_new$317 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$19  (.A(\c$4188 ),
    .B(\s$4191 ),
    .COUT(\final_adder.$signal$40 ),
    .SUM(\final_adder.$signal$1109 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$190  (.A(\final_adder.$signal$1154 ),
    .B(\final_adder.$signal$1155 ),
    .X(\final_adder.p_new$318 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$191  (.A1(\final_adder.$signal$1155 ),
    .A2(\final_adder.$signal$130 ),
    .B1(\final_adder.$signal$132 ),
    .X(\final_adder.g_new$319 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$192  (.A(\final_adder.$signal$1152 ),
    .B(\final_adder.$signal$1153 ),
    .X(\final_adder.p_new$320 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$193  (.A1(\final_adder.$signal$1153 ),
    .A2(\final_adder.$signal$126 ),
    .B1(\final_adder.$signal$128 ),
    .X(\final_adder.g_new$321 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$194  (.A(\final_adder.$signal$1150 ),
    .B(\final_adder.$signal$1151 ),
    .X(\final_adder.p_new$322 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$195  (.A1(\final_adder.$signal$1151 ),
    .A2(\final_adder.$signal$122 ),
    .B1(\final_adder.$signal$124 ),
    .X(\final_adder.g_new$323 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$196  (.A(\final_adder.$signal$1148 ),
    .B(\final_adder.$signal$1149 ),
    .X(\final_adder.p_new$324 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$197  (.A1(\final_adder.$signal$1149 ),
    .A2(\final_adder.$signal$118 ),
    .B1(\final_adder.$signal$120 ),
    .X(\final_adder.g_new$325 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$198  (.A(\final_adder.$signal$1146 ),
    .B(\final_adder.$signal$1147 ),
    .X(\final_adder.p_new$326 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$199  (.A1(\final_adder.$signal$1147 ),
    .A2(\final_adder.$signal$114 ),
    .B1(\final_adder.$signal$116 ),
    .X(\final_adder.g_new$327 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$2  (.A(\c$4154 ),
    .B(\s$4157 ),
    .COUT(\final_adder.$signal$6 ),
    .SUM(\final_adder.$signal$1092 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$20  (.A(\c$4190 ),
    .B(\s$4193 ),
    .COUT(\final_adder.$signal$42 ),
    .SUM(\final_adder.$signal$1110 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$200  (.A(\final_adder.$signal$111 ),
    .B(\final_adder.$signal$113 ),
    .X(\final_adder.p_new$328 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$201  (.A1(\final_adder.$signal$113 ),
    .A2(\final_adder.$signal$110 ),
    .B1(\final_adder.$signal$112 ),
    .X(\final_adder.g_new$329 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$202  (.A(\final_adder.$signal$107 ),
    .B(\final_adder.$signal$109 ),
    .X(\final_adder.p_new$330 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$203  (.A1(\final_adder.$signal$109 ),
    .A2(\final_adder.$signal$106 ),
    .B1(\final_adder.$signal$108 ),
    .X(\final_adder.g_new$331 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$204  (.A(\final_adder.$signal$103 ),
    .B(\final_adder.$signal$105 ),
    .X(\final_adder.p_new$332 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$205  (.A1(\final_adder.$signal$105 ),
    .A2(\final_adder.$signal$102 ),
    .B1(\final_adder.$signal$104 ),
    .X(\final_adder.g_new$333 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$206  (.A(\final_adder.$signal$1138 ),
    .B(\final_adder.$signal$101 ),
    .X(\final_adder.p_new$334 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$207  (.A1(\final_adder.$signal$101 ),
    .A2(\final_adder.$signal$98 ),
    .B1(\final_adder.$signal$100 ),
    .X(\final_adder.g_new$335 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$208  (.A(\final_adder.$signal$1136 ),
    .B(\final_adder.$signal$1137 ),
    .X(\final_adder.p_new$336 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$209  (.A1(\final_adder.$signal$1137 ),
    .A2(\final_adder.$signal$94 ),
    .B1(\final_adder.$signal$96 ),
    .X(\final_adder.g_new$337 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$21  (.A(\c$4192 ),
    .B(\s$4195 ),
    .COUT(\final_adder.$signal$44 ),
    .SUM(\final_adder.$signal$1111 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$210  (.A(\final_adder.$signal$1134 ),
    .B(\final_adder.$signal$1135 ),
    .X(\final_adder.p_new$338 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$211  (.A1(\final_adder.$signal$1135 ),
    .A2(\final_adder.$signal$90 ),
    .B1(\final_adder.$signal$92 ),
    .X(\final_adder.g_new$339 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$212  (.A(\final_adder.$signal$1132 ),
    .B(\final_adder.$signal$1133 ),
    .X(\final_adder.p_new$340 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$213  (.A1(\final_adder.$signal$1133 ),
    .A2(\final_adder.$signal$86 ),
    .B1(\final_adder.$signal$88 ),
    .X(\final_adder.g_new$341 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$214  (.A(\final_adder.$signal$1130 ),
    .B(\final_adder.$signal$1131 ),
    .X(\final_adder.p_new$342 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$215  (.A1(\final_adder.$signal$1131 ),
    .A2(\final_adder.$signal$82 ),
    .B1(\final_adder.$signal$84 ),
    .X(\final_adder.g_new$343 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$216  (.A(\final_adder.$signal$1128 ),
    .B(\final_adder.$signal$1129 ),
    .X(\final_adder.p_new$344 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$217  (.A1(\final_adder.$signal$1129 ),
    .A2(\final_adder.$signal$78 ),
    .B1(\final_adder.$signal$80 ),
    .X(\final_adder.g_new$345 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$218  (.A(\final_adder.$signal$1126 ),
    .B(\final_adder.$signal$1127 ),
    .X(\final_adder.p_new$346 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$219  (.A1(\final_adder.$signal$1127 ),
    .A2(\final_adder.$signal$74 ),
    .B1(\final_adder.$signal$76 ),
    .X(\final_adder.g_new$347 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$22  (.A(\c$4194 ),
    .B(\s$4197 ),
    .COUT(\final_adder.$signal$46 ),
    .SUM(\final_adder.$signal$1112 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$220  (.A(\final_adder.$signal$1124 ),
    .B(\final_adder.$signal$1125 ),
    .X(\final_adder.p_new$348 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$221  (.A1(\final_adder.$signal$1125 ),
    .A2(\final_adder.$signal$70 ),
    .B1(\final_adder.$signal$72 ),
    .X(\final_adder.g_new$349 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$222  (.A(\final_adder.$signal$1122 ),
    .B(\final_adder.$signal$1123 ),
    .X(\final_adder.p_new$350 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$223  (.A1(\final_adder.$signal$1123 ),
    .A2(\final_adder.$signal$66 ),
    .B1(\final_adder.$signal$68 ),
    .X(\final_adder.g_new$351 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$224  (.A(\final_adder.$signal$1120 ),
    .B(\final_adder.$signal$1121 ),
    .X(\final_adder.p_new$352 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$225  (.A1(\final_adder.$signal$1121 ),
    .A2(\final_adder.$signal$62 ),
    .B1(\final_adder.$signal$64 ),
    .X(\final_adder.g_new$353 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$226  (.A(\final_adder.$signal$1118 ),
    .B(\final_adder.$signal$1119 ),
    .X(\final_adder.p_new$354 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$227  (.A1(\final_adder.$signal$1119 ),
    .A2(\final_adder.$signal$58 ),
    .B1(\final_adder.$signal$60 ),
    .X(\final_adder.g_new$355 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$228  (.A(\final_adder.$signal$1116 ),
    .B(\final_adder.$signal$1117 ),
    .X(\final_adder.p_new$356 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$229  (.A1(\final_adder.$signal$1117 ),
    .A2(\final_adder.$signal$54 ),
    .B1(\final_adder.$signal$56 ),
    .X(\final_adder.g_new$357 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$23  (.A(\c$4196 ),
    .B(\s$4199 ),
    .COUT(\final_adder.$signal$48 ),
    .SUM(\final_adder.$signal$1113 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$230  (.A(\final_adder.$signal$1114 ),
    .B(\final_adder.$signal$1115 ),
    .X(\final_adder.p_new$358 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$231  (.A1(\final_adder.$signal$1115 ),
    .A2(\final_adder.$signal$50 ),
    .B1(\final_adder.$signal$52 ),
    .X(\final_adder.g_new$359 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$232  (.A(\final_adder.$signal$1112 ),
    .B(\final_adder.$signal$1113 ),
    .X(\final_adder.p_new$360 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$233  (.A1(\final_adder.$signal$1113 ),
    .A2(\final_adder.$signal$46 ),
    .B1(\final_adder.$signal$48 ),
    .X(\final_adder.g_new$361 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$234  (.A(\final_adder.$signal$1110 ),
    .B(\final_adder.$signal$1111 ),
    .X(\final_adder.p_new$362 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$235  (.A1(\final_adder.$signal$1111 ),
    .A2(\final_adder.$signal$42 ),
    .B1(\final_adder.$signal$44 ),
    .X(\final_adder.g_new$363 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$236  (.A(\final_adder.$signal$1108 ),
    .B(\final_adder.$signal$1109 ),
    .X(\final_adder.p_new$364 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$237  (.A1(\final_adder.$signal$1109 ),
    .A2(\final_adder.$signal$38 ),
    .B1(\final_adder.$signal$40 ),
    .X(\final_adder.g_new$365 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$238  (.A(\final_adder.$signal$1106 ),
    .B(\final_adder.$signal$1107 ),
    .X(\final_adder.p_new$366 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$239  (.A1(\final_adder.$signal$1107 ),
    .A2(\final_adder.$signal$34 ),
    .B1(\final_adder.$signal$36 ),
    .X(\final_adder.g_new$367 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$24  (.A(\c$4198 ),
    .B(\s$4201 ),
    .COUT(\final_adder.$signal$50 ),
    .SUM(\final_adder.$signal$1114 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$240  (.A(\final_adder.$signal$1104 ),
    .B(\final_adder.$signal$1105 ),
    .X(\final_adder.p_new$368 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$241  (.A1(\final_adder.$signal$1105 ),
    .A2(\final_adder.$signal$30 ),
    .B1(\final_adder.$signal$32 ),
    .X(\final_adder.g_new$369 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$242  (.A(\final_adder.$signal$1102 ),
    .B(\final_adder.$signal$1103 ),
    .X(\final_adder.p_new$370 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$243  (.A1(\final_adder.$signal$1103 ),
    .A2(\final_adder.$signal$26 ),
    .B1(\final_adder.$signal$28 ),
    .X(\final_adder.g_new$371 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$244  (.A(\final_adder.$signal$1100 ),
    .B(\final_adder.$signal$1101 ),
    .X(\final_adder.p_new$372 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$245  (.A1(\final_adder.$signal$1101 ),
    .A2(\final_adder.$signal$22 ),
    .B1(\final_adder.$signal$24 ),
    .X(\final_adder.g_new$373 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$246  (.A(\final_adder.$signal$1098 ),
    .B(\final_adder.$signal$1099 ),
    .X(\final_adder.p_new$374 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$247  (.A1(\final_adder.$signal$1099 ),
    .A2(\final_adder.$signal$18 ),
    .B1(\final_adder.$signal$20 ),
    .X(\final_adder.g_new$375 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$248  (.A(\final_adder.$signal$1096 ),
    .B(\final_adder.$signal$1097 ),
    .X(\final_adder.p_new$376 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$249  (.A1(\final_adder.$signal$1097 ),
    .A2(\final_adder.$signal$14 ),
    .B1(\final_adder.$signal$16 ),
    .X(\final_adder.g_new$377 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$25  (.A(\c$4200 ),
    .B(\s$4203 ),
    .COUT(\final_adder.$signal$52 ),
    .SUM(\final_adder.$signal$1115 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$250  (.A(\final_adder.$signal$1094 ),
    .B(\final_adder.$signal$1095 ),
    .X(\final_adder.p_new$378 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$251  (.A1(\final_adder.$signal$1095 ),
    .A2(\final_adder.$signal$10 ),
    .B1(\final_adder.$signal$12 ),
    .X(\final_adder.g_new$379 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$252  (.A(\final_adder.$signal$1092 ),
    .B(\final_adder.$signal$1093 ),
    .X(\final_adder.p_new$380 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$253  (.A1(\final_adder.$signal$1093 ),
    .A2(\final_adder.$signal$6 ),
    .B1(\final_adder.$signal$8 ),
    .X(\final_adder.g_new$381 ));
 sky130_fd_sc_hd__a21o_4 \final_adder.U$$255  (.A1(\final_adder.$signal$1091 ),
    .A2(\final_adder.$signal ),
    .B1(\final_adder.$signal$4 ),
    .X(\final_adder.g_new$383 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$258  (.A(\final_adder.p_new$260 ),
    .B(\final_adder.p_new$258 ),
    .X(\final_adder.p_new$386 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$259  (.A1(\final_adder.p_new$258 ),
    .A2(\final_adder.g_new$261 ),
    .B1(\final_adder.g_new$259 ),
    .X(\final_adder.g_new$387 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$26  (.A(\c$4202 ),
    .B(\s$4205 ),
    .COUT(\final_adder.$signal$54 ),
    .SUM(\final_adder.$signal$1116 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$260  (.A(\final_adder.p_new$262 ),
    .B(\final_adder.p_new$260 ),
    .X(\final_adder.p_new$388 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$261  (.A1(\final_adder.p_new$260 ),
    .A2(\final_adder.g_new$263 ),
    .B1(\final_adder.g_new$261 ),
    .X(\final_adder.g_new$389 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$262  (.A(\final_adder.p_new$264 ),
    .B(\final_adder.p_new$262 ),
    .X(\final_adder.p_new$390 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$263  (.A1(\final_adder.p_new$262 ),
    .A2(\final_adder.g_new$265 ),
    .B1(\final_adder.g_new$263 ),
    .X(\final_adder.g_new$391 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$264  (.A(\final_adder.p_new$266 ),
    .B(\final_adder.p_new$264 ),
    .X(\final_adder.p_new$392 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$265  (.A1(\final_adder.p_new$264 ),
    .A2(\final_adder.g_new$267 ),
    .B1(\final_adder.g_new$265 ),
    .X(\final_adder.g_new$393 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$266  (.A(\final_adder.p_new$268 ),
    .B(\final_adder.p_new$266 ),
    .X(\final_adder.p_new$394 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$267  (.A1(\final_adder.p_new$266 ),
    .A2(\final_adder.g_new$269 ),
    .B1(\final_adder.g_new$267 ),
    .X(\final_adder.g_new$395 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$268  (.A(\final_adder.p_new$270 ),
    .B(\final_adder.p_new$268 ),
    .X(\final_adder.p_new$396 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$269  (.A1(\final_adder.p_new$268 ),
    .A2(\final_adder.g_new$271 ),
    .B1(\final_adder.g_new$269 ),
    .X(\final_adder.g_new$397 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$27  (.A(\c$4204 ),
    .B(\s$4207 ),
    .COUT(\final_adder.$signal$56 ),
    .SUM(\final_adder.$signal$1117 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$270  (.A(\final_adder.p_new$272 ),
    .B(\final_adder.p_new$270 ),
    .X(\final_adder.p_new$398 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$271  (.A1(\final_adder.p_new$270 ),
    .A2(\final_adder.g_new$273 ),
    .B1(\final_adder.g_new$271 ),
    .X(\final_adder.g_new$399 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$272  (.A(\final_adder.p_new$274 ),
    .B(\final_adder.p_new$272 ),
    .X(\final_adder.p_new$400 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$273  (.A1(\final_adder.p_new$272 ),
    .A2(\final_adder.g_new$275 ),
    .B1(\final_adder.g_new$273 ),
    .X(\final_adder.g_new$401 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$274  (.A(\final_adder.p_new$276 ),
    .B(\final_adder.p_new$274 ),
    .X(\final_adder.p_new$402 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$275  (.A1(\final_adder.p_new$274 ),
    .A2(\final_adder.g_new$277 ),
    .B1(\final_adder.g_new$275 ),
    .X(\final_adder.g_new$403 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$276  (.A(\final_adder.p_new$278 ),
    .B(\final_adder.p_new$276 ),
    .X(\final_adder.p_new$404 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$277  (.A1(\final_adder.p_new$276 ),
    .A2(\final_adder.g_new$279 ),
    .B1(\final_adder.g_new$277 ),
    .X(\final_adder.g_new$405 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$278  (.A(\final_adder.p_new$280 ),
    .B(\final_adder.p_new$278 ),
    .X(\final_adder.p_new$406 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$279  (.A1(\final_adder.p_new$278 ),
    .A2(\final_adder.g_new$281 ),
    .B1(\final_adder.g_new$279 ),
    .X(\final_adder.g_new$407 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$28  (.A(\c$4206 ),
    .B(\s$4209 ),
    .COUT(\final_adder.$signal$58 ),
    .SUM(\final_adder.$signal$1118 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$280  (.A(\final_adder.p_new$282 ),
    .B(\final_adder.p_new$280 ),
    .X(\final_adder.p_new$408 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$281  (.A1(\final_adder.p_new$280 ),
    .A2(\final_adder.g_new$283 ),
    .B1(\final_adder.g_new$281 ),
    .X(\final_adder.g_new$409 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$282  (.A(\final_adder.p_new$284 ),
    .B(\final_adder.p_new$282 ),
    .X(\final_adder.p_new$410 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$283  (.A1(\final_adder.p_new$282 ),
    .A2(\final_adder.g_new$285 ),
    .B1(\final_adder.g_new$283 ),
    .X(\final_adder.g_new$411 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$284  (.A(\final_adder.p_new$286 ),
    .B(\final_adder.p_new$284 ),
    .X(\final_adder.p_new$412 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$285  (.A1(\final_adder.p_new$284 ),
    .A2(\final_adder.g_new$287 ),
    .B1(\final_adder.g_new$285 ),
    .X(\final_adder.g_new$413 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$286  (.A(\final_adder.p_new$288 ),
    .B(\final_adder.p_new$286 ),
    .X(\final_adder.p_new$414 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$287  (.A1(\final_adder.p_new$286 ),
    .A2(\final_adder.g_new$289 ),
    .B1(\final_adder.g_new$287 ),
    .X(\final_adder.g_new$415 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$288  (.A(\final_adder.p_new$290 ),
    .B(\final_adder.p_new$288 ),
    .X(\final_adder.p_new$416 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$289  (.A1(\final_adder.p_new$288 ),
    .A2(\final_adder.g_new$291 ),
    .B1(\final_adder.g_new$289 ),
    .X(\final_adder.g_new$417 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$29  (.A(\c$4208 ),
    .B(\s$4211 ),
    .COUT(\final_adder.$signal$60 ),
    .SUM(\final_adder.$signal$1119 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$290  (.A(\final_adder.p_new$292 ),
    .B(\final_adder.p_new$290 ),
    .X(\final_adder.p_new$418 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$291  (.A1(\final_adder.p_new$290 ),
    .A2(\final_adder.g_new$293 ),
    .B1(\final_adder.g_new$291 ),
    .X(\final_adder.g_new$419 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$292  (.A(\final_adder.p_new$294 ),
    .B(\final_adder.p_new$292 ),
    .X(\final_adder.p_new$420 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$293  (.A1(\final_adder.p_new$292 ),
    .A2(\final_adder.g_new$295 ),
    .B1(\final_adder.g_new$293 ),
    .X(\final_adder.g_new$421 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$294  (.A(\final_adder.p_new$296 ),
    .B(\final_adder.p_new$294 ),
    .X(\final_adder.p_new$422 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$295  (.A1(\final_adder.p_new$294 ),
    .A2(\final_adder.g_new$297 ),
    .B1(\final_adder.g_new$295 ),
    .X(\final_adder.g_new$423 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$296  (.A(\final_adder.p_new$298 ),
    .B(\final_adder.p_new$296 ),
    .X(\final_adder.p_new$424 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$297  (.A1(\final_adder.p_new$296 ),
    .A2(\final_adder.g_new$299 ),
    .B1(\final_adder.g_new$297 ),
    .X(\final_adder.g_new$425 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$298  (.A(\final_adder.p_new$300 ),
    .B(\final_adder.p_new$298 ),
    .X(\final_adder.p_new$426 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$299  (.A1(\final_adder.p_new$298 ),
    .A2(\final_adder.g_new$301 ),
    .B1(\final_adder.g_new$299 ),
    .X(\final_adder.g_new$427 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$3  (.A(\c$4156 ),
    .B(\s$4159 ),
    .COUT(\final_adder.$signal$8 ),
    .SUM(\final_adder.$signal$1093 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$30  (.A(\c$4210 ),
    .B(\s$4213 ),
    .COUT(\final_adder.$signal$62 ),
    .SUM(\final_adder.$signal$1120 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$300  (.A(\final_adder.p_new$302 ),
    .B(\final_adder.p_new$300 ),
    .X(\final_adder.p_new$428 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$301  (.A1(\final_adder.p_new$300 ),
    .A2(\final_adder.g_new$303 ),
    .B1(\final_adder.g_new$301 ),
    .X(\final_adder.g_new$429 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$302  (.A(\final_adder.p_new$304 ),
    .B(\final_adder.p_new$302 ),
    .X(\final_adder.p_new$430 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$303  (.A1(\final_adder.p_new$302 ),
    .A2(\final_adder.g_new$305 ),
    .B1(\final_adder.g_new$303 ),
    .X(\final_adder.g_new$431 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$304  (.A(\final_adder.p_new$306 ),
    .B(\final_adder.p_new$304 ),
    .X(\final_adder.p_new$432 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$305  (.A1(\final_adder.p_new$304 ),
    .A2(\final_adder.g_new$307 ),
    .B1(\final_adder.g_new$305 ),
    .X(\final_adder.g_new$433 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$306  (.A(\final_adder.p_new$308 ),
    .B(\final_adder.p_new$306 ),
    .X(\final_adder.p_new$434 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$307  (.A1(\final_adder.p_new$306 ),
    .A2(\final_adder.g_new$309 ),
    .B1(\final_adder.g_new$307 ),
    .X(\final_adder.g_new$435 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$308  (.A(\final_adder.p_new$310 ),
    .B(\final_adder.p_new$308 ),
    .X(\final_adder.p_new$436 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$309  (.A1(\final_adder.p_new$308 ),
    .A2(\final_adder.g_new$311 ),
    .B1(\final_adder.g_new$309 ),
    .X(\final_adder.g_new$437 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$31  (.A(\c$4212 ),
    .B(\s$4215 ),
    .COUT(\final_adder.$signal$64 ),
    .SUM(\final_adder.$signal$1121 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$310  (.A(\final_adder.p_new$312 ),
    .B(\final_adder.p_new$310 ),
    .X(\final_adder.p_new$438 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$311  (.A1(\final_adder.p_new$310 ),
    .A2(\final_adder.g_new$313 ),
    .B1(\final_adder.g_new$311 ),
    .X(\final_adder.g_new$439 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$312  (.A(\final_adder.p_new$314 ),
    .B(\final_adder.p_new$312 ),
    .X(\final_adder.p_new$440 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$313  (.A1(\final_adder.p_new$312 ),
    .A2(\final_adder.g_new$315 ),
    .B1(\final_adder.g_new$313 ),
    .X(\final_adder.g_new$441 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$314  (.A(\final_adder.p_new$316 ),
    .B(\final_adder.p_new$314 ),
    .X(\final_adder.p_new$442 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$315  (.A1(\final_adder.p_new$314 ),
    .A2(\final_adder.g_new$317 ),
    .B1(\final_adder.g_new$315 ),
    .X(\final_adder.g_new$443 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$316  (.A(\final_adder.p_new$318 ),
    .B(\final_adder.p_new$316 ),
    .X(\final_adder.p_new$444 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$317  (.A1(\final_adder.p_new$316 ),
    .A2(\final_adder.g_new$319 ),
    .B1(\final_adder.g_new$317 ),
    .X(\final_adder.g_new$445 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$318  (.A(\final_adder.p_new$320 ),
    .B(\final_adder.p_new$318 ),
    .X(\final_adder.p_new$446 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$319  (.A1(\final_adder.p_new$318 ),
    .A2(\final_adder.g_new$321 ),
    .B1(\final_adder.g_new$319 ),
    .X(\final_adder.g_new$447 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$32  (.A(\c$4214 ),
    .B(\s$4217 ),
    .COUT(\final_adder.$signal$66 ),
    .SUM(\final_adder.$signal$1122 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$320  (.A(\final_adder.p_new$322 ),
    .B(\final_adder.p_new$320 ),
    .X(\final_adder.p_new$448 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$321  (.A1(\final_adder.p_new$320 ),
    .A2(\final_adder.g_new$323 ),
    .B1(\final_adder.g_new$321 ),
    .X(\final_adder.g_new$449 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$322  (.A(\final_adder.p_new$324 ),
    .B(\final_adder.p_new$322 ),
    .X(\final_adder.p_new$450 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$323  (.A1(\final_adder.p_new$322 ),
    .A2(\final_adder.g_new$325 ),
    .B1(\final_adder.g_new$323 ),
    .X(\final_adder.g_new$451 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$324  (.A(\final_adder.p_new$326 ),
    .B(\final_adder.p_new$324 ),
    .X(\final_adder.p_new$452 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$325  (.A1(\final_adder.p_new$324 ),
    .A2(\final_adder.g_new$327 ),
    .B1(\final_adder.g_new$325 ),
    .X(\final_adder.g_new$453 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$326  (.A(\final_adder.p_new$328 ),
    .B(\final_adder.p_new$326 ),
    .X(\final_adder.p_new$454 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$327  (.A1(\final_adder.p_new$326 ),
    .A2(\final_adder.g_new$329 ),
    .B1(\final_adder.g_new$327 ),
    .X(\final_adder.g_new$455 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$328  (.A(\final_adder.p_new$330 ),
    .B(\final_adder.p_new$328 ),
    .X(\final_adder.p_new$456 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$329  (.A1(\final_adder.p_new$328 ),
    .A2(\final_adder.g_new$331 ),
    .B1(\final_adder.g_new$329 ),
    .X(\final_adder.g_new$457 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$33  (.A(\c$4216 ),
    .B(\s$4219 ),
    .COUT(\final_adder.$signal$68 ),
    .SUM(\final_adder.$signal$1123 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$330  (.A(\final_adder.p_new$332 ),
    .B(\final_adder.p_new$330 ),
    .X(\final_adder.p_new$458 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$331  (.A1(\final_adder.p_new$330 ),
    .A2(\final_adder.g_new$333 ),
    .B1(\final_adder.g_new$331 ),
    .X(\final_adder.g_new$459 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$332  (.A(\final_adder.p_new$334 ),
    .B(\final_adder.p_new$332 ),
    .X(\final_adder.p_new$460 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$333  (.A1(\final_adder.p_new$332 ),
    .A2(\final_adder.g_new$335 ),
    .B1(\final_adder.g_new$333 ),
    .X(\final_adder.g_new$461 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$334  (.A(\final_adder.p_new$336 ),
    .B(\final_adder.p_new$334 ),
    .X(\final_adder.p_new$462 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$335  (.A1(\final_adder.p_new$334 ),
    .A2(\final_adder.g_new$337 ),
    .B1(\final_adder.g_new$335 ),
    .X(\final_adder.g_new$463 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$336  (.A(\final_adder.p_new$338 ),
    .B(\final_adder.p_new$336 ),
    .X(\final_adder.p_new$464 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$337  (.A1(\final_adder.p_new$336 ),
    .A2(\final_adder.g_new$339 ),
    .B1(\final_adder.g_new$337 ),
    .X(\final_adder.g_new$465 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$338  (.A(\final_adder.p_new$340 ),
    .B(\final_adder.p_new$338 ),
    .X(\final_adder.p_new$466 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$339  (.A1(\final_adder.p_new$338 ),
    .A2(\final_adder.g_new$341 ),
    .B1(\final_adder.g_new$339 ),
    .X(\final_adder.g_new$467 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$34  (.A(\c$4218 ),
    .B(\s$4221 ),
    .COUT(\final_adder.$signal$70 ),
    .SUM(\final_adder.$signal$1124 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$340  (.A(\final_adder.p_new$342 ),
    .B(\final_adder.p_new$340 ),
    .X(\final_adder.p_new$468 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$341  (.A1(\final_adder.p_new$340 ),
    .A2(\final_adder.g_new$343 ),
    .B1(\final_adder.g_new$341 ),
    .X(\final_adder.g_new$469 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$342  (.A(\final_adder.p_new$344 ),
    .B(\final_adder.p_new$342 ),
    .X(\final_adder.p_new$470 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$343  (.A1(\final_adder.p_new$342 ),
    .A2(\final_adder.g_new$345 ),
    .B1(\final_adder.g_new$343 ),
    .X(\final_adder.g_new$471 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$344  (.A(\final_adder.p_new$346 ),
    .B(\final_adder.p_new$344 ),
    .X(\final_adder.p_new$472 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$345  (.A1(\final_adder.p_new$344 ),
    .A2(\final_adder.g_new$347 ),
    .B1(\final_adder.g_new$345 ),
    .X(\final_adder.g_new$473 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$346  (.A(\final_adder.p_new$348 ),
    .B(\final_adder.p_new$346 ),
    .X(\final_adder.p_new$474 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$347  (.A1(\final_adder.p_new$346 ),
    .A2(\final_adder.g_new$349 ),
    .B1(\final_adder.g_new$347 ),
    .X(\final_adder.g_new$475 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$348  (.A(\final_adder.p_new$350 ),
    .B(\final_adder.p_new$348 ),
    .X(\final_adder.p_new$476 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$349  (.A1(\final_adder.p_new$348 ),
    .A2(\final_adder.g_new$351 ),
    .B1(\final_adder.g_new$349 ),
    .X(\final_adder.g_new$477 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$35  (.A(\c$4220 ),
    .B(\s$4223 ),
    .COUT(\final_adder.$signal$72 ),
    .SUM(\final_adder.$signal$1125 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$350  (.A(\final_adder.p_new$352 ),
    .B(\final_adder.p_new$350 ),
    .X(\final_adder.p_new$478 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$351  (.A1(\final_adder.p_new$350 ),
    .A2(\final_adder.g_new$353 ),
    .B1(\final_adder.g_new$351 ),
    .X(\final_adder.g_new$479 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$352  (.A(\final_adder.p_new$354 ),
    .B(\final_adder.p_new$352 ),
    .X(\final_adder.p_new$480 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$353  (.A1(\final_adder.p_new$352 ),
    .A2(\final_adder.g_new$355 ),
    .B1(\final_adder.g_new$353 ),
    .X(\final_adder.g_new$481 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$354  (.A(\final_adder.p_new$356 ),
    .B(\final_adder.p_new$354 ),
    .X(\final_adder.p_new$482 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$355  (.A1(\final_adder.p_new$354 ),
    .A2(\final_adder.g_new$357 ),
    .B1(\final_adder.g_new$355 ),
    .X(\final_adder.g_new$483 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$356  (.A(\final_adder.p_new$358 ),
    .B(\final_adder.p_new$356 ),
    .X(\final_adder.p_new$484 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$357  (.A1(\final_adder.p_new$356 ),
    .A2(\final_adder.g_new$359 ),
    .B1(\final_adder.g_new$357 ),
    .X(\final_adder.g_new$485 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$358  (.A(\final_adder.p_new$360 ),
    .B(\final_adder.p_new$358 ),
    .X(\final_adder.p_new$486 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$359  (.A1(\final_adder.p_new$358 ),
    .A2(\final_adder.g_new$361 ),
    .B1(\final_adder.g_new$359 ),
    .X(\final_adder.g_new$487 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$36  (.A(\c$4222 ),
    .B(\s$4225 ),
    .COUT(\final_adder.$signal$74 ),
    .SUM(\final_adder.$signal$1126 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$360  (.A(\final_adder.p_new$362 ),
    .B(\final_adder.p_new$360 ),
    .X(\final_adder.p_new$488 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$361  (.A1(\final_adder.p_new$360 ),
    .A2(\final_adder.g_new$363 ),
    .B1(\final_adder.g_new$361 ),
    .X(\final_adder.g_new$489 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$362  (.A(\final_adder.p_new$364 ),
    .B(\final_adder.p_new$362 ),
    .X(\final_adder.p_new$490 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$363  (.A1(\final_adder.p_new$362 ),
    .A2(\final_adder.g_new$365 ),
    .B1(\final_adder.g_new$363 ),
    .X(\final_adder.g_new$491 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$364  (.A(\final_adder.p_new$366 ),
    .B(\final_adder.p_new$364 ),
    .X(\final_adder.p_new$492 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$365  (.A1(\final_adder.p_new$364 ),
    .A2(\final_adder.g_new$367 ),
    .B1(\final_adder.g_new$365 ),
    .X(\final_adder.g_new$493 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$366  (.A(\final_adder.p_new$368 ),
    .B(\final_adder.p_new$366 ),
    .X(\final_adder.p_new$494 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$367  (.A1(\final_adder.p_new$366 ),
    .A2(\final_adder.g_new$369 ),
    .B1(\final_adder.g_new$367 ),
    .X(\final_adder.g_new$495 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$368  (.A(\final_adder.p_new$370 ),
    .B(\final_adder.p_new$368 ),
    .X(\final_adder.p_new$496 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$369  (.A1(\final_adder.p_new$368 ),
    .A2(\final_adder.g_new$371 ),
    .B1(\final_adder.g_new$369 ),
    .X(\final_adder.g_new$497 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$37  (.A(\c$4224 ),
    .B(\s$4227 ),
    .COUT(\final_adder.$signal$76 ),
    .SUM(\final_adder.$signal$1127 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$370  (.A(\final_adder.p_new$372 ),
    .B(\final_adder.p_new$370 ),
    .X(\final_adder.p_new$498 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$371  (.A1(\final_adder.p_new$370 ),
    .A2(\final_adder.g_new$373 ),
    .B1(\final_adder.g_new$371 ),
    .X(\final_adder.g_new$499 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$372  (.A(\final_adder.p_new$374 ),
    .B(\final_adder.p_new$372 ),
    .X(\final_adder.p_new$500 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$373  (.A1(\final_adder.p_new$372 ),
    .A2(\final_adder.g_new$375 ),
    .B1(\final_adder.g_new$373 ),
    .X(\final_adder.g_new$501 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$374  (.A(\final_adder.p_new$376 ),
    .B(\final_adder.p_new$374 ),
    .X(\final_adder.p_new$502 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$375  (.A1(\final_adder.p_new$374 ),
    .A2(\final_adder.g_new$377 ),
    .B1(\final_adder.g_new$375 ),
    .X(\final_adder.g_new$503 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$376  (.A(\final_adder.p_new$378 ),
    .B(\final_adder.p_new$376 ),
    .X(\final_adder.p_new$504 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$377  (.A1(\final_adder.p_new$376 ),
    .A2(\final_adder.g_new$379 ),
    .B1(\final_adder.g_new$377 ),
    .X(\final_adder.g_new$505 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$378  (.A(\final_adder.p_new$380 ),
    .B(\final_adder.p_new$378 ),
    .X(\final_adder.p_new$506 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$379  (.A1(\final_adder.p_new$378 ),
    .A2(\final_adder.g_new$381 ),
    .B1(\final_adder.g_new$379 ),
    .X(\final_adder.g_new$507 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$38  (.A(\c$4226 ),
    .B(\s$4229 ),
    .COUT(\final_adder.$signal$78 ),
    .SUM(\final_adder.$signal$1128 ));
 sky130_fd_sc_hd__a21o_4 \final_adder.U$$381  (.A1(\final_adder.p_new$380 ),
    .A2(\final_adder.g_new$383 ),
    .B1(\final_adder.g_new$381 ),
    .X(\final_adder.g_new$509 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$384  (.A(\final_adder.p_new$390 ),
    .B(\final_adder.p_new$386 ),
    .X(\final_adder.p_new$512 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$385  (.A1(\final_adder.p_new$386 ),
    .A2(\final_adder.g_new$391 ),
    .B1(\final_adder.g_new$387 ),
    .X(\final_adder.g_new$513 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$386  (.A(\final_adder.p_new$392 ),
    .B(\final_adder.p_new$388 ),
    .X(\final_adder.p_new$514 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$387  (.A1(\final_adder.p_new$388 ),
    .A2(\final_adder.g_new$393 ),
    .B1(\final_adder.g_new$389 ),
    .X(\final_adder.g_new$515 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$388  (.A(\final_adder.p_new$394 ),
    .B(\final_adder.p_new$390 ),
    .X(\final_adder.p_new$516 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$389  (.A1(\final_adder.p_new$390 ),
    .A2(\final_adder.g_new$395 ),
    .B1(\final_adder.g_new$391 ),
    .X(\final_adder.g_new$517 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$39  (.A(\c$4228 ),
    .B(\s$4231 ),
    .COUT(\final_adder.$signal$80 ),
    .SUM(\final_adder.$signal$1129 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$390  (.A(\final_adder.p_new$396 ),
    .B(\final_adder.p_new$392 ),
    .X(\final_adder.p_new$518 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$391  (.A1(\final_adder.p_new$392 ),
    .A2(\final_adder.g_new$397 ),
    .B1(\final_adder.g_new$393 ),
    .X(\final_adder.g_new$519 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$392  (.A(\final_adder.p_new$398 ),
    .B(\final_adder.p_new$394 ),
    .X(\final_adder.p_new$520 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$393  (.A1(\final_adder.p_new$394 ),
    .A2(\final_adder.g_new$399 ),
    .B1(\final_adder.g_new$395 ),
    .X(\final_adder.g_new$521 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$394  (.A(\final_adder.p_new$400 ),
    .B(\final_adder.p_new$396 ),
    .X(\final_adder.p_new$522 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$395  (.A1(\final_adder.p_new$396 ),
    .A2(\final_adder.g_new$401 ),
    .B1(\final_adder.g_new$397 ),
    .X(\final_adder.g_new$523 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$396  (.A(\final_adder.p_new$402 ),
    .B(\final_adder.p_new$398 ),
    .X(\final_adder.p_new$524 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$397  (.A1(\final_adder.p_new$398 ),
    .A2(\final_adder.g_new$403 ),
    .B1(\final_adder.g_new$399 ),
    .X(\final_adder.g_new$525 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$398  (.A(\final_adder.p_new$404 ),
    .B(\final_adder.p_new$400 ),
    .X(\final_adder.p_new$526 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$399  (.A1(\final_adder.p_new$400 ),
    .A2(\final_adder.g_new$405 ),
    .B1(\final_adder.g_new$401 ),
    .X(\final_adder.g_new$527 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$4  (.A(\c$4158 ),
    .B(\s$4161 ),
    .COUT(\final_adder.$signal$10 ),
    .SUM(\final_adder.$signal$1094 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$40  (.A(\c$4230 ),
    .B(\s$4233 ),
    .COUT(\final_adder.$signal$82 ),
    .SUM(\final_adder.$signal$1130 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$400  (.A(\final_adder.p_new$406 ),
    .B(\final_adder.p_new$402 ),
    .X(\final_adder.p_new$528 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$401  (.A1(\final_adder.p_new$402 ),
    .A2(\final_adder.g_new$407 ),
    .B1(\final_adder.g_new$403 ),
    .X(\final_adder.g_new$529 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$402  (.A(\final_adder.p_new$408 ),
    .B(\final_adder.p_new$404 ),
    .X(\final_adder.p_new$530 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$403  (.A1(\final_adder.p_new$404 ),
    .A2(\final_adder.g_new$409 ),
    .B1(\final_adder.g_new$405 ),
    .X(\final_adder.g_new$531 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$404  (.A(\final_adder.p_new$410 ),
    .B(\final_adder.p_new$406 ),
    .X(\final_adder.p_new$532 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$405  (.A1(\final_adder.p_new$406 ),
    .A2(\final_adder.g_new$411 ),
    .B1(\final_adder.g_new$407 ),
    .X(\final_adder.g_new$533 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$406  (.A(\final_adder.p_new$412 ),
    .B(\final_adder.p_new$408 ),
    .X(\final_adder.p_new$534 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$407  (.A1(\final_adder.p_new$408 ),
    .A2(\final_adder.g_new$413 ),
    .B1(\final_adder.g_new$409 ),
    .X(\final_adder.g_new$535 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$408  (.A(\final_adder.p_new$414 ),
    .B(\final_adder.p_new$410 ),
    .X(\final_adder.p_new$536 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$409  (.A1(\final_adder.p_new$410 ),
    .A2(\final_adder.g_new$415 ),
    .B1(\final_adder.g_new$411 ),
    .X(\final_adder.g_new$537 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$41  (.A(\c$4232 ),
    .B(\s$4235 ),
    .COUT(\final_adder.$signal$84 ),
    .SUM(\final_adder.$signal$1131 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$410  (.A(\final_adder.p_new$416 ),
    .B(\final_adder.p_new$412 ),
    .X(\final_adder.p_new$538 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$411  (.A1(\final_adder.p_new$412 ),
    .A2(\final_adder.g_new$417 ),
    .B1(\final_adder.g_new$413 ),
    .X(\final_adder.g_new$539 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$412  (.A(\final_adder.p_new$418 ),
    .B(\final_adder.p_new$414 ),
    .X(\final_adder.p_new$540 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$413  (.A1(\final_adder.p_new$414 ),
    .A2(\final_adder.g_new$419 ),
    .B1(\final_adder.g_new$415 ),
    .X(\final_adder.g_new$541 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$414  (.A(\final_adder.p_new$420 ),
    .B(\final_adder.p_new$416 ),
    .X(\final_adder.p_new$542 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$415  (.A1(\final_adder.p_new$416 ),
    .A2(\final_adder.g_new$421 ),
    .B1(\final_adder.g_new$417 ),
    .X(\final_adder.g_new$543 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$416  (.A(\final_adder.p_new$422 ),
    .B(\final_adder.p_new$418 ),
    .X(\final_adder.p_new$544 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$417  (.A1(\final_adder.p_new$418 ),
    .A2(\final_adder.g_new$423 ),
    .B1(\final_adder.g_new$419 ),
    .X(\final_adder.g_new$545 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$418  (.A(\final_adder.p_new$424 ),
    .B(\final_adder.p_new$420 ),
    .X(\final_adder.p_new$546 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$419  (.A1(\final_adder.p_new$420 ),
    .A2(\final_adder.g_new$425 ),
    .B1(\final_adder.g_new$421 ),
    .X(\final_adder.g_new$547 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$42  (.A(\c$4234 ),
    .B(\s$4237 ),
    .COUT(\final_adder.$signal$86 ),
    .SUM(\final_adder.$signal$1132 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$420  (.A(\final_adder.p_new$426 ),
    .B(\final_adder.p_new$422 ),
    .X(\final_adder.p_new$548 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$421  (.A1(\final_adder.p_new$422 ),
    .A2(\final_adder.g_new$427 ),
    .B1(\final_adder.g_new$423 ),
    .X(\final_adder.g_new$549 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$422  (.A(\final_adder.p_new$428 ),
    .B(\final_adder.p_new$424 ),
    .X(\final_adder.p_new$550 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$423  (.A1(\final_adder.p_new$424 ),
    .A2(\final_adder.g_new$429 ),
    .B1(\final_adder.g_new$425 ),
    .X(\final_adder.g_new$551 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$424  (.A(\final_adder.p_new$430 ),
    .B(\final_adder.p_new$426 ),
    .X(\final_adder.p_new$552 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$425  (.A1(\final_adder.p_new$426 ),
    .A2(\final_adder.g_new$431 ),
    .B1(\final_adder.g_new$427 ),
    .X(\final_adder.g_new$553 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$426  (.A(\final_adder.p_new$432 ),
    .B(\final_adder.p_new$428 ),
    .X(\final_adder.p_new$554 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$427  (.A1(\final_adder.p_new$428 ),
    .A2(\final_adder.g_new$433 ),
    .B1(\final_adder.g_new$429 ),
    .X(\final_adder.g_new$555 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$428  (.A(\final_adder.p_new$434 ),
    .B(\final_adder.p_new$430 ),
    .X(\final_adder.p_new$556 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$429  (.A1(\final_adder.p_new$430 ),
    .A2(\final_adder.g_new$435 ),
    .B1(\final_adder.g_new$431 ),
    .X(\final_adder.g_new$557 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$43  (.A(\c$4236 ),
    .B(\s$4239 ),
    .COUT(\final_adder.$signal$88 ),
    .SUM(\final_adder.$signal$1133 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$430  (.A(\final_adder.p_new$436 ),
    .B(\final_adder.p_new$432 ),
    .X(\final_adder.p_new$558 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$431  (.A1(\final_adder.p_new$432 ),
    .A2(\final_adder.g_new$437 ),
    .B1(\final_adder.g_new$433 ),
    .X(\final_adder.g_new$559 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$432  (.A(\final_adder.p_new$438 ),
    .B(\final_adder.p_new$434 ),
    .X(\final_adder.p_new$560 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$433  (.A1(\final_adder.p_new$434 ),
    .A2(\final_adder.g_new$439 ),
    .B1(\final_adder.g_new$435 ),
    .X(\final_adder.g_new$561 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$434  (.A(\final_adder.p_new$440 ),
    .B(\final_adder.p_new$436 ),
    .X(\final_adder.p_new$562 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$435  (.A1(\final_adder.p_new$436 ),
    .A2(\final_adder.g_new$441 ),
    .B1(\final_adder.g_new$437 ),
    .X(\final_adder.g_new$563 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$436  (.A(\final_adder.p_new$442 ),
    .B(\final_adder.p_new$438 ),
    .X(\final_adder.p_new$564 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$437  (.A1(\final_adder.p_new$438 ),
    .A2(\final_adder.g_new$443 ),
    .B1(\final_adder.g_new$439 ),
    .X(\final_adder.g_new$565 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$438  (.A(\final_adder.p_new$444 ),
    .B(\final_adder.p_new$440 ),
    .X(\final_adder.p_new$566 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$439  (.A1(\final_adder.p_new$440 ),
    .A2(\final_adder.g_new$445 ),
    .B1(\final_adder.g_new$441 ),
    .X(\final_adder.g_new$567 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$44  (.A(\c$4238 ),
    .B(\s$4241 ),
    .COUT(\final_adder.$signal$90 ),
    .SUM(\final_adder.$signal$1134 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$440  (.A(\final_adder.p_new$446 ),
    .B(\final_adder.p_new$442 ),
    .X(\final_adder.p_new$568 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$441  (.A1(\final_adder.p_new$442 ),
    .A2(\final_adder.g_new$447 ),
    .B1(\final_adder.g_new$443 ),
    .X(\final_adder.g_new$569 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$442  (.A(\final_adder.p_new$448 ),
    .B(\final_adder.p_new$444 ),
    .X(\final_adder.p_new$570 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$443  (.A1(\final_adder.p_new$444 ),
    .A2(\final_adder.g_new$449 ),
    .B1(\final_adder.g_new$445 ),
    .X(\final_adder.g_new$571 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$444  (.A(\final_adder.p_new$450 ),
    .B(\final_adder.p_new$446 ),
    .X(\final_adder.p_new$572 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$445  (.A1(\final_adder.p_new$446 ),
    .A2(\final_adder.g_new$451 ),
    .B1(\final_adder.g_new$447 ),
    .X(\final_adder.g_new$573 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$446  (.A(\final_adder.p_new$452 ),
    .B(\final_adder.p_new$448 ),
    .X(\final_adder.p_new$574 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$447  (.A1(\final_adder.p_new$448 ),
    .A2(\final_adder.g_new$453 ),
    .B1(\final_adder.g_new$449 ),
    .X(\final_adder.g_new$575 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$448  (.A(\final_adder.p_new$454 ),
    .B(\final_adder.p_new$450 ),
    .X(\final_adder.p_new$576 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$449  (.A1(\final_adder.p_new$450 ),
    .A2(\final_adder.g_new$455 ),
    .B1(\final_adder.g_new$451 ),
    .X(\final_adder.g_new$577 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$45  (.A(\c$4240 ),
    .B(\s$4243 ),
    .COUT(\final_adder.$signal$92 ),
    .SUM(\final_adder.$signal$1135 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$450  (.A(\final_adder.p_new$456 ),
    .B(\final_adder.p_new$452 ),
    .X(\final_adder.p_new$578 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$451  (.A1(\final_adder.p_new$452 ),
    .A2(\final_adder.g_new$457 ),
    .B1(\final_adder.g_new$453 ),
    .X(\final_adder.g_new$579 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$452  (.A(\final_adder.p_new$458 ),
    .B(\final_adder.p_new$454 ),
    .X(\final_adder.p_new$580 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$453  (.A1(\final_adder.p_new$454 ),
    .A2(\final_adder.g_new$459 ),
    .B1(\final_adder.g_new$455 ),
    .X(\final_adder.g_new$581 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$454  (.A(\final_adder.p_new$460 ),
    .B(\final_adder.p_new$456 ),
    .X(\final_adder.p_new$582 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$455  (.A1(\final_adder.p_new$456 ),
    .A2(\final_adder.g_new$461 ),
    .B1(\final_adder.g_new$457 ),
    .X(\final_adder.g_new$583 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$456  (.A(\final_adder.p_new$462 ),
    .B(\final_adder.p_new$458 ),
    .X(\final_adder.p_new$584 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$457  (.A1(\final_adder.p_new$458 ),
    .A2(\final_adder.g_new$463 ),
    .B1(\final_adder.g_new$459 ),
    .X(\final_adder.g_new$585 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$458  (.A(\final_adder.p_new$464 ),
    .B(\final_adder.p_new$460 ),
    .X(\final_adder.p_new$586 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$459  (.A1(\final_adder.p_new$460 ),
    .A2(\final_adder.g_new$465 ),
    .B1(\final_adder.g_new$461 ),
    .X(\final_adder.g_new$587 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$46  (.A(\c$4242 ),
    .B(\s$4245 ),
    .COUT(\final_adder.$signal$94 ),
    .SUM(\final_adder.$signal$1136 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$460  (.A(\final_adder.p_new$466 ),
    .B(\final_adder.p_new$462 ),
    .X(\final_adder.p_new$588 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$461  (.A1(\final_adder.p_new$462 ),
    .A2(\final_adder.g_new$467 ),
    .B1(\final_adder.g_new$463 ),
    .X(\final_adder.g_new$589 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$462  (.A(\final_adder.p_new$468 ),
    .B(\final_adder.p_new$464 ),
    .X(\final_adder.p_new$590 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$463  (.A1(\final_adder.p_new$464 ),
    .A2(\final_adder.g_new$469 ),
    .B1(\final_adder.g_new$465 ),
    .X(\final_adder.g_new$591 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$464  (.A(\final_adder.p_new$470 ),
    .B(\final_adder.p_new$466 ),
    .X(\final_adder.p_new$592 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$465  (.A1(\final_adder.p_new$466 ),
    .A2(\final_adder.g_new$471 ),
    .B1(\final_adder.g_new$467 ),
    .X(\final_adder.g_new$593 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$466  (.A(\final_adder.p_new$472 ),
    .B(\final_adder.p_new$468 ),
    .X(\final_adder.p_new$594 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$467  (.A1(\final_adder.p_new$468 ),
    .A2(\final_adder.g_new$473 ),
    .B1(\final_adder.g_new$469 ),
    .X(\final_adder.g_new$595 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$468  (.A(\final_adder.p_new$474 ),
    .B(\final_adder.p_new$470 ),
    .X(\final_adder.p_new$596 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$469  (.A1(\final_adder.p_new$470 ),
    .A2(\final_adder.g_new$475 ),
    .B1(\final_adder.g_new$471 ),
    .X(\final_adder.g_new$597 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$47  (.A(\c$4244 ),
    .B(\s$4247 ),
    .COUT(\final_adder.$signal$96 ),
    .SUM(\final_adder.$signal$1137 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$470  (.A(\final_adder.p_new$476 ),
    .B(\final_adder.p_new$472 ),
    .X(\final_adder.p_new$598 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$471  (.A1(\final_adder.p_new$472 ),
    .A2(\final_adder.g_new$477 ),
    .B1(\final_adder.g_new$473 ),
    .X(\final_adder.g_new$599 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$472  (.A(\final_adder.p_new$478 ),
    .B(\final_adder.p_new$474 ),
    .X(\final_adder.p_new$600 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$473  (.A1(\final_adder.p_new$474 ),
    .A2(\final_adder.g_new$479 ),
    .B1(\final_adder.g_new$475 ),
    .X(\final_adder.g_new$601 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$474  (.A(\final_adder.p_new$480 ),
    .B(\final_adder.p_new$476 ),
    .X(\final_adder.p_new$602 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$475  (.A1(\final_adder.p_new$476 ),
    .A2(\final_adder.g_new$481 ),
    .B1(\final_adder.g_new$477 ),
    .X(\final_adder.g_new$603 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$476  (.A(\final_adder.p_new$482 ),
    .B(\final_adder.p_new$478 ),
    .X(\final_adder.p_new$604 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$477  (.A1(\final_adder.p_new$478 ),
    .A2(\final_adder.g_new$483 ),
    .B1(\final_adder.g_new$479 ),
    .X(\final_adder.g_new$605 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$478  (.A(\final_adder.p_new$484 ),
    .B(\final_adder.p_new$480 ),
    .X(\final_adder.p_new$606 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$479  (.A1(\final_adder.p_new$480 ),
    .A2(\final_adder.g_new$485 ),
    .B1(\final_adder.g_new$481 ),
    .X(\final_adder.g_new$607 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$48  (.A(\c$4246 ),
    .B(\s$4249 ),
    .COUT(\final_adder.$signal$98 ),
    .SUM(\final_adder.$signal$1138 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$480  (.A(\final_adder.p_new$486 ),
    .B(\final_adder.p_new$482 ),
    .X(\final_adder.p_new$608 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$481  (.A1(\final_adder.p_new$482 ),
    .A2(\final_adder.g_new$487 ),
    .B1(\final_adder.g_new$483 ),
    .X(\final_adder.g_new$609 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$482  (.A(\final_adder.p_new$488 ),
    .B(\final_adder.p_new$484 ),
    .X(\final_adder.p_new$610 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$483  (.A1(\final_adder.p_new$484 ),
    .A2(\final_adder.g_new$489 ),
    .B1(\final_adder.g_new$485 ),
    .X(\final_adder.g_new$611 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$484  (.A(\final_adder.p_new$490 ),
    .B(\final_adder.p_new$486 ),
    .X(\final_adder.p_new$612 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$485  (.A1(\final_adder.p_new$486 ),
    .A2(\final_adder.g_new$491 ),
    .B1(\final_adder.g_new$487 ),
    .X(\final_adder.g_new$613 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$486  (.A(\final_adder.p_new$492 ),
    .B(\final_adder.p_new$488 ),
    .X(\final_adder.p_new$614 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$487  (.A1(\final_adder.p_new$488 ),
    .A2(\final_adder.g_new$493 ),
    .B1(\final_adder.g_new$489 ),
    .X(\final_adder.g_new$615 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$488  (.A(\final_adder.p_new$494 ),
    .B(\final_adder.p_new$490 ),
    .X(\final_adder.p_new$616 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$489  (.A1(\final_adder.p_new$490 ),
    .A2(\final_adder.g_new$495 ),
    .B1(\final_adder.g_new$491 ),
    .X(\final_adder.g_new$617 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$49  (.A(\c$4248 ),
    .B(\s$4251 ),
    .COUT(\final_adder.$signal$100 ),
    .SUM(\final_adder.$signal$101 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$490  (.A(\final_adder.p_new$496 ),
    .B(\final_adder.p_new$492 ),
    .X(\final_adder.p_new$618 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$491  (.A1(\final_adder.p_new$492 ),
    .A2(\final_adder.g_new$497 ),
    .B1(\final_adder.g_new$493 ),
    .X(\final_adder.g_new$619 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$492  (.A(\final_adder.p_new$498 ),
    .B(\final_adder.p_new$494 ),
    .X(\final_adder.p_new$620 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$493  (.A1(\final_adder.p_new$494 ),
    .A2(\final_adder.g_new$499 ),
    .B1(\final_adder.g_new$495 ),
    .X(\final_adder.g_new$621 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$494  (.A(\final_adder.p_new$500 ),
    .B(\final_adder.p_new$496 ),
    .X(\final_adder.p_new$622 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$495  (.A1(\final_adder.p_new$496 ),
    .A2(\final_adder.g_new$501 ),
    .B1(\final_adder.g_new$497 ),
    .X(\final_adder.g_new$623 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$496  (.A(\final_adder.p_new$502 ),
    .B(\final_adder.p_new$498 ),
    .X(\final_adder.p_new$624 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$497  (.A1(\final_adder.p_new$498 ),
    .A2(\final_adder.g_new$503 ),
    .B1(\final_adder.g_new$499 ),
    .X(\final_adder.g_new$625 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$498  (.A(\final_adder.p_new$504 ),
    .B(\final_adder.p_new$500 ),
    .X(\final_adder.p_new$626 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$499  (.A1(\final_adder.p_new$500 ),
    .A2(\final_adder.g_new$505 ),
    .B1(\final_adder.g_new$501 ),
    .X(\final_adder.g_new$627 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$5  (.A(\c$4160 ),
    .B(\s$4163 ),
    .COUT(\final_adder.$signal$12 ),
    .SUM(\final_adder.$signal$1095 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$50  (.A(\c$4250 ),
    .B(\s$4253 ),
    .COUT(\final_adder.$signal$102 ),
    .SUM(\final_adder.$signal$103 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$500  (.A(\final_adder.p_new$506 ),
    .B(\final_adder.p_new$502 ),
    .X(\final_adder.p_new$628 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$501  (.A1(\final_adder.p_new$502 ),
    .A2(\final_adder.g_new$507 ),
    .B1(\final_adder.g_new$503 ),
    .X(\final_adder.g_new$629 ));
 sky130_fd_sc_hd__a21o_4 \final_adder.U$$503  (.A1(\final_adder.p_new$504 ),
    .A2(\final_adder.g_new$509 ),
    .B1(\final_adder.g_new$505 ),
    .X(\final_adder.g_new$631 ));
 sky130_fd_sc_hd__a21o_4 \final_adder.U$$505  (.A1(\final_adder.p_new$506 ),
    .A2(\final_adder.g_new$383 ),
    .B1(\final_adder.g_new$507 ),
    .X(\final_adder.g_new$633 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$508  (.A(\final_adder.p_new$520 ),
    .B(\final_adder.p_new$512 ),
    .X(\final_adder.p_new$636 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$509  (.A1(\final_adder.p_new$512 ),
    .A2(\final_adder.g_new$521 ),
    .B1(\final_adder.g_new$513 ),
    .X(\final_adder.g_new$637 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$51  (.A(\c$4252 ),
    .B(\s$4255 ),
    .COUT(\final_adder.$signal$104 ),
    .SUM(\final_adder.$signal$105 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$510  (.A(\final_adder.p_new$522 ),
    .B(\final_adder.p_new$514 ),
    .X(\final_adder.p_new$638 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$511  (.A1(\final_adder.p_new$514 ),
    .A2(\final_adder.g_new$523 ),
    .B1(\final_adder.g_new$515 ),
    .X(\final_adder.g_new$639 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$512  (.A(\final_adder.p_new$524 ),
    .B(\final_adder.p_new$516 ),
    .X(\final_adder.p_new$640 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$513  (.A1(\final_adder.p_new$516 ),
    .A2(\final_adder.g_new$525 ),
    .B1(\final_adder.g_new$517 ),
    .X(\final_adder.g_new$641 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$514  (.A(\final_adder.p_new$526 ),
    .B(\final_adder.p_new$518 ),
    .X(\final_adder.p_new$642 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$515  (.A1(\final_adder.p_new$518 ),
    .A2(\final_adder.g_new$527 ),
    .B1(\final_adder.g_new$519 ),
    .X(\final_adder.g_new$643 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$516  (.A(\final_adder.p_new$528 ),
    .B(\final_adder.p_new$520 ),
    .X(\final_adder.p_new$644 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$517  (.A1(\final_adder.p_new$520 ),
    .A2(\final_adder.g_new$529 ),
    .B1(\final_adder.g_new$521 ),
    .X(\final_adder.g_new$645 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$518  (.A(\final_adder.p_new$530 ),
    .B(\final_adder.p_new$522 ),
    .X(\final_adder.p_new$646 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$519  (.A1(\final_adder.p_new$522 ),
    .A2(\final_adder.g_new$531 ),
    .B1(\final_adder.g_new$523 ),
    .X(\final_adder.g_new$647 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$52  (.A(\c$4254 ),
    .B(\s$4257 ),
    .COUT(\final_adder.$signal$106 ),
    .SUM(\final_adder.$signal$107 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$520  (.A(\final_adder.p_new$532 ),
    .B(\final_adder.p_new$524 ),
    .X(\final_adder.p_new$648 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$521  (.A1(\final_adder.p_new$524 ),
    .A2(\final_adder.g_new$533 ),
    .B1(\final_adder.g_new$525 ),
    .X(\final_adder.g_new$649 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$522  (.A(\final_adder.p_new$534 ),
    .B(\final_adder.p_new$526 ),
    .X(\final_adder.p_new$650 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$523  (.A1(\final_adder.p_new$526 ),
    .A2(\final_adder.g_new$535 ),
    .B1(\final_adder.g_new$527 ),
    .X(\final_adder.g_new$651 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$524  (.A(\final_adder.p_new$536 ),
    .B(\final_adder.p_new$528 ),
    .X(\final_adder.p_new$652 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$525  (.A1(\final_adder.p_new$528 ),
    .A2(\final_adder.g_new$537 ),
    .B1(\final_adder.g_new$529 ),
    .X(\final_adder.g_new$653 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$526  (.A(\final_adder.p_new$538 ),
    .B(\final_adder.p_new$530 ),
    .X(\final_adder.p_new$654 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$527  (.A1(\final_adder.p_new$530 ),
    .A2(\final_adder.g_new$539 ),
    .B1(\final_adder.g_new$531 ),
    .X(\final_adder.g_new$655 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$528  (.A(\final_adder.p_new$540 ),
    .B(\final_adder.p_new$532 ),
    .X(\final_adder.p_new$656 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$529  (.A1(\final_adder.p_new$532 ),
    .A2(\final_adder.g_new$541 ),
    .B1(\final_adder.g_new$533 ),
    .X(\final_adder.g_new$657 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$53  (.A(\c$4256 ),
    .B(\s$4259 ),
    .COUT(\final_adder.$signal$108 ),
    .SUM(\final_adder.$signal$109 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$530  (.A(\final_adder.p_new$542 ),
    .B(\final_adder.p_new$534 ),
    .X(\final_adder.p_new$658 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$531  (.A1(\final_adder.p_new$534 ),
    .A2(\final_adder.g_new$543 ),
    .B1(\final_adder.g_new$535 ),
    .X(\final_adder.g_new$659 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$532  (.A(\final_adder.p_new$544 ),
    .B(\final_adder.p_new$536 ),
    .X(\final_adder.p_new$660 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$533  (.A1(\final_adder.p_new$536 ),
    .A2(\final_adder.g_new$545 ),
    .B1(\final_adder.g_new$537 ),
    .X(\final_adder.g_new$661 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$534  (.A(\final_adder.p_new$546 ),
    .B(\final_adder.p_new$538 ),
    .X(\final_adder.p_new$662 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$535  (.A1(\final_adder.p_new$538 ),
    .A2(\final_adder.g_new$547 ),
    .B1(\final_adder.g_new$539 ),
    .X(\final_adder.g_new$663 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$536  (.A(\final_adder.p_new$548 ),
    .B(\final_adder.p_new$540 ),
    .X(\final_adder.p_new$664 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$537  (.A1(\final_adder.p_new$540 ),
    .A2(\final_adder.g_new$549 ),
    .B1(\final_adder.g_new$541 ),
    .X(\final_adder.g_new$665 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$538  (.A(\final_adder.p_new$550 ),
    .B(\final_adder.p_new$542 ),
    .X(\final_adder.p_new$666 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$539  (.A1(\final_adder.p_new$542 ),
    .A2(\final_adder.g_new$551 ),
    .B1(\final_adder.g_new$543 ),
    .X(\final_adder.g_new$667 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$54  (.A(\c$4258 ),
    .B(\s$4261 ),
    .COUT(\final_adder.$signal$110 ),
    .SUM(\final_adder.$signal$111 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$540  (.A(\final_adder.p_new$552 ),
    .B(\final_adder.p_new$544 ),
    .X(\final_adder.p_new$668 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$541  (.A1(\final_adder.p_new$544 ),
    .A2(\final_adder.g_new$553 ),
    .B1(\final_adder.g_new$545 ),
    .X(\final_adder.g_new$669 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$542  (.A(\final_adder.p_new$554 ),
    .B(\final_adder.p_new$546 ),
    .X(\final_adder.p_new$670 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$543  (.A1(\final_adder.p_new$546 ),
    .A2(\final_adder.g_new$555 ),
    .B1(\final_adder.g_new$547 ),
    .X(\final_adder.g_new$671 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$544  (.A(\final_adder.p_new$556 ),
    .B(\final_adder.p_new$548 ),
    .X(\final_adder.p_new$672 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$545  (.A1(\final_adder.p_new$548 ),
    .A2(\final_adder.g_new$557 ),
    .B1(\final_adder.g_new$549 ),
    .X(\final_adder.g_new$673 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$546  (.A(\final_adder.p_new$558 ),
    .B(\final_adder.p_new$550 ),
    .X(\final_adder.p_new$674 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$547  (.A1(\final_adder.p_new$550 ),
    .A2(\final_adder.g_new$559 ),
    .B1(\final_adder.g_new$551 ),
    .X(\final_adder.g_new$675 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$548  (.A(\final_adder.p_new$560 ),
    .B(\final_adder.p_new$552 ),
    .X(\final_adder.p_new$676 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$549  (.A1(\final_adder.p_new$552 ),
    .A2(\final_adder.g_new$561 ),
    .B1(\final_adder.g_new$553 ),
    .X(\final_adder.g_new$677 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$55  (.A(\c$4260 ),
    .B(\s$4263 ),
    .COUT(\final_adder.$signal$112 ),
    .SUM(\final_adder.$signal$113 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$550  (.A(\final_adder.p_new$562 ),
    .B(\final_adder.p_new$554 ),
    .X(\final_adder.p_new$678 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$551  (.A1(\final_adder.p_new$554 ),
    .A2(\final_adder.g_new$563 ),
    .B1(\final_adder.g_new$555 ),
    .X(\final_adder.g_new$679 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$552  (.A(\final_adder.p_new$564 ),
    .B(\final_adder.p_new$556 ),
    .X(\final_adder.p_new$680 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$553  (.A1(\final_adder.p_new$556 ),
    .A2(\final_adder.g_new$565 ),
    .B1(\final_adder.g_new$557 ),
    .X(\final_adder.g_new$681 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$554  (.A(\final_adder.p_new$566 ),
    .B(\final_adder.p_new$558 ),
    .X(\final_adder.p_new$682 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$555  (.A1(\final_adder.p_new$558 ),
    .A2(\final_adder.g_new$567 ),
    .B1(\final_adder.g_new$559 ),
    .X(\final_adder.g_new$683 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$556  (.A(\final_adder.p_new$568 ),
    .B(\final_adder.p_new$560 ),
    .X(\final_adder.p_new$684 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$557  (.A1(\final_adder.p_new$560 ),
    .A2(\final_adder.g_new$569 ),
    .B1(\final_adder.g_new$561 ),
    .X(\final_adder.g_new$685 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$558  (.A(\final_adder.p_new$570 ),
    .B(\final_adder.p_new$562 ),
    .X(\final_adder.p_new$686 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$559  (.A1(\final_adder.p_new$562 ),
    .A2(\final_adder.g_new$571 ),
    .B1(\final_adder.g_new$563 ),
    .X(\final_adder.g_new$687 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$56  (.A(\c$4262 ),
    .B(\s$4265 ),
    .COUT(\final_adder.$signal$114 ),
    .SUM(\final_adder.$signal$1146 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$560  (.A(\final_adder.p_new$572 ),
    .B(\final_adder.p_new$564 ),
    .X(\final_adder.p_new$688 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$561  (.A1(\final_adder.p_new$564 ),
    .A2(\final_adder.g_new$573 ),
    .B1(\final_adder.g_new$565 ),
    .X(\final_adder.g_new$689 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$562  (.A(\final_adder.p_new$574 ),
    .B(\final_adder.p_new$566 ),
    .X(\final_adder.p_new$690 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$563  (.A1(\final_adder.p_new$566 ),
    .A2(\final_adder.g_new$575 ),
    .B1(\final_adder.g_new$567 ),
    .X(\final_adder.g_new$691 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$564  (.A(\final_adder.p_new$576 ),
    .B(\final_adder.p_new$568 ),
    .X(\final_adder.p_new$692 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$565  (.A1(\final_adder.p_new$568 ),
    .A2(\final_adder.g_new$577 ),
    .B1(\final_adder.g_new$569 ),
    .X(\final_adder.g_new$693 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$566  (.A(\final_adder.p_new$578 ),
    .B(\final_adder.p_new$570 ),
    .X(\final_adder.p_new$694 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$567  (.A1(\final_adder.p_new$570 ),
    .A2(\final_adder.g_new$579 ),
    .B1(\final_adder.g_new$571 ),
    .X(\final_adder.g_new$695 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$568  (.A(\final_adder.p_new$580 ),
    .B(\final_adder.p_new$572 ),
    .X(\final_adder.p_new$696 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$569  (.A1(\final_adder.p_new$572 ),
    .A2(\final_adder.g_new$581 ),
    .B1(\final_adder.g_new$573 ),
    .X(\final_adder.g_new$697 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$57  (.A(\c$4264 ),
    .B(\s$4267 ),
    .COUT(\final_adder.$signal$116 ),
    .SUM(\final_adder.$signal$1147 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$570  (.A(\final_adder.p_new$582 ),
    .B(\final_adder.p_new$574 ),
    .X(\final_adder.p_new$698 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$571  (.A1(\final_adder.p_new$574 ),
    .A2(\final_adder.g_new$583 ),
    .B1(\final_adder.g_new$575 ),
    .X(\final_adder.g_new$699 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$572  (.A(\final_adder.p_new$584 ),
    .B(\final_adder.p_new$576 ),
    .X(\final_adder.p_new$700 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$573  (.A1(\final_adder.p_new$576 ),
    .A2(\final_adder.g_new$585 ),
    .B1(\final_adder.g_new$577 ),
    .X(\final_adder.g_new$701 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$574  (.A(\final_adder.p_new$586 ),
    .B(\final_adder.p_new$578 ),
    .X(\final_adder.p_new$702 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$575  (.A1(\final_adder.p_new$578 ),
    .A2(\final_adder.g_new$587 ),
    .B1(\final_adder.g_new$579 ),
    .X(\final_adder.g_new$703 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$576  (.A(\final_adder.p_new$588 ),
    .B(\final_adder.p_new$580 ),
    .X(\final_adder.p_new$704 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$577  (.A1(\final_adder.p_new$580 ),
    .A2(\final_adder.g_new$589 ),
    .B1(\final_adder.g_new$581 ),
    .X(\final_adder.g_new$705 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$578  (.A(\final_adder.p_new$590 ),
    .B(\final_adder.p_new$582 ),
    .X(\final_adder.p_new$706 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$579  (.A1(\final_adder.p_new$582 ),
    .A2(\final_adder.g_new$591 ),
    .B1(\final_adder.g_new$583 ),
    .X(\final_adder.g_new$707 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$58  (.A(\c$4266 ),
    .B(\s$4269 ),
    .COUT(\final_adder.$signal$118 ),
    .SUM(\final_adder.$signal$1148 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$580  (.A(\final_adder.p_new$592 ),
    .B(\final_adder.p_new$584 ),
    .X(\final_adder.p_new$708 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$581  (.A1(\final_adder.p_new$584 ),
    .A2(\final_adder.g_new$593 ),
    .B1(\final_adder.g_new$585 ),
    .X(\final_adder.g_new$709 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$582  (.A(\final_adder.p_new$594 ),
    .B(\final_adder.p_new$586 ),
    .X(\final_adder.p_new$710 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$583  (.A1(\final_adder.p_new$586 ),
    .A2(\final_adder.g_new$595 ),
    .B1(\final_adder.g_new$587 ),
    .X(\final_adder.g_new$711 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$584  (.A(\final_adder.p_new$596 ),
    .B(\final_adder.p_new$588 ),
    .X(\final_adder.p_new$712 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$585  (.A1(\final_adder.p_new$588 ),
    .A2(\final_adder.g_new$597 ),
    .B1(\final_adder.g_new$589 ),
    .X(\final_adder.g_new$713 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$586  (.A(\final_adder.p_new$598 ),
    .B(\final_adder.p_new$590 ),
    .X(\final_adder.p_new$714 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$587  (.A1(\final_adder.p_new$590 ),
    .A2(\final_adder.g_new$599 ),
    .B1(\final_adder.g_new$591 ),
    .X(\final_adder.g_new$715 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$588  (.A(\final_adder.p_new$600 ),
    .B(\final_adder.p_new$592 ),
    .X(\final_adder.p_new$716 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$589  (.A1(\final_adder.p_new$592 ),
    .A2(\final_adder.g_new$601 ),
    .B1(\final_adder.g_new$593 ),
    .X(\final_adder.g_new$717 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$59  (.A(\c$4268 ),
    .B(\s$4271 ),
    .COUT(\final_adder.$signal$120 ),
    .SUM(\final_adder.$signal$1149 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$590  (.A(\final_adder.p_new$602 ),
    .B(\final_adder.p_new$594 ),
    .X(\final_adder.p_new$718 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$591  (.A1(\final_adder.p_new$594 ),
    .A2(\final_adder.g_new$603 ),
    .B1(\final_adder.g_new$595 ),
    .X(\final_adder.g_new$719 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$592  (.A(\final_adder.p_new$604 ),
    .B(\final_adder.p_new$596 ),
    .X(\final_adder.p_new$720 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$593  (.A1(\final_adder.p_new$596 ),
    .A2(\final_adder.g_new$605 ),
    .B1(\final_adder.g_new$597 ),
    .X(\final_adder.g_new$721 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$594  (.A(\final_adder.p_new$606 ),
    .B(\final_adder.p_new$598 ),
    .X(\final_adder.p_new$722 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$595  (.A1(\final_adder.p_new$598 ),
    .A2(\final_adder.g_new$607 ),
    .B1(\final_adder.g_new$599 ),
    .X(\final_adder.g_new$723 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$596  (.A(\final_adder.p_new$608 ),
    .B(\final_adder.p_new$600 ),
    .X(\final_adder.p_new$724 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$597  (.A1(\final_adder.p_new$600 ),
    .A2(\final_adder.g_new$609 ),
    .B1(\final_adder.g_new$601 ),
    .X(\final_adder.g_new$725 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$598  (.A(\final_adder.p_new$610 ),
    .B(\final_adder.p_new$602 ),
    .X(\final_adder.p_new$726 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$599  (.A1(\final_adder.p_new$602 ),
    .A2(\final_adder.g_new$611 ),
    .B1(\final_adder.g_new$603 ),
    .X(\final_adder.g_new$727 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$6  (.A(\c$4162 ),
    .B(\s$4165 ),
    .COUT(\final_adder.$signal$14 ),
    .SUM(\final_adder.$signal$1096 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$60  (.A(\c$4270 ),
    .B(\s$4273 ),
    .COUT(\final_adder.$signal$122 ),
    .SUM(\final_adder.$signal$1150 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$600  (.A(\final_adder.p_new$612 ),
    .B(\final_adder.p_new$604 ),
    .X(\final_adder.p_new$728 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$601  (.A1(\final_adder.p_new$604 ),
    .A2(\final_adder.g_new$613 ),
    .B1(\final_adder.g_new$605 ),
    .X(\final_adder.g_new$729 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$602  (.A(\final_adder.p_new$614 ),
    .B(\final_adder.p_new$606 ),
    .X(\final_adder.p_new$730 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$603  (.A1(\final_adder.p_new$606 ),
    .A2(\final_adder.g_new$615 ),
    .B1(\final_adder.g_new$607 ),
    .X(\final_adder.g_new$731 ));
 sky130_fd_sc_hd__and2_2 \final_adder.U$$604  (.A(\final_adder.p_new$616 ),
    .B(\final_adder.p_new$608 ),
    .X(\final_adder.p_new$732 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$605  (.A1(\final_adder.p_new$608 ),
    .A2(\final_adder.g_new$617 ),
    .B1(\final_adder.g_new$609 ),
    .X(\final_adder.g_new$733 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$606  (.A(\final_adder.p_new$618 ),
    .B(\final_adder.p_new$610 ),
    .X(\final_adder.p_new$734 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$607  (.A1(\final_adder.p_new$610 ),
    .A2(\final_adder.g_new$619 ),
    .B1(\final_adder.g_new$611 ),
    .X(\final_adder.g_new$735 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$608  (.A(\final_adder.p_new$620 ),
    .B(\final_adder.p_new$612 ),
    .X(\final_adder.p_new$736 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$609  (.A1(\final_adder.p_new$612 ),
    .A2(\final_adder.g_new$621 ),
    .B1(\final_adder.g_new$613 ),
    .X(\final_adder.g_new$737 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$61  (.A(\c$4272 ),
    .B(\s$4275 ),
    .COUT(\final_adder.$signal$124 ),
    .SUM(\final_adder.$signal$1151 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$610  (.A(\final_adder.p_new$622 ),
    .B(\final_adder.p_new$614 ),
    .X(\final_adder.p_new$738 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$611  (.A1(\final_adder.p_new$614 ),
    .A2(\final_adder.g_new$623 ),
    .B1(\final_adder.g_new$615 ),
    .X(\final_adder.g_new$739 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$612  (.A(\final_adder.p_new$624 ),
    .B(\final_adder.p_new$616 ),
    .X(\final_adder.p_new$740 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$613  (.A1(\final_adder.p_new$616 ),
    .A2(\final_adder.g_new$625 ),
    .B1(\final_adder.g_new$617 ),
    .X(\final_adder.g_new$741 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$614  (.A(\final_adder.p_new$626 ),
    .B(\final_adder.p_new$618 ),
    .X(\final_adder.p_new$742 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$615  (.A1(\final_adder.p_new$618 ),
    .A2(\final_adder.g_new$627 ),
    .B1(\final_adder.g_new$619 ),
    .X(\final_adder.g_new$743 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$616  (.A(\final_adder.p_new$628 ),
    .B(\final_adder.p_new$620 ),
    .X(\final_adder.p_new$744 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$617  (.A1(\final_adder.p_new$620 ),
    .A2(\final_adder.g_new$629 ),
    .B1(\final_adder.g_new$621 ),
    .X(\final_adder.g_new$745 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$619  (.A1(\final_adder.p_new$622 ),
    .A2(\final_adder.g_new$631 ),
    .B1(\final_adder.g_new$623 ),
    .X(\final_adder.g_new$747 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$62  (.A(\c$4274 ),
    .B(\s$4277 ),
    .COUT(\final_adder.$signal$126 ),
    .SUM(\final_adder.$signal$1152 ));
 sky130_fd_sc_hd__a21o_4 \final_adder.U$$621  (.A1(\final_adder.p_new$624 ),
    .A2(\final_adder.g_new$633 ),
    .B1(\final_adder.g_new$625 ),
    .X(\final_adder.g_new$749 ));
 sky130_fd_sc_hd__a21o_4 \final_adder.U$$623  (.A1(\final_adder.p_new$626 ),
    .A2(\final_adder.g_new$509 ),
    .B1(\final_adder.g_new$627 ),
    .X(\final_adder.g_new$751 ));
 sky130_fd_sc_hd__a21o_4 \final_adder.U$$625  (.A1(\final_adder.p_new$628 ),
    .A2(\final_adder.g_new$383 ),
    .B1(\final_adder.g_new$629 ),
    .X(\final_adder.g_new$753 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$628  (.A(\final_adder.p_new$652 ),
    .B(\final_adder.p_new$636 ),
    .X(\final_adder.p_new$756 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$629  (.A1(\final_adder.p_new$636 ),
    .A2(\final_adder.g_new$653 ),
    .B1(\final_adder.g_new$637 ),
    .X(\final_adder.g_new$757 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$63  (.A(\c$4276 ),
    .B(\s$4279 ),
    .COUT(\final_adder.$signal$128 ),
    .SUM(\final_adder.$signal$1153 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$630  (.A(\final_adder.p_new$654 ),
    .B(\final_adder.p_new$638 ),
    .X(\final_adder.p_new$758 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$631  (.A1(\final_adder.p_new$638 ),
    .A2(\final_adder.g_new$655 ),
    .B1(\final_adder.g_new$639 ),
    .X(\final_adder.g_new$759 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$632  (.A(\final_adder.p_new$656 ),
    .B(\final_adder.p_new$640 ),
    .X(\final_adder.p_new$760 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$633  (.A1(\final_adder.p_new$640 ),
    .A2(\final_adder.g_new$657 ),
    .B1(\final_adder.g_new$641 ),
    .X(\final_adder.g_new$761 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$634  (.A(\final_adder.p_new$658 ),
    .B(\final_adder.p_new$642 ),
    .X(\final_adder.p_new$762 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$635  (.A1(\final_adder.p_new$642 ),
    .A2(\final_adder.g_new$659 ),
    .B1(\final_adder.g_new$643 ),
    .X(\final_adder.g_new$763 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$636  (.A(\final_adder.p_new$660 ),
    .B(\final_adder.p_new$644 ),
    .X(\final_adder.p_new$764 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$637  (.A1(\final_adder.p_new$644 ),
    .A2(\final_adder.g_new$661 ),
    .B1(\final_adder.g_new$645 ),
    .X(\final_adder.g_new$765 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$638  (.A(\final_adder.p_new$662 ),
    .B(\final_adder.p_new$646 ),
    .X(\final_adder.p_new$766 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$639  (.A1(\final_adder.p_new$646 ),
    .A2(\final_adder.g_new$663 ),
    .B1(\final_adder.g_new$647 ),
    .X(\final_adder.g_new$767 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$64  (.A(\c$4278 ),
    .B(\s$4281 ),
    .COUT(\final_adder.$signal$130 ),
    .SUM(\final_adder.$signal$1154 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$640  (.A(\final_adder.p_new$664 ),
    .B(\final_adder.p_new$648 ),
    .X(\final_adder.p_new$768 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$641  (.A1(\final_adder.p_new$648 ),
    .A2(\final_adder.g_new$665 ),
    .B1(\final_adder.g_new$649 ),
    .X(\final_adder.g_new$769 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$642  (.A(\final_adder.p_new$666 ),
    .B(\final_adder.p_new$650 ),
    .X(\final_adder.p_new$770 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$643  (.A1(\final_adder.p_new$650 ),
    .A2(\final_adder.g_new$667 ),
    .B1(\final_adder.g_new$651 ),
    .X(\final_adder.g_new$771 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$644  (.A(\final_adder.p_new$668 ),
    .B(\final_adder.p_new$652 ),
    .X(\final_adder.p_new$772 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$645  (.A1(\final_adder.p_new$652 ),
    .A2(\final_adder.g_new$669 ),
    .B1(\final_adder.g_new$653 ),
    .X(\final_adder.g_new$773 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$646  (.A(\final_adder.p_new$670 ),
    .B(\final_adder.p_new$654 ),
    .X(\final_adder.p_new$774 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$647  (.A1(\final_adder.p_new$654 ),
    .A2(\final_adder.g_new$671 ),
    .B1(\final_adder.g_new$655 ),
    .X(\final_adder.g_new$775 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$648  (.A(\final_adder.p_new$672 ),
    .B(\final_adder.p_new$656 ),
    .X(\final_adder.p_new$776 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$649  (.A1(\final_adder.p_new$656 ),
    .A2(\final_adder.g_new$673 ),
    .B1(\final_adder.g_new$657 ),
    .X(\final_adder.g_new$777 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$65  (.A(\c$4280 ),
    .B(\s$4283 ),
    .COUT(\final_adder.$signal$132 ),
    .SUM(\final_adder.$signal$1155 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$650  (.A(\final_adder.p_new$674 ),
    .B(\final_adder.p_new$658 ),
    .X(\final_adder.p_new$778 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$651  (.A1(\final_adder.p_new$658 ),
    .A2(\final_adder.g_new$675 ),
    .B1(\final_adder.g_new$659 ),
    .X(\final_adder.g_new$779 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$652  (.A(\final_adder.p_new$676 ),
    .B(\final_adder.p_new$660 ),
    .X(\final_adder.p_new$780 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$653  (.A1(\final_adder.p_new$660 ),
    .A2(\final_adder.g_new$677 ),
    .B1(\final_adder.g_new$661 ),
    .X(\final_adder.g_new$781 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$654  (.A(\final_adder.p_new$678 ),
    .B(\final_adder.p_new$662 ),
    .X(\final_adder.p_new$782 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$655  (.A1(\final_adder.p_new$662 ),
    .A2(\final_adder.g_new$679 ),
    .B1(\final_adder.g_new$663 ),
    .X(\final_adder.g_new$783 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$656  (.A(\final_adder.p_new$680 ),
    .B(\final_adder.p_new$664 ),
    .X(\final_adder.p_new$784 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$657  (.A1(\final_adder.p_new$664 ),
    .A2(\final_adder.g_new$681 ),
    .B1(\final_adder.g_new$665 ),
    .X(\final_adder.g_new$785 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$658  (.A(\final_adder.p_new$682 ),
    .B(\final_adder.p_new$666 ),
    .X(\final_adder.p_new$786 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$659  (.A1(\final_adder.p_new$666 ),
    .A2(\final_adder.g_new$683 ),
    .B1(\final_adder.g_new$667 ),
    .X(\final_adder.g_new$787 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$66  (.A(\c$4282 ),
    .B(\s$4285 ),
    .COUT(\final_adder.$signal$134 ),
    .SUM(\final_adder.$signal$1156 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$660  (.A(\final_adder.p_new$684 ),
    .B(\final_adder.p_new$668 ),
    .X(\final_adder.p_new$788 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$661  (.A1(\final_adder.p_new$668 ),
    .A2(\final_adder.g_new$685 ),
    .B1(\final_adder.g_new$669 ),
    .X(\final_adder.g_new$789 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$662  (.A(\final_adder.p_new$686 ),
    .B(\final_adder.p_new$670 ),
    .X(\final_adder.p_new$790 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$663  (.A1(\final_adder.p_new$670 ),
    .A2(\final_adder.g_new$687 ),
    .B1(\final_adder.g_new$671 ),
    .X(\final_adder.g_new$791 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$664  (.A(\final_adder.p_new$688 ),
    .B(\final_adder.p_new$672 ),
    .X(\final_adder.p_new$792 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$665  (.A1(\final_adder.p_new$672 ),
    .A2(\final_adder.g_new$689 ),
    .B1(\final_adder.g_new$673 ),
    .X(\final_adder.g_new$793 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$666  (.A(\final_adder.p_new$690 ),
    .B(\final_adder.p_new$674 ),
    .X(\final_adder.p_new$794 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$667  (.A1(\final_adder.p_new$674 ),
    .A2(\final_adder.g_new$691 ),
    .B1(\final_adder.g_new$675 ),
    .X(\final_adder.g_new$795 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$668  (.A(\final_adder.p_new$692 ),
    .B(\final_adder.p_new$676 ),
    .X(\final_adder.p_new$796 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$669  (.A1(\final_adder.p_new$676 ),
    .A2(\final_adder.g_new$693 ),
    .B1(\final_adder.g_new$677 ),
    .X(\final_adder.g_new$797 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$67  (.A(\c$4284 ),
    .B(\s$4287 ),
    .COUT(\final_adder.$signal$136 ),
    .SUM(\final_adder.$signal$1157 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$670  (.A(\final_adder.p_new$694 ),
    .B(\final_adder.p_new$678 ),
    .X(\final_adder.p_new$798 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$671  (.A1(\final_adder.p_new$678 ),
    .A2(\final_adder.g_new$695 ),
    .B1(\final_adder.g_new$679 ),
    .X(\final_adder.g_new$799 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$672  (.A(\final_adder.p_new$696 ),
    .B(\final_adder.p_new$680 ),
    .X(\final_adder.p_new$800 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$673  (.A1(\final_adder.p_new$680 ),
    .A2(\final_adder.g_new$697 ),
    .B1(\final_adder.g_new$681 ),
    .X(\final_adder.g_new$801 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$674  (.A(\final_adder.p_new$698 ),
    .B(\final_adder.p_new$682 ),
    .X(\final_adder.p_new$802 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$675  (.A1(\final_adder.p_new$682 ),
    .A2(\final_adder.g_new$699 ),
    .B1(\final_adder.g_new$683 ),
    .X(\final_adder.g_new$803 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$676  (.A(\final_adder.p_new$700 ),
    .B(\final_adder.p_new$684 ),
    .X(\final_adder.p_new$804 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$677  (.A1(\final_adder.p_new$684 ),
    .A2(\final_adder.g_new$701 ),
    .B1(\final_adder.g_new$685 ),
    .X(\final_adder.g_new$805 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$678  (.A(\final_adder.p_new$702 ),
    .B(\final_adder.p_new$686 ),
    .X(\final_adder.p_new$806 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$679  (.A1(\final_adder.p_new$686 ),
    .A2(\final_adder.g_new$703 ),
    .B1(\final_adder.g_new$687 ),
    .X(\final_adder.g_new$807 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$68  (.A(\c$4286 ),
    .B(\s$4289 ),
    .COUT(\final_adder.$signal$138 ),
    .SUM(\final_adder.$signal$1158 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$680  (.A(\final_adder.p_new$704 ),
    .B(\final_adder.p_new$688 ),
    .X(\final_adder.p_new$808 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$681  (.A1(\final_adder.p_new$688 ),
    .A2(\final_adder.g_new$705 ),
    .B1(\final_adder.g_new$689 ),
    .X(\final_adder.g_new$809 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$682  (.A(\final_adder.p_new$706 ),
    .B(\final_adder.p_new$690 ),
    .X(\final_adder.p_new$810 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$683  (.A1(\final_adder.p_new$690 ),
    .A2(\final_adder.g_new$707 ),
    .B1(\final_adder.g_new$691 ),
    .X(\final_adder.g_new$811 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$684  (.A(\final_adder.p_new$708 ),
    .B(\final_adder.p_new$692 ),
    .X(\final_adder.p_new$812 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$685  (.A1(\final_adder.p_new$692 ),
    .A2(\final_adder.g_new$709 ),
    .B1(\final_adder.g_new$693 ),
    .X(\final_adder.g_new$813 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$686  (.A(\final_adder.p_new$710 ),
    .B(\final_adder.p_new$694 ),
    .X(\final_adder.p_new$814 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$687  (.A1(\final_adder.p_new$694 ),
    .A2(\final_adder.g_new$711 ),
    .B1(\final_adder.g_new$695 ),
    .X(\final_adder.g_new$815 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$688  (.A(\final_adder.p_new$712 ),
    .B(\final_adder.p_new$696 ),
    .X(\final_adder.p_new$816 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$689  (.A1(\final_adder.p_new$696 ),
    .A2(\final_adder.g_new$713 ),
    .B1(\final_adder.g_new$697 ),
    .X(\final_adder.g_new$817 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$69  (.A(\c$4288 ),
    .B(\s$4291 ),
    .COUT(\final_adder.$signal$140 ),
    .SUM(\final_adder.$signal$1159 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$690  (.A(\final_adder.p_new$714 ),
    .B(\final_adder.p_new$698 ),
    .X(\final_adder.p_new$818 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$691  (.A1(\final_adder.p_new$698 ),
    .A2(\final_adder.g_new$715 ),
    .B1(\final_adder.g_new$699 ),
    .X(\final_adder.g_new$819 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$692  (.A(\final_adder.p_new$716 ),
    .B(\final_adder.p_new$700 ),
    .X(\final_adder.p_new$820 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$693  (.A1(\final_adder.p_new$700 ),
    .A2(\final_adder.g_new$717 ),
    .B1(\final_adder.g_new$701 ),
    .X(\final_adder.g_new$821 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$694  (.A(\final_adder.p_new$718 ),
    .B(\final_adder.p_new$702 ),
    .X(\final_adder.p_new$822 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$695  (.A1(\final_adder.p_new$702 ),
    .A2(\final_adder.g_new$719 ),
    .B1(\final_adder.g_new$703 ),
    .X(\final_adder.g_new$823 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$696  (.A(\final_adder.p_new$720 ),
    .B(\final_adder.p_new$704 ),
    .X(\final_adder.p_new$824 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$697  (.A1(\final_adder.p_new$704 ),
    .A2(\final_adder.g_new$721 ),
    .B1(\final_adder.g_new$705 ),
    .X(\final_adder.g_new$825 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$698  (.A(\final_adder.p_new$722 ),
    .B(\final_adder.p_new$706 ),
    .X(\final_adder.p_new$826 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$699  (.A1(\final_adder.p_new$706 ),
    .A2(\final_adder.g_new$723 ),
    .B1(\final_adder.g_new$707 ),
    .X(\final_adder.g_new$827 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$7  (.A(\c$4164 ),
    .B(\s$4167 ),
    .COUT(\final_adder.$signal$16 ),
    .SUM(\final_adder.$signal$1097 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$70  (.A(\c$4290 ),
    .B(\s$4293 ),
    .COUT(\final_adder.$signal$142 ),
    .SUM(\final_adder.$signal$1160 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$700  (.A(\final_adder.p_new$724 ),
    .B(\final_adder.p_new$708 ),
    .X(\final_adder.p_new$828 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$701  (.A1(\final_adder.p_new$708 ),
    .A2(\final_adder.g_new$725 ),
    .B1(\final_adder.g_new$709 ),
    .X(\final_adder.g_new$829 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$702  (.A(\final_adder.p_new$726 ),
    .B(\final_adder.p_new$710 ),
    .X(\final_adder.p_new$830 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$703  (.A1(\final_adder.p_new$710 ),
    .A2(\final_adder.g_new$727 ),
    .B1(\final_adder.g_new$711 ),
    .X(\final_adder.g_new$831 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$704  (.A(\final_adder.p_new$728 ),
    .B(\final_adder.p_new$712 ),
    .X(\final_adder.p_new$832 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$705  (.A1(\final_adder.p_new$712 ),
    .A2(\final_adder.g_new$729 ),
    .B1(\final_adder.g_new$713 ),
    .X(\final_adder.g_new$833 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$706  (.A(\final_adder.p_new$730 ),
    .B(\final_adder.p_new$714 ),
    .X(\final_adder.p_new$834 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$707  (.A1(\final_adder.p_new$714 ),
    .A2(\final_adder.g_new$731 ),
    .B1(\final_adder.g_new$715 ),
    .X(\final_adder.g_new$835 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$708  (.A(\final_adder.p_new$732 ),
    .B(\final_adder.p_new$716 ),
    .X(\final_adder.p_new$836 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$709  (.A1(\final_adder.p_new$716 ),
    .A2(\final_adder.g_new$733 ),
    .B1(\final_adder.g_new$717 ),
    .X(\final_adder.g_new$837 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$71  (.A(\c$4292 ),
    .B(\s$4295 ),
    .COUT(\final_adder.$signal$144 ),
    .SUM(\final_adder.$signal$1161 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$710  (.A(\final_adder.p_new$734 ),
    .B(\final_adder.p_new$718 ),
    .X(\final_adder.p_new$838 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$711  (.A1(\final_adder.p_new$718 ),
    .A2(\final_adder.g_new$735 ),
    .B1(\final_adder.g_new$719 ),
    .X(\final_adder.g_new$839 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$712  (.A(\final_adder.p_new$736 ),
    .B(\final_adder.p_new$720 ),
    .X(\final_adder.p_new$840 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$713  (.A1(\final_adder.p_new$720 ),
    .A2(\final_adder.g_new$737 ),
    .B1(\final_adder.g_new$721 ),
    .X(\final_adder.g_new$841 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$714  (.A(\final_adder.p_new$738 ),
    .B(\final_adder.p_new$722 ),
    .X(\final_adder.p_new$842 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$715  (.A1(\final_adder.p_new$722 ),
    .A2(\final_adder.g_new$739 ),
    .B1(\final_adder.g_new$723 ),
    .X(\final_adder.g_new$843 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$716  (.A(\final_adder.p_new$740 ),
    .B(\final_adder.p_new$724 ),
    .X(\final_adder.p_new$844 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$717  (.A1(\final_adder.p_new$724 ),
    .A2(\final_adder.g_new$741 ),
    .B1(\final_adder.g_new$725 ),
    .X(\final_adder.g_new$845 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$718  (.A(\final_adder.p_new$742 ),
    .B(\final_adder.p_new$726 ),
    .X(\final_adder.p_new$846 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$719  (.A1(\final_adder.p_new$726 ),
    .A2(\final_adder.g_new$743 ),
    .B1(\final_adder.g_new$727 ),
    .X(\final_adder.g_new$847 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$72  (.A(\c$4294 ),
    .B(\s$4297 ),
    .COUT(\final_adder.$signal$146 ),
    .SUM(\final_adder.$signal$1162 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$720  (.A(\final_adder.p_new$744 ),
    .B(\final_adder.p_new$728 ),
    .X(\final_adder.p_new$848 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$721  (.A1(\final_adder.p_new$728 ),
    .A2(\final_adder.g_new$745 ),
    .B1(\final_adder.g_new$729 ),
    .X(\final_adder.g_new$849 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$723  (.A1(\final_adder.p_new$730 ),
    .A2(\final_adder.g_new$747 ),
    .B1(\final_adder.g_new$731 ),
    .X(\final_adder.g_new$851 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$725  (.A1(\final_adder.p_new$732 ),
    .A2(\final_adder.g_new$749 ),
    .B1(\final_adder.g_new$733 ),
    .X(\final_adder.g_new$853 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$727  (.A1(\final_adder.p_new$734 ),
    .A2(\final_adder.g_new$751 ),
    .B1(\final_adder.g_new$735 ),
    .X(\final_adder.g_new$855 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$729  (.A1(\final_adder.p_new$736 ),
    .A2(\final_adder.g_new$753 ),
    .B1(\final_adder.g_new$737 ),
    .X(\final_adder.g_new$857 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$73  (.A(\c$4296 ),
    .B(\s$4299 ),
    .COUT(\final_adder.$signal$148 ),
    .SUM(\final_adder.$signal$1163 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$731  (.A1(\final_adder.p_new$738 ),
    .A2(\final_adder.g_new$631 ),
    .B1(\final_adder.g_new$739 ),
    .X(\final_adder.g_new$859 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$733  (.A1(\final_adder.p_new$740 ),
    .A2(\final_adder.g_new$633 ),
    .B1(\final_adder.g_new$741 ),
    .X(\final_adder.g_new$861 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$735  (.A1(\final_adder.p_new$742 ),
    .A2(\final_adder.g_new$509 ),
    .B1(\final_adder.g_new$743 ),
    .X(\final_adder.g_new$863 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$737  (.A1(\final_adder.p_new$744 ),
    .A2(\final_adder.g_new$383 ),
    .B1(\final_adder.g_new$745 ),
    .X(\final_adder.g_new$865 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$74  (.A(\c$4298 ),
    .B(\s$4301 ),
    .COUT(\final_adder.$signal$150 ),
    .SUM(\final_adder.$signal$1164 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$740  (.A(\final_adder.p_new$788 ),
    .B(\final_adder.p_new$756 ),
    .X(\final_adder.p_new$868 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$741  (.A1(\final_adder.p_new$756 ),
    .A2(\final_adder.g_new$789 ),
    .B1(\final_adder.g_new$757 ),
    .X(\final_adder.g_new$869 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$742  (.A(\final_adder.p_new$790 ),
    .B(\final_adder.p_new$758 ),
    .X(\final_adder.p_new$870 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$743  (.A1(\final_adder.p_new$758 ),
    .A2(\final_adder.g_new$791 ),
    .B1(\final_adder.g_new$759 ),
    .X(\final_adder.g_new$871 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$744  (.A(\final_adder.p_new$792 ),
    .B(\final_adder.p_new$760 ),
    .X(\final_adder.p_new$872 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$745  (.A1(\final_adder.p_new$760 ),
    .A2(\final_adder.g_new$793 ),
    .B1(\final_adder.g_new$761 ),
    .X(\final_adder.g_new$873 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$746  (.A(\final_adder.p_new$794 ),
    .B(\final_adder.p_new$762 ),
    .X(\final_adder.p_new$874 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$747  (.A1(\final_adder.p_new$762 ),
    .A2(\final_adder.g_new$795 ),
    .B1(\final_adder.g_new$763 ),
    .X(\final_adder.g_new$875 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$748  (.A(\final_adder.p_new$796 ),
    .B(\final_adder.p_new$764 ),
    .X(\final_adder.p_new$876 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$749  (.A1(\final_adder.p_new$764 ),
    .A2(\final_adder.g_new$797 ),
    .B1(\final_adder.g_new$765 ),
    .X(\final_adder.g_new$877 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$75  (.A(\c$4300 ),
    .B(\s$4303 ),
    .COUT(\final_adder.$signal$152 ),
    .SUM(\final_adder.$signal$1165 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$750  (.A(\final_adder.p_new$798 ),
    .B(\final_adder.p_new$766 ),
    .X(\final_adder.p_new$878 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$751  (.A1(\final_adder.p_new$766 ),
    .A2(\final_adder.g_new$799 ),
    .B1(\final_adder.g_new$767 ),
    .X(\final_adder.g_new$879 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$752  (.A(\final_adder.p_new$800 ),
    .B(\final_adder.p_new$768 ),
    .X(\final_adder.p_new$880 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$753  (.A1(\final_adder.p_new$768 ),
    .A2(\final_adder.g_new$801 ),
    .B1(\final_adder.g_new$769 ),
    .X(\final_adder.g_new$881 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$754  (.A(\final_adder.p_new$802 ),
    .B(\final_adder.p_new$770 ),
    .X(\final_adder.p_new$882 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$755  (.A1(\final_adder.p_new$770 ),
    .A2(\final_adder.g_new$803 ),
    .B1(\final_adder.g_new$771 ),
    .X(\final_adder.g_new$883 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$756  (.A(\final_adder.p_new$804 ),
    .B(\final_adder.p_new$772 ),
    .X(\final_adder.p_new$884 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$757  (.A1(\final_adder.p_new$772 ),
    .A2(\final_adder.g_new$805 ),
    .B1(\final_adder.g_new$773 ),
    .X(\final_adder.g_new$885 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$758  (.A(\final_adder.p_new$806 ),
    .B(\final_adder.p_new$774 ),
    .X(\final_adder.p_new$886 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$759  (.A1(\final_adder.p_new$774 ),
    .A2(\final_adder.g_new$807 ),
    .B1(\final_adder.g_new$775 ),
    .X(\final_adder.g_new$887 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$76  (.A(\c$4302 ),
    .B(\s$4305 ),
    .COUT(\final_adder.$signal$154 ),
    .SUM(\final_adder.$signal$1166 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$760  (.A(\final_adder.p_new$808 ),
    .B(\final_adder.p_new$776 ),
    .X(\final_adder.p_new$888 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$761  (.A1(\final_adder.p_new$776 ),
    .A2(\final_adder.g_new$809 ),
    .B1(\final_adder.g_new$777 ),
    .X(\final_adder.g_new$889 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$762  (.A(\final_adder.p_new$810 ),
    .B(\final_adder.p_new$778 ),
    .X(\final_adder.p_new$890 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$763  (.A1(\final_adder.p_new$778 ),
    .A2(\final_adder.g_new$811 ),
    .B1(\final_adder.g_new$779 ),
    .X(\final_adder.g_new$891 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$764  (.A(\final_adder.p_new$812 ),
    .B(\final_adder.p_new$780 ),
    .X(\final_adder.p_new$892 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$765  (.A1(\final_adder.p_new$780 ),
    .A2(\final_adder.g_new$813 ),
    .B1(\final_adder.g_new$781 ),
    .X(\final_adder.g_new$893 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$766  (.A(\final_adder.p_new$814 ),
    .B(\final_adder.p_new$782 ),
    .X(\final_adder.p_new$894 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$767  (.A1(\final_adder.p_new$782 ),
    .A2(\final_adder.g_new$815 ),
    .B1(\final_adder.g_new$783 ),
    .X(\final_adder.g_new$895 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$768  (.A(\final_adder.p_new$816 ),
    .B(\final_adder.p_new$784 ),
    .X(\final_adder.p_new$896 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$769  (.A1(\final_adder.p_new$784 ),
    .A2(\final_adder.g_new$817 ),
    .B1(\final_adder.g_new$785 ),
    .X(\final_adder.g_new$897 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$77  (.A(\c$4304 ),
    .B(\s$4307 ),
    .COUT(\final_adder.$signal$156 ),
    .SUM(\final_adder.$signal$1167 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$770  (.A(\final_adder.p_new$818 ),
    .B(\final_adder.p_new$786 ),
    .X(\final_adder.p_new$898 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$771  (.A1(\final_adder.p_new$786 ),
    .A2(\final_adder.g_new$819 ),
    .B1(\final_adder.g_new$787 ),
    .X(\final_adder.g_new$899 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$772  (.A(\final_adder.p_new$820 ),
    .B(\final_adder.p_new$788 ),
    .X(\final_adder.p_new$900 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$773  (.A1(\final_adder.p_new$788 ),
    .A2(\final_adder.g_new$821 ),
    .B1(\final_adder.g_new$789 ),
    .X(\final_adder.g_new$901 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$774  (.A(\final_adder.p_new$822 ),
    .B(\final_adder.p_new$790 ),
    .X(\final_adder.p_new$902 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$775  (.A1(\final_adder.p_new$790 ),
    .A2(\final_adder.g_new$823 ),
    .B1(\final_adder.g_new$791 ),
    .X(\final_adder.g_new$903 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$776  (.A(\final_adder.p_new$824 ),
    .B(\final_adder.p_new$792 ),
    .X(\final_adder.p_new$904 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$777  (.A1(\final_adder.p_new$792 ),
    .A2(\final_adder.g_new$825 ),
    .B1(\final_adder.g_new$793 ),
    .X(\final_adder.g_new$905 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$778  (.A(\final_adder.p_new$826 ),
    .B(\final_adder.p_new$794 ),
    .X(\final_adder.p_new$906 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$779  (.A1(\final_adder.p_new$794 ),
    .A2(\final_adder.g_new$827 ),
    .B1(\final_adder.g_new$795 ),
    .X(\final_adder.g_new$907 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$78  (.A(\c$4306 ),
    .B(\s$4309 ),
    .COUT(\final_adder.$signal$158 ),
    .SUM(\final_adder.$signal$1168 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$780  (.A(\final_adder.p_new$828 ),
    .B(\final_adder.p_new$796 ),
    .X(\final_adder.p_new$908 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$781  (.A1(\final_adder.p_new$796 ),
    .A2(\final_adder.g_new$829 ),
    .B1(\final_adder.g_new$797 ),
    .X(\final_adder.g_new$909 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$782  (.A(\final_adder.p_new$830 ),
    .B(\final_adder.p_new$798 ),
    .X(\final_adder.p_new$910 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$783  (.A1(\final_adder.p_new$798 ),
    .A2(\final_adder.g_new$831 ),
    .B1(\final_adder.g_new$799 ),
    .X(\final_adder.g_new$911 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$784  (.A(\final_adder.p_new$832 ),
    .B(\final_adder.p_new$800 ),
    .X(\final_adder.p_new$912 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$785  (.A1(\final_adder.p_new$800 ),
    .A2(\final_adder.g_new$833 ),
    .B1(\final_adder.g_new$801 ),
    .X(\final_adder.g_new$913 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$786  (.A(\final_adder.p_new$834 ),
    .B(\final_adder.p_new$802 ),
    .X(\final_adder.p_new$914 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$787  (.A1(\final_adder.p_new$802 ),
    .A2(\final_adder.g_new$835 ),
    .B1(\final_adder.g_new$803 ),
    .X(\final_adder.g_new$915 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$788  (.A(\final_adder.p_new$836 ),
    .B(\final_adder.p_new$804 ),
    .X(\final_adder.p_new$916 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$789  (.A1(\final_adder.p_new$804 ),
    .A2(\final_adder.g_new$837 ),
    .B1(\final_adder.g_new$805 ),
    .X(\final_adder.g_new$917 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$79  (.A(\c$4308 ),
    .B(\s$4311 ),
    .COUT(\final_adder.$signal$160 ),
    .SUM(\final_adder.$signal$1169 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$790  (.A(\final_adder.p_new$838 ),
    .B(\final_adder.p_new$806 ),
    .X(\final_adder.p_new$918 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$791  (.A1(\final_adder.p_new$806 ),
    .A2(\final_adder.g_new$839 ),
    .B1(\final_adder.g_new$807 ),
    .X(\final_adder.g_new$919 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$792  (.A(\final_adder.p_new$840 ),
    .B(\final_adder.p_new$808 ),
    .X(\final_adder.p_new$920 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$793  (.A1(\final_adder.p_new$808 ),
    .A2(\final_adder.g_new$841 ),
    .B1(\final_adder.g_new$809 ),
    .X(\final_adder.g_new$921 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$794  (.A(\final_adder.p_new$842 ),
    .B(\final_adder.p_new$810 ),
    .X(\final_adder.p_new$922 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$795  (.A1(\final_adder.p_new$810 ),
    .A2(\final_adder.g_new$843 ),
    .B1(\final_adder.g_new$811 ),
    .X(\final_adder.g_new$923 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$796  (.A(\final_adder.p_new$844 ),
    .B(\final_adder.p_new$812 ),
    .X(\final_adder.p_new$924 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$797  (.A1(\final_adder.p_new$812 ),
    .A2(\final_adder.g_new$845 ),
    .B1(\final_adder.g_new$813 ),
    .X(\final_adder.g_new$925 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$798  (.A(\final_adder.p_new$846 ),
    .B(\final_adder.p_new$814 ),
    .X(\final_adder.p_new$926 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$799  (.A1(\final_adder.p_new$814 ),
    .A2(\final_adder.g_new$847 ),
    .B1(\final_adder.g_new$815 ),
    .X(\final_adder.g_new$927 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$8  (.A(\c$4166 ),
    .B(\s$4169 ),
    .COUT(\final_adder.$signal$18 ),
    .SUM(\final_adder.$signal$1098 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$80  (.A(\c$4310 ),
    .B(\s$4313 ),
    .COUT(\final_adder.$signal$162 ),
    .SUM(\final_adder.$signal$1170 ));
 sky130_fd_sc_hd__and2_1 \final_adder.U$$800  (.A(\final_adder.p_new$848 ),
    .B(\final_adder.p_new$816 ),
    .X(\final_adder.p_new$928 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$801  (.A1(\final_adder.p_new$816 ),
    .A2(\final_adder.g_new$849 ),
    .B1(\final_adder.g_new$817 ),
    .X(\final_adder.g_new$929 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$803  (.A1(\final_adder.p_new$818 ),
    .A2(\final_adder.g_new$851 ),
    .B1(\final_adder.g_new$819 ),
    .X(\final_adder.g_new$931 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$805  (.A1(\final_adder.p_new$820 ),
    .A2(\final_adder.g_new$853 ),
    .B1(\final_adder.g_new$821 ),
    .X(\final_adder.g_new$933 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$807  (.A1(\final_adder.p_new$822 ),
    .A2(\final_adder.g_new$855 ),
    .B1(\final_adder.g_new$823 ),
    .X(\final_adder.g_new$935 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$809  (.A1(\final_adder.p_new$824 ),
    .A2(\final_adder.g_new$857 ),
    .B1(\final_adder.g_new$825 ),
    .X(\final_adder.g_new$937 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$81  (.A(\c$4312 ),
    .B(\s$4315 ),
    .COUT(\final_adder.$signal$164 ),
    .SUM(\final_adder.$signal$1171 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$811  (.A1(\final_adder.p_new$826 ),
    .A2(\final_adder.g_new$859 ),
    .B1(\final_adder.g_new$827 ),
    .X(\final_adder.g_new$939 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$813  (.A1(\final_adder.p_new$828 ),
    .A2(\final_adder.g_new$861 ),
    .B1(\final_adder.g_new$829 ),
    .X(\final_adder.g_new$941 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$815  (.A1(\final_adder.p_new$830 ),
    .A2(\final_adder.g_new$863 ),
    .B1(\final_adder.g_new$831 ),
    .X(\final_adder.g_new$943 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$817  (.A1(\final_adder.p_new$832 ),
    .A2(\final_adder.g_new$865 ),
    .B1(\final_adder.g_new$833 ),
    .X(\final_adder.g_new$945 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$819  (.A1(\final_adder.p_new$834 ),
    .A2(\final_adder.g_new$747 ),
    .B1(\final_adder.g_new$835 ),
    .X(\final_adder.g_new$947 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$82  (.A(\c$4314 ),
    .B(\s$4317 ),
    .COUT(\final_adder.$signal$166 ),
    .SUM(\final_adder.$signal$1172 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$821  (.A1(\final_adder.p_new$836 ),
    .A2(\final_adder.g_new$749 ),
    .B1(\final_adder.g_new$837 ),
    .X(\final_adder.g_new$949 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$823  (.A1(\final_adder.p_new$838 ),
    .A2(\final_adder.g_new$751 ),
    .B1(\final_adder.g_new$839 ),
    .X(\final_adder.g_new$951 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$825  (.A1(\final_adder.p_new$840 ),
    .A2(\final_adder.g_new$753 ),
    .B1(\final_adder.g_new$841 ),
    .X(\final_adder.g_new$953 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$827  (.A1(\final_adder.p_new$842 ),
    .A2(\final_adder.g_new$631 ),
    .B1(\final_adder.g_new$843 ),
    .X(\final_adder.g_new$955 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$829  (.A1(\final_adder.p_new$844 ),
    .A2(\final_adder.g_new$633 ),
    .B1(\final_adder.g_new$845 ),
    .X(\final_adder.g_new$957 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$83  (.A(\c$4316 ),
    .B(\s$4319 ),
    .COUT(\final_adder.$signal$168 ),
    .SUM(\final_adder.$signal$1173 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$831  (.A1(\final_adder.p_new$846 ),
    .A2(\final_adder.g_new$509 ),
    .B1(\final_adder.g_new$847 ),
    .X(\final_adder.g_new$959 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$833  (.A1(\final_adder.p_new$848 ),
    .A2(\final_adder.g_new$383 ),
    .B1(\final_adder.g_new$849 ),
    .X(\final_adder.g_new$961 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$837  (.A1(\final_adder.p_new$868 ),
    .A2(\final_adder.g_new$933 ),
    .B1(\final_adder.g_new$869 ),
    .X(\final_adder.g_new$965 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$839  (.A1(\final_adder.p_new$870 ),
    .A2(\final_adder.g_new$935 ),
    .B1(\final_adder.g_new$871 ),
    .X(\final_adder.g_new$967 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$84  (.A(\c$4318 ),
    .B(\s$4321 ),
    .COUT(\final_adder.$signal$170 ),
    .SUM(\final_adder.$signal$1174 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$841  (.A1(\final_adder.p_new$872 ),
    .A2(\final_adder.g_new$937 ),
    .B1(\final_adder.g_new$873 ),
    .X(\final_adder.g_new$969 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$843  (.A1(\final_adder.p_new$874 ),
    .A2(\final_adder.g_new$939 ),
    .B1(\final_adder.g_new$875 ),
    .X(\final_adder.g_new$971 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$845  (.A1(\final_adder.p_new$876 ),
    .A2(\final_adder.g_new$941 ),
    .B1(\final_adder.g_new$877 ),
    .X(\final_adder.g_new$973 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$847  (.A1(\final_adder.p_new$878 ),
    .A2(\final_adder.g_new$943 ),
    .B1(\final_adder.g_new$879 ),
    .X(\final_adder.g_new$975 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$849  (.A1(\final_adder.p_new$880 ),
    .A2(\final_adder.g_new$945 ),
    .B1(\final_adder.g_new$881 ),
    .X(\final_adder.g_new$977 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$85  (.A(\c$4320 ),
    .B(\s$4323 ),
    .COUT(\final_adder.$signal$172 ),
    .SUM(\final_adder.$signal$1175 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$851  (.A1(\final_adder.p_new$882 ),
    .A2(\final_adder.g_new$947 ),
    .B1(\final_adder.g_new$883 ),
    .X(\final_adder.g_new$979 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$853  (.A1(\final_adder.p_new$884 ),
    .A2(\final_adder.g_new$949 ),
    .B1(\final_adder.g_new$885 ),
    .X(\final_adder.g_new$981 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$855  (.A1(\final_adder.p_new$886 ),
    .A2(\final_adder.g_new$951 ),
    .B1(\final_adder.g_new$887 ),
    .X(\final_adder.g_new$983 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$857  (.A1(\final_adder.p_new$888 ),
    .A2(\final_adder.g_new$953 ),
    .B1(\final_adder.g_new$889 ),
    .X(\final_adder.g_new$985 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$859  (.A1(\final_adder.p_new$890 ),
    .A2(\final_adder.g_new$955 ),
    .B1(\final_adder.g_new$891 ),
    .X(\final_adder.g_new$987 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$86  (.A(\c$4322 ),
    .B(\s$4325 ),
    .COUT(\final_adder.$signal$174 ),
    .SUM(\final_adder.$signal$1176 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$861  (.A1(\final_adder.p_new$892 ),
    .A2(\final_adder.g_new$957 ),
    .B1(\final_adder.g_new$893 ),
    .X(\final_adder.g_new$989 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$863  (.A1(\final_adder.p_new$894 ),
    .A2(\final_adder.g_new$959 ),
    .B1(\final_adder.g_new$895 ),
    .X(\final_adder.g_new$991 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$865  (.A1(\final_adder.p_new$896 ),
    .A2(\final_adder.g_new$961 ),
    .B1(\final_adder.g_new$897 ),
    .X(\final_adder.g_new$993 ));
 sky130_fd_sc_hd__a21o_2 \final_adder.U$$867  (.A1(\final_adder.p_new$898 ),
    .A2(\final_adder.g_new$851 ),
    .B1(\final_adder.g_new$899 ),
    .X(\final_adder.g_new$995 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$869  (.A1(\final_adder.p_new$900 ),
    .A2(\final_adder.g_new$853 ),
    .B1(\final_adder.g_new$901 ),
    .X(\final_adder.g_new$997 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$87  (.A(\c$4324 ),
    .B(\s$4327 ),
    .COUT(\final_adder.$signal$176 ),
    .SUM(\final_adder.$signal$1177 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$871  (.A1(\final_adder.p_new$902 ),
    .A2(\final_adder.g_new$855 ),
    .B1(\final_adder.g_new$903 ),
    .X(\final_adder.g_new$999 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$873  (.A1(\final_adder.p_new$904 ),
    .A2(\final_adder.g_new$857 ),
    .B1(\final_adder.g_new$905 ),
    .X(\final_adder.g_new$1001 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$875  (.A1(\final_adder.p_new$906 ),
    .A2(\final_adder.g_new$859 ),
    .B1(\final_adder.g_new$907 ),
    .X(\final_adder.g_new$1003 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$877  (.A1(\final_adder.p_new$908 ),
    .A2(\final_adder.g_new$861 ),
    .B1(\final_adder.g_new$909 ),
    .X(\final_adder.g_new$1005 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$879  (.A1(\final_adder.p_new$910 ),
    .A2(\final_adder.g_new$863 ),
    .B1(\final_adder.g_new$911 ),
    .X(\final_adder.g_new$1007 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$88  (.A(\c$4326 ),
    .B(\s$4329 ),
    .COUT(\final_adder.$signal$178 ),
    .SUM(\final_adder.$signal$1178 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$881  (.A1(\final_adder.p_new$912 ),
    .A2(\final_adder.g_new$865 ),
    .B1(\final_adder.g_new$913 ),
    .X(\final_adder.g_new$1009 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$883  (.A1(\final_adder.p_new$914 ),
    .A2(\final_adder.g_new$747 ),
    .B1(\final_adder.g_new$915 ),
    .X(\final_adder.g_new$1011 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$885  (.A1(\final_adder.p_new$916 ),
    .A2(\final_adder.g_new$749 ),
    .B1(\final_adder.g_new$917 ),
    .X(\final_adder.g_new$1013 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$887  (.A1(\final_adder.p_new$918 ),
    .A2(\final_adder.g_new$751 ),
    .B1(\final_adder.g_new$919 ),
    .X(\final_adder.g_new$1015 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$889  (.A1(\final_adder.p_new$920 ),
    .A2(\final_adder.g_new$753 ),
    .B1(\final_adder.g_new$921 ),
    .X(\final_adder.g_new$1017 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$89  (.A(\c$4328 ),
    .B(\s$4331 ),
    .COUT(\final_adder.$signal$180 ),
    .SUM(\final_adder.$signal$1179 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$891  (.A1(\final_adder.p_new$922 ),
    .A2(\final_adder.g_new$631 ),
    .B1(\final_adder.g_new$923 ),
    .X(\final_adder.g_new$1019 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$893  (.A1(\final_adder.p_new$924 ),
    .A2(\final_adder.g_new$633 ),
    .B1(\final_adder.g_new$925 ),
    .X(\final_adder.g_new$1021 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$895  (.A1(\final_adder.p_new$926 ),
    .A2(\final_adder.g_new$509 ),
    .B1(\final_adder.g_new$927 ),
    .X(\final_adder.g_new$1023 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$897  (.A1(\final_adder.p_new$928 ),
    .A2(\final_adder.g_new$383 ),
    .B1(\final_adder.g_new$929 ),
    .X(\final_adder.g_new$1025 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$898  (.A1(\final_adder.$signal$1216 ),
    .A2(\final_adder.g_new$965 ),
    .B1(\final_adder.$signal$254 ),
    .X(\final_adder.g_new$1026 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$899  (.A1(\final_adder.$signal$1214 ),
    .A2(\final_adder.g_new$967 ),
    .B1(\final_adder.$signal$250 ),
    .X(\final_adder.g_new$1027 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$9  (.A(\c$4168 ),
    .B(\s$4171 ),
    .COUT(\final_adder.$signal$20 ),
    .SUM(\final_adder.$signal$1099 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$90  (.A(\c$4330 ),
    .B(\s$4333 ),
    .COUT(\final_adder.$signal$182 ),
    .SUM(\final_adder.$signal$1180 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$900  (.A1(\final_adder.$signal$1212 ),
    .A2(\final_adder.g_new$969 ),
    .B1(\final_adder.$signal$246 ),
    .X(\final_adder.g_new$1028 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$901  (.A1(\final_adder.$signal$1210 ),
    .A2(\final_adder.g_new$971 ),
    .B1(\final_adder.$signal$242 ),
    .X(\final_adder.g_new$1029 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$902  (.A1(\final_adder.$signal$1208 ),
    .A2(\final_adder.g_new$973 ),
    .B1(\final_adder.$signal$238 ),
    .X(\final_adder.g_new$1030 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$903  (.A1(\final_adder.$signal$1206 ),
    .A2(\final_adder.g_new$975 ),
    .B1(\final_adder.$signal$234 ),
    .X(\final_adder.g_new$1031 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$904  (.A1(\final_adder.$signal$1204 ),
    .A2(\final_adder.g_new$977 ),
    .B1(\final_adder.$signal$230 ),
    .X(\final_adder.g_new$1032 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$905  (.A1(\final_adder.$signal$1202 ),
    .A2(\final_adder.g_new$979 ),
    .B1(\final_adder.$signal$226 ),
    .X(\final_adder.g_new$1033 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$906  (.A1(\final_adder.$signal$1200 ),
    .A2(\final_adder.g_new$981 ),
    .B1(\final_adder.$signal$222 ),
    .X(\final_adder.g_new$1034 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$907  (.A1(\final_adder.$signal$1198 ),
    .A2(\final_adder.g_new$983 ),
    .B1(\final_adder.$signal$218 ),
    .X(\final_adder.g_new$1035 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$908  (.A1(\final_adder.$signal$1196 ),
    .A2(\final_adder.g_new$985 ),
    .B1(\final_adder.$signal$214 ),
    .X(\final_adder.g_new$1036 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$909  (.A1(\final_adder.$signal$1194 ),
    .A2(\final_adder.g_new$987 ),
    .B1(\final_adder.$signal$210 ),
    .X(\final_adder.g_new$1037 ));
 sky130_fd_sc_hd__ha_2 \final_adder.U$$91  (.A(\c$4332 ),
    .B(\s$4335 ),
    .COUT(\final_adder.$signal$184 ),
    .SUM(\final_adder.$signal$1181 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$910  (.A1(\final_adder.$signal$1192 ),
    .A2(\final_adder.g_new$989 ),
    .B1(\final_adder.$signal$206 ),
    .X(\final_adder.g_new$1038 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$911  (.A1(\final_adder.$signal$1190 ),
    .A2(\final_adder.g_new$991 ),
    .B1(\final_adder.$signal$202 ),
    .X(\final_adder.g_new$1039 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$912  (.A1(\final_adder.$signal$1188 ),
    .A2(\final_adder.g_new$993 ),
    .B1(\final_adder.$signal$198 ),
    .X(\final_adder.g_new$1040 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$913  (.A1(\final_adder.$signal$1186 ),
    .A2(\final_adder.g_new$995 ),
    .B1(\final_adder.$signal$194 ),
    .X(\final_adder.g_new$1041 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$914  (.A1(\final_adder.$signal$1184 ),
    .A2(\final_adder.g_new$997 ),
    .B1(\final_adder.$signal$190 ),
    .X(\final_adder.g_new$1042 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$915  (.A1(\final_adder.$signal$1182 ),
    .A2(\final_adder.g_new$999 ),
    .B1(\final_adder.$signal$186 ),
    .X(\final_adder.g_new$1043 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$916  (.A1(\final_adder.$signal$1180 ),
    .A2(\final_adder.g_new$1001 ),
    .B1(\final_adder.$signal$182 ),
    .X(\final_adder.g_new$1044 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$917  (.A1(\final_adder.$signal$1178 ),
    .A2(\final_adder.g_new$1003 ),
    .B1(\final_adder.$signal$178 ),
    .X(\final_adder.g_new$1045 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$918  (.A1(\final_adder.$signal$1176 ),
    .A2(\final_adder.g_new$1005 ),
    .B1(\final_adder.$signal$174 ),
    .X(\final_adder.g_new$1046 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$919  (.A1(\final_adder.$signal$1174 ),
    .A2(\final_adder.g_new$1007 ),
    .B1(\final_adder.$signal$170 ),
    .X(\final_adder.g_new$1047 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$92  (.A(\c$4334 ),
    .B(\s$4337 ),
    .COUT(\final_adder.$signal$186 ),
    .SUM(\final_adder.$signal$1182 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$920  (.A1(\final_adder.$signal$1172 ),
    .A2(\final_adder.g_new$1009 ),
    .B1(\final_adder.$signal$166 ),
    .X(\final_adder.g_new$1048 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$921  (.A1(\final_adder.$signal$1170 ),
    .A2(\final_adder.g_new$1011 ),
    .B1(\final_adder.$signal$162 ),
    .X(\final_adder.g_new$1049 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$922  (.A1(\final_adder.$signal$1168 ),
    .A2(\final_adder.g_new$1013 ),
    .B1(\final_adder.$signal$158 ),
    .X(\final_adder.g_new$1050 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$923  (.A1(\final_adder.$signal$1166 ),
    .A2(\final_adder.g_new$1015 ),
    .B1(\final_adder.$signal$154 ),
    .X(\final_adder.g_new$1051 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$924  (.A1(\final_adder.$signal$1164 ),
    .A2(\final_adder.g_new$1017 ),
    .B1(\final_adder.$signal$150 ),
    .X(\final_adder.g_new$1052 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$925  (.A1(\final_adder.$signal$1162 ),
    .A2(\final_adder.g_new$1019 ),
    .B1(\final_adder.$signal$146 ),
    .X(\final_adder.g_new$1053 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$926  (.A1(\final_adder.$signal$1160 ),
    .A2(\final_adder.g_new$1021 ),
    .B1(\final_adder.$signal$142 ),
    .X(\final_adder.g_new$1054 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$927  (.A1(\final_adder.$signal$1158 ),
    .A2(\final_adder.g_new$1023 ),
    .B1(\final_adder.$signal$138 ),
    .X(\final_adder.g_new$1055 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$928  (.A1(\final_adder.$signal$1156 ),
    .A2(\final_adder.g_new$1025 ),
    .B1(\final_adder.$signal$134 ),
    .X(\final_adder.g_new$1056 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$929  (.A1(\final_adder.$signal$1154 ),
    .A2(\final_adder.g_new$931 ),
    .B1(\final_adder.$signal$130 ),
    .X(\final_adder.g_new$1057 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$93  (.A(\c$4336 ),
    .B(\s$4339 ),
    .COUT(\final_adder.$signal$188 ),
    .SUM(\final_adder.$signal$1183 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$930  (.A1(\final_adder.$signal$1152 ),
    .A2(\final_adder.g_new$933 ),
    .B1(\final_adder.$signal$126 ),
    .X(\final_adder.g_new$1058 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$931  (.A1(\final_adder.$signal$1150 ),
    .A2(\final_adder.g_new$935 ),
    .B1(\final_adder.$signal$122 ),
    .X(\final_adder.g_new$1059 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$932  (.A1(\final_adder.$signal$1148 ),
    .A2(\final_adder.g_new$937 ),
    .B1(\final_adder.$signal$118 ),
    .X(\final_adder.g_new$1060 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$933  (.A1(\final_adder.$signal$1146 ),
    .A2(\final_adder.g_new$939 ),
    .B1(\final_adder.$signal$114 ),
    .X(\final_adder.g_new$1061 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$934  (.A1(\final_adder.$signal$111 ),
    .A2(\final_adder.g_new$941 ),
    .B1(\final_adder.$signal$110 ),
    .X(\final_adder.g_new$1062 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$935  (.A1(\final_adder.$signal$107 ),
    .A2(\final_adder.g_new$943 ),
    .B1(\final_adder.$signal$106 ),
    .X(\final_adder.g_new$1063 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$936  (.A1(\final_adder.$signal$103 ),
    .A2(\final_adder.g_new$945 ),
    .B1(\final_adder.$signal$102 ),
    .X(\final_adder.g_new$1064 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$937  (.A1(\final_adder.$signal$1138 ),
    .A2(\final_adder.g_new$947 ),
    .B1(\final_adder.$signal$98 ),
    .X(\final_adder.g_new$1065 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$938  (.A1(\final_adder.$signal$1136 ),
    .A2(\final_adder.g_new$949 ),
    .B1(\final_adder.$signal$94 ),
    .X(\final_adder.g_new$1066 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$939  (.A1(\final_adder.$signal$1134 ),
    .A2(\final_adder.g_new$951 ),
    .B1(\final_adder.$signal$90 ),
    .X(\final_adder.g_new$1067 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$94  (.A(\c$4338 ),
    .B(\s$4341 ),
    .COUT(\final_adder.$signal$190 ),
    .SUM(\final_adder.$signal$1184 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$940  (.A1(\final_adder.$signal$1132 ),
    .A2(\final_adder.g_new$953 ),
    .B1(\final_adder.$signal$86 ),
    .X(\final_adder.g_new$1068 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$941  (.A1(\final_adder.$signal$1130 ),
    .A2(\final_adder.g_new$955 ),
    .B1(\final_adder.$signal$82 ),
    .X(\final_adder.g_new$1069 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$942  (.A1(\final_adder.$signal$1128 ),
    .A2(\final_adder.g_new$957 ),
    .B1(\final_adder.$signal$78 ),
    .X(\final_adder.g_new$1070 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$943  (.A1(\final_adder.$signal$1126 ),
    .A2(\final_adder.g_new$959 ),
    .B1(\final_adder.$signal$74 ),
    .X(\final_adder.g_new$1071 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$944  (.A1(\final_adder.$signal$1124 ),
    .A2(\final_adder.g_new$961 ),
    .B1(\final_adder.$signal$70 ),
    .X(\final_adder.g_new$1072 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$945  (.A1(\final_adder.$signal$1122 ),
    .A2(\final_adder.g_new$851 ),
    .B1(\final_adder.$signal$66 ),
    .X(\final_adder.g_new$1073 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$946  (.A1(\final_adder.$signal$1120 ),
    .A2(\final_adder.g_new$853 ),
    .B1(\final_adder.$signal$62 ),
    .X(\final_adder.g_new$1074 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$947  (.A1(\final_adder.$signal$1118 ),
    .A2(\final_adder.g_new$855 ),
    .B1(\final_adder.$signal$58 ),
    .X(\final_adder.g_new$1075 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$948  (.A1(\final_adder.$signal$1116 ),
    .A2(\final_adder.g_new$857 ),
    .B1(\final_adder.$signal$54 ),
    .X(\final_adder.g_new$1076 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$949  (.A1(\final_adder.$signal$1114 ),
    .A2(\final_adder.g_new$859 ),
    .B1(\final_adder.$signal$50 ),
    .X(\final_adder.g_new$1077 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$95  (.A(\c$4340 ),
    .B(\s$4343 ),
    .COUT(\final_adder.$signal$192 ),
    .SUM(\final_adder.$signal$1185 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$950  (.A1(\final_adder.$signal$1112 ),
    .A2(\final_adder.g_new$861 ),
    .B1(\final_adder.$signal$46 ),
    .X(\final_adder.g_new$1078 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$951  (.A1(\final_adder.$signal$1110 ),
    .A2(\final_adder.g_new$863 ),
    .B1(\final_adder.$signal$42 ),
    .X(\final_adder.g_new$1079 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$952  (.A1(\final_adder.$signal$1108 ),
    .A2(\final_adder.g_new$865 ),
    .B1(\final_adder.$signal$38 ),
    .X(\final_adder.g_new$1080 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$953  (.A1(\final_adder.$signal$1106 ),
    .A2(\final_adder.g_new$747 ),
    .B1(\final_adder.$signal$34 ),
    .X(\final_adder.g_new$1081 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$954  (.A1(\final_adder.$signal$1104 ),
    .A2(\final_adder.g_new$749 ),
    .B1(\final_adder.$signal$30 ),
    .X(\final_adder.g_new$1082 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$955  (.A1(\final_adder.$signal$1102 ),
    .A2(\final_adder.g_new$751 ),
    .B1(\final_adder.$signal$26 ),
    .X(\final_adder.g_new$1083 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$956  (.A1(\final_adder.$signal$1100 ),
    .A2(\final_adder.g_new$753 ),
    .B1(\final_adder.$signal$22 ),
    .X(\final_adder.g_new$1084 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$957  (.A1(\final_adder.$signal$1098 ),
    .A2(\final_adder.g_new$631 ),
    .B1(\final_adder.$signal$18 ),
    .X(\final_adder.g_new$1085 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$958  (.A1(\final_adder.$signal$1096 ),
    .A2(\final_adder.g_new$633 ),
    .B1(\final_adder.$signal$14 ),
    .X(\final_adder.g_new$1086 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$959  (.A1(\final_adder.$signal$1094 ),
    .A2(\final_adder.g_new$509 ),
    .B1(\final_adder.$signal$10 ),
    .X(\final_adder.g_new$1087 ));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$96  (.A(\c$4342 ),
    .B(\s$4345 ),
    .COUT(\final_adder.$signal$194 ),
    .SUM(\final_adder.$signal$1186 ));
 sky130_fd_sc_hd__a21o_1 \final_adder.U$$960  (.A1(\final_adder.$signal$1092 ),
    .A2(\final_adder.g_new$383 ),
    .B1(\final_adder.$signal$6 ),
    .X(\final_adder.g_new$1088 ));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$961  (.A(\final_adder.$signal$1 ),
    .B(net1890),
    .X(net257));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$962  (.A(\final_adder.$signal$1091 ),
    .B(\final_adder.$signal ),
    .X(net296));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$963  (.A(\final_adder.$signal$1092 ),
    .B(\final_adder.g_new$383 ),
    .X(net307));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$964  (.A(\final_adder.$signal$1093 ),
    .B(\final_adder.g_new$1088 ),
    .X(net318));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$965  (.A(\final_adder.$signal$1094 ),
    .B(\final_adder.g_new$509 ),
    .X(net329));
 sky130_fd_sc_hd__xor2_1 \final_adder.U$$966  (.A(\final_adder.$signal$1095 ),
    .B(\final_adder.g_new$1087 ),
    .X(net340));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$967  (.A(\final_adder.$signal$1096 ),
    .B(\final_adder.g_new$633 ),
    .X(net351));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$968  (.A(\final_adder.$signal$1097 ),
    .B(\final_adder.g_new$1086 ),
    .X(net362));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$969  (.A(\final_adder.$signal$1098 ),
    .B(\final_adder.g_new$631 ),
    .X(net373));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$97  (.A(\c$4344 ),
    .B(\s$4347 ),
    .COUT(\final_adder.$signal$196 ),
    .SUM(\final_adder.$signal$1187 ));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$970  (.A(\final_adder.$signal$1099 ),
    .B(\final_adder.g_new$1085 ),
    .X(net384));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$971  (.A(\final_adder.$signal$1100 ),
    .B(\final_adder.g_new$753 ),
    .X(net268));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$972  (.A(\final_adder.$signal$1101 ),
    .B(\final_adder.g_new$1084 ),
    .X(net279));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$973  (.A(\final_adder.$signal$1102 ),
    .B(\final_adder.g_new$751 ),
    .X(net288));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$974  (.A(\final_adder.$signal$1103 ),
    .B(\final_adder.g_new$1083 ),
    .X(net289));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$975  (.A(\final_adder.$signal$1104 ),
    .B(\final_adder.g_new$749 ),
    .X(net290));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$976  (.A(\final_adder.$signal$1105 ),
    .B(\final_adder.g_new$1082 ),
    .X(net291));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$977  (.A(\final_adder.$signal$1106 ),
    .B(\final_adder.g_new$747 ),
    .X(net292));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$978  (.A(\final_adder.$signal$1107 ),
    .B(\final_adder.g_new$1081 ),
    .X(net293));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$979  (.A(\final_adder.$signal$1108 ),
    .B(\final_adder.g_new$865 ),
    .X(net294));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$98  (.A(\c$4346 ),
    .B(\s$4349 ),
    .COUT(\final_adder.$signal$198 ),
    .SUM(\final_adder.$signal$1188 ));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$980  (.A(\final_adder.$signal$1109 ),
    .B(\final_adder.g_new$1080 ),
    .X(net295));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$981  (.A(\final_adder.$signal$1110 ),
    .B(\final_adder.g_new$863 ),
    .X(net297));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$982  (.A(\final_adder.$signal$1111 ),
    .B(\final_adder.g_new$1079 ),
    .X(net298));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$983  (.A(\final_adder.$signal$1112 ),
    .B(\final_adder.g_new$861 ),
    .X(net299));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$984  (.A(\final_adder.$signal$1113 ),
    .B(\final_adder.g_new$1078 ),
    .X(net300));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$985  (.A(\final_adder.$signal$1114 ),
    .B(\final_adder.g_new$859 ),
    .X(net301));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$986  (.A(\final_adder.$signal$1115 ),
    .B(\final_adder.g_new$1077 ),
    .X(net302));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$987  (.A(\final_adder.$signal$1116 ),
    .B(\final_adder.g_new$857 ),
    .X(net303));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$988  (.A(\final_adder.$signal$1117 ),
    .B(\final_adder.g_new$1076 ),
    .X(net304));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$989  (.A(\final_adder.$signal$1118 ),
    .B(\final_adder.g_new$855 ),
    .X(net305));
 sky130_fd_sc_hd__ha_1 \final_adder.U$$99  (.A(\c$4348 ),
    .B(\s$4351 ),
    .COUT(\final_adder.$signal$200 ),
    .SUM(\final_adder.$signal$1189 ));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$990  (.A(\final_adder.$signal$1119 ),
    .B(\final_adder.g_new$1075 ),
    .X(net306));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$991  (.A(\final_adder.$signal$1120 ),
    .B(\final_adder.g_new$853 ),
    .X(net308));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$992  (.A(\final_adder.$signal$1121 ),
    .B(\final_adder.g_new$1074 ),
    .X(net309));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$993  (.A(\final_adder.$signal$1122 ),
    .B(\final_adder.g_new$851 ),
    .X(net310));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$994  (.A(\final_adder.$signal$1123 ),
    .B(\final_adder.g_new$1073 ),
    .X(net311));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$995  (.A(\final_adder.$signal$1124 ),
    .B(\final_adder.g_new$961 ),
    .X(net312));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$996  (.A(\final_adder.$signal$1125 ),
    .B(\final_adder.g_new$1072 ),
    .X(net313));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$997  (.A(\final_adder.$signal$1126 ),
    .B(\final_adder.g_new$959 ),
    .X(net314));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$998  (.A(\final_adder.$signal$1127 ),
    .B(\final_adder.g_new$1071 ),
    .X(net315));
 sky130_fd_sc_hd__xor2_2 \final_adder.U$$999  (.A(\final_adder.$signal$1128 ),
    .B(\final_adder.g_new$957 ),
    .X(net316));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(a[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_6 input3 (.A(a[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(a[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(a[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(a[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_8 input7 (.A(a[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(a[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(a[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input10 (.A(a[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(a[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(a[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(a[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(a[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(a[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_8 input16 (.A(a[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(a[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_6 input18 (.A(a[25]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(a[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_6 input20 (.A(a[27]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(a[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(a[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_4 input23 (.A(a[2]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(a[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(a[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 input26 (.A(a[32]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(a[33]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(a[34]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(a[35]),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(a[36]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(a[37]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(a[38]),
    .X(net32));
 sky130_fd_sc_hd__buf_6 input33 (.A(a[39]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(a[3]),
    .X(net34));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(a[40]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(a[41]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 input37 (.A(a[42]),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(a[43]),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(a[44]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(a[45]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(a[46]),
    .X(net41));
 sky130_fd_sc_hd__buf_4 input42 (.A(a[47]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(a[48]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(a[49]),
    .X(net44));
 sky130_fd_sc_hd__buf_4 input45 (.A(a[4]),
    .X(net45));
 sky130_fd_sc_hd__buf_2 input46 (.A(a[50]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(a[51]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(a[52]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(a[53]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(a[54]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(a[55]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(a[56]),
    .X(net52));
 sky130_fd_sc_hd__dlymetal6s2s_1 input53 (.A(a[57]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(a[58]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 input55 (.A(a[59]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(a[5]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(a[60]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 input58 (.A(a[61]),
    .X(net58));
 sky130_fd_sc_hd__dlymetal6s2s_1 input59 (.A(a[62]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(a[63]),
    .X(net60));
 sky130_fd_sc_hd__buf_2 input61 (.A(a[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(a[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(a[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_6 input64 (.A(a[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_2 input65 (.A(b[0]),
    .X(net65));
 sky130_fd_sc_hd__buf_6 input66 (.A(b[10]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 input67 (.A(b[11]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(b[12]),
    .X(net68));
 sky130_fd_sc_hd__buf_4 input69 (.A(b[13]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input70 (.A(b[14]),
    .X(net70));
 sky130_fd_sc_hd__buf_6 input71 (.A(b[15]),
    .X(net71));
 sky130_fd_sc_hd__buf_8 input72 (.A(b[16]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 input73 (.A(b[17]),
    .X(net73));
 sky130_fd_sc_hd__buf_8 input74 (.A(b[18]),
    .X(net74));
 sky130_fd_sc_hd__buf_4 input75 (.A(b[19]),
    .X(net75));
 sky130_fd_sc_hd__buf_6 input76 (.A(b[1]),
    .X(net76));
 sky130_fd_sc_hd__buf_6 input77 (.A(b[20]),
    .X(net77));
 sky130_fd_sc_hd__buf_4 input78 (.A(b[21]),
    .X(net78));
 sky130_fd_sc_hd__buf_4 input79 (.A(b[22]),
    .X(net79));
 sky130_fd_sc_hd__buf_4 input80 (.A(b[23]),
    .X(net80));
 sky130_fd_sc_hd__buf_6 input81 (.A(b[24]),
    .X(net81));
 sky130_fd_sc_hd__dlymetal6s2s_1 input82 (.A(b[25]),
    .X(net82));
 sky130_fd_sc_hd__buf_6 input83 (.A(b[26]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 input84 (.A(b[27]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(b[28]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(b[29]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 input87 (.A(b[2]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 input88 (.A(b[30]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(b[31]),
    .X(net89));
 sky130_fd_sc_hd__dlymetal6s2s_1 input90 (.A(b[32]),
    .X(net90));
 sky130_fd_sc_hd__buf_6 input91 (.A(b[33]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_4 input92 (.A(b[34]),
    .X(net92));
 sky130_fd_sc_hd__dlymetal6s2s_1 input93 (.A(b[35]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_4 input94 (.A(b[36]),
    .X(net94));
 sky130_fd_sc_hd__buf_2 input95 (.A(b[37]),
    .X(net95));
 sky130_fd_sc_hd__buf_4 input96 (.A(b[38]),
    .X(net96));
 sky130_fd_sc_hd__dlymetal6s2s_1 input97 (.A(b[39]),
    .X(net97));
 sky130_fd_sc_hd__buf_4 input98 (.A(b[3]),
    .X(net98));
 sky130_fd_sc_hd__dlymetal6s2s_1 input99 (.A(b[40]),
    .X(net99));
 sky130_fd_sc_hd__dlymetal6s2s_1 input100 (.A(b[41]),
    .X(net100));
 sky130_fd_sc_hd__buf_4 input101 (.A(b[42]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_4 input102 (.A(b[43]),
    .X(net102));
 sky130_fd_sc_hd__buf_2 input103 (.A(b[44]),
    .X(net103));
 sky130_fd_sc_hd__buf_6 input104 (.A(b[45]),
    .X(net104));
 sky130_fd_sc_hd__buf_6 input105 (.A(b[46]),
    .X(net105));
 sky130_fd_sc_hd__buf_6 input106 (.A(b[47]),
    .X(net106));
 sky130_fd_sc_hd__buf_6 input107 (.A(b[48]),
    .X(net107));
 sky130_fd_sc_hd__buf_4 input108 (.A(b[49]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 input109 (.A(b[4]),
    .X(net109));
 sky130_fd_sc_hd__buf_6 input110 (.A(b[50]),
    .X(net110));
 sky130_fd_sc_hd__buf_6 input111 (.A(b[51]),
    .X(net111));
 sky130_fd_sc_hd__buf_4 input112 (.A(b[52]),
    .X(net112));
 sky130_fd_sc_hd__buf_2 input113 (.A(b[53]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(b[54]),
    .X(net114));
 sky130_fd_sc_hd__buf_2 input115 (.A(b[55]),
    .X(net115));
 sky130_fd_sc_hd__buf_2 input116 (.A(b[56]),
    .X(net116));
 sky130_fd_sc_hd__buf_2 input117 (.A(b[57]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(b[58]),
    .X(net118));
 sky130_fd_sc_hd__buf_2 input119 (.A(b[59]),
    .X(net119));
 sky130_fd_sc_hd__buf_2 input120 (.A(b[5]),
    .X(net120));
 sky130_fd_sc_hd__dlymetal6s2s_1 input121 (.A(b[60]),
    .X(net121));
 sky130_fd_sc_hd__buf_6 input122 (.A(b[61]),
    .X(net122));
 sky130_fd_sc_hd__buf_4 input123 (.A(b[62]),
    .X(net123));
 sky130_fd_sc_hd__buf_4 input124 (.A(b[63]),
    .X(net124));
 sky130_fd_sc_hd__buf_4 input125 (.A(b[6]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 input126 (.A(b[7]),
    .X(net126));
 sky130_fd_sc_hd__buf_6 input127 (.A(b[8]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 input128 (.A(b[9]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(c[0]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(c[100]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(c[101]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(c[102]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(c[103]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(c[104]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(c[105]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(c[106]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(c[107]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(c[108]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(c[109]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(c[10]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(c[110]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 input142 (.A(c[111]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(c[112]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(c[113]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 input145 (.A(c[114]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 input146 (.A(c[115]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 input147 (.A(c[116]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(c[117]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(c[118]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 input150 (.A(c[119]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(c[11]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(c[120]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 input153 (.A(c[121]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(c[122]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 input155 (.A(c[123]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 input156 (.A(c[124]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 input157 (.A(c[125]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 input158 (.A(c[126]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 input159 (.A(c[127]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 input160 (.A(c[12]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(c[13]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 input162 (.A(c[14]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 input163 (.A(c[15]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(c[16]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 input165 (.A(c[17]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(c[18]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(c[19]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 input168 (.A(c[1]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 input169 (.A(c[20]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(c[21]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 input171 (.A(c[22]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 input172 (.A(c[23]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 input173 (.A(c[24]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 input174 (.A(c[25]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(c[26]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(c[27]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(c[28]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(c[29]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(c[2]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(c[30]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 input181 (.A(c[31]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 input182 (.A(c[32]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(c[33]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(c[34]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(c[35]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(c[36]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(c[37]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(c[38]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 input189 (.A(c[39]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 input190 (.A(c[3]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(c[40]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(c[41]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 input193 (.A(c[42]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(c[43]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 input195 (.A(c[44]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 input196 (.A(c[45]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 input197 (.A(c[46]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 input198 (.A(c[47]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 input199 (.A(c[48]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 input200 (.A(c[49]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 input201 (.A(c[4]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 input202 (.A(c[50]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 input203 (.A(c[51]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 input204 (.A(c[52]),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 input205 (.A(c[53]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 input206 (.A(c[54]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 input207 (.A(c[55]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 input208 (.A(c[56]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 input209 (.A(c[57]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_1 input210 (.A(c[58]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_1 input211 (.A(c[59]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 input212 (.A(c[5]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 input213 (.A(c[60]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 input214 (.A(c[61]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 input215 (.A(c[62]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_1 input216 (.A(c[63]),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_1 input217 (.A(c[64]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_1 input218 (.A(c[65]),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_1 input219 (.A(c[66]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_1 input220 (.A(c[67]),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_1 input221 (.A(c[68]),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_1 input222 (.A(c[69]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_1 input223 (.A(c[6]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_1 input224 (.A(c[70]),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_1 input225 (.A(c[71]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 input226 (.A(c[72]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 input227 (.A(c[73]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 input228 (.A(c[74]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_1 input229 (.A(c[75]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 input230 (.A(c[76]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_1 input231 (.A(c[77]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_1 input232 (.A(c[78]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 input233 (.A(c[79]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 input234 (.A(c[7]),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 input235 (.A(c[80]),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 input236 (.A(c[81]),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_1 input237 (.A(c[82]),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 input238 (.A(c[83]),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 input239 (.A(c[84]),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 input240 (.A(c[85]),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 input241 (.A(c[86]),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_1 input242 (.A(c[87]),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 input243 (.A(c[88]),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 input244 (.A(c[89]),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_1 input245 (.A(c[8]),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_1 input246 (.A(c[90]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_1 input247 (.A(c[91]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_1 input248 (.A(c[92]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 input249 (.A(c[93]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 input250 (.A(c[94]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 input251 (.A(c[95]),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 input252 (.A(c[96]),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_1 input253 (.A(c[97]),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 input254 (.A(c[98]),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_1 input255 (.A(c[99]),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_1 input256 (.A(c[9]),
    .X(net256));
 sky130_fd_sc_hd__buf_2 output257 (.A(net257),
    .X(o[0]));
 sky130_fd_sc_hd__buf_2 output258 (.A(net258),
    .X(o[100]));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .X(o[101]));
 sky130_fd_sc_hd__buf_2 output260 (.A(net260),
    .X(o[102]));
 sky130_fd_sc_hd__buf_2 output261 (.A(net261),
    .X(o[103]));
 sky130_fd_sc_hd__buf_2 output262 (.A(net262),
    .X(o[104]));
 sky130_fd_sc_hd__buf_2 output263 (.A(net263),
    .X(o[105]));
 sky130_fd_sc_hd__buf_2 output264 (.A(net264),
    .X(o[106]));
 sky130_fd_sc_hd__buf_2 output265 (.A(net265),
    .X(o[107]));
 sky130_fd_sc_hd__buf_2 output266 (.A(net266),
    .X(o[108]));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .X(o[109]));
 sky130_fd_sc_hd__buf_2 output268 (.A(net268),
    .X(o[10]));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .X(o[110]));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .X(o[111]));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .X(o[112]));
 sky130_fd_sc_hd__buf_2 output272 (.A(net272),
    .X(o[113]));
 sky130_fd_sc_hd__buf_2 output273 (.A(net273),
    .X(o[114]));
 sky130_fd_sc_hd__buf_2 output274 (.A(net274),
    .X(o[115]));
 sky130_fd_sc_hd__buf_2 output275 (.A(net275),
    .X(o[116]));
 sky130_fd_sc_hd__buf_2 output276 (.A(net276),
    .X(o[117]));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .X(o[118]));
 sky130_fd_sc_hd__buf_2 output278 (.A(net278),
    .X(o[119]));
 sky130_fd_sc_hd__buf_2 output279 (.A(net279),
    .X(o[11]));
 sky130_fd_sc_hd__buf_2 output280 (.A(net280),
    .X(o[120]));
 sky130_fd_sc_hd__buf_2 output281 (.A(net281),
    .X(o[121]));
 sky130_fd_sc_hd__buf_2 output282 (.A(net282),
    .X(o[122]));
 sky130_fd_sc_hd__buf_2 output283 (.A(net283),
    .X(o[123]));
 sky130_fd_sc_hd__buf_2 output284 (.A(net284),
    .X(o[124]));
 sky130_fd_sc_hd__buf_2 output285 (.A(net285),
    .X(o[125]));
 sky130_fd_sc_hd__buf_2 output286 (.A(net286),
    .X(o[126]));
 sky130_fd_sc_hd__buf_2 output287 (.A(net287),
    .X(o[127]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(o[12]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(o[13]));
 sky130_fd_sc_hd__buf_2 output290 (.A(net290),
    .X(o[14]));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .X(o[15]));
 sky130_fd_sc_hd__buf_2 output292 (.A(net292),
    .X(o[16]));
 sky130_fd_sc_hd__buf_2 output293 (.A(net293),
    .X(o[17]));
 sky130_fd_sc_hd__buf_2 output294 (.A(net294),
    .X(o[18]));
 sky130_fd_sc_hd__buf_2 output295 (.A(net295),
    .X(o[19]));
 sky130_fd_sc_hd__buf_2 output296 (.A(net296),
    .X(o[1]));
 sky130_fd_sc_hd__buf_2 output297 (.A(net297),
    .X(o[20]));
 sky130_fd_sc_hd__buf_2 output298 (.A(net298),
    .X(o[21]));
 sky130_fd_sc_hd__buf_2 output299 (.A(net299),
    .X(o[22]));
 sky130_fd_sc_hd__buf_2 output300 (.A(net300),
    .X(o[23]));
 sky130_fd_sc_hd__buf_2 output301 (.A(net301),
    .X(o[24]));
 sky130_fd_sc_hd__buf_2 output302 (.A(net302),
    .X(o[25]));
 sky130_fd_sc_hd__buf_2 output303 (.A(net303),
    .X(o[26]));
 sky130_fd_sc_hd__buf_2 output304 (.A(net304),
    .X(o[27]));
 sky130_fd_sc_hd__buf_2 output305 (.A(net305),
    .X(o[28]));
 sky130_fd_sc_hd__buf_2 output306 (.A(net306),
    .X(o[29]));
 sky130_fd_sc_hd__buf_2 output307 (.A(net307),
    .X(o[2]));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .X(o[30]));
 sky130_fd_sc_hd__buf_2 output309 (.A(net309),
    .X(o[31]));
 sky130_fd_sc_hd__buf_2 output310 (.A(net310),
    .X(o[32]));
 sky130_fd_sc_hd__buf_2 output311 (.A(net311),
    .X(o[33]));
 sky130_fd_sc_hd__buf_2 output312 (.A(net312),
    .X(o[34]));
 sky130_fd_sc_hd__buf_2 output313 (.A(net313),
    .X(o[35]));
 sky130_fd_sc_hd__buf_2 output314 (.A(net314),
    .X(o[36]));
 sky130_fd_sc_hd__buf_2 output315 (.A(net315),
    .X(o[37]));
 sky130_fd_sc_hd__buf_2 output316 (.A(net316),
    .X(o[38]));
 sky130_fd_sc_hd__buf_2 output317 (.A(net317),
    .X(o[39]));
 sky130_fd_sc_hd__buf_2 output318 (.A(net318),
    .X(o[3]));
 sky130_fd_sc_hd__buf_2 output319 (.A(net319),
    .X(o[40]));
 sky130_fd_sc_hd__buf_2 output320 (.A(net320),
    .X(o[41]));
 sky130_fd_sc_hd__buf_2 output321 (.A(net321),
    .X(o[42]));
 sky130_fd_sc_hd__buf_2 output322 (.A(net322),
    .X(o[43]));
 sky130_fd_sc_hd__buf_2 output323 (.A(net323),
    .X(o[44]));
 sky130_fd_sc_hd__buf_2 output324 (.A(net324),
    .X(o[45]));
 sky130_fd_sc_hd__buf_2 output325 (.A(net325),
    .X(o[46]));
 sky130_fd_sc_hd__buf_2 output326 (.A(net326),
    .X(o[47]));
 sky130_fd_sc_hd__buf_2 output327 (.A(net327),
    .X(o[48]));
 sky130_fd_sc_hd__buf_2 output328 (.A(net328),
    .X(o[49]));
 sky130_fd_sc_hd__buf_2 output329 (.A(net329),
    .X(o[4]));
 sky130_fd_sc_hd__buf_2 output330 (.A(net330),
    .X(o[50]));
 sky130_fd_sc_hd__buf_2 output331 (.A(net331),
    .X(o[51]));
 sky130_fd_sc_hd__buf_2 output332 (.A(net332),
    .X(o[52]));
 sky130_fd_sc_hd__buf_2 output333 (.A(net333),
    .X(o[53]));
 sky130_fd_sc_hd__buf_2 output334 (.A(net334),
    .X(o[54]));
 sky130_fd_sc_hd__buf_2 output335 (.A(net335),
    .X(o[55]));
 sky130_fd_sc_hd__buf_2 output336 (.A(net336),
    .X(o[56]));
 sky130_fd_sc_hd__buf_2 output337 (.A(net337),
    .X(o[57]));
 sky130_fd_sc_hd__buf_2 output338 (.A(net338),
    .X(o[58]));
 sky130_fd_sc_hd__buf_2 output339 (.A(net339),
    .X(o[59]));
 sky130_fd_sc_hd__buf_2 output340 (.A(net340),
    .X(o[5]));
 sky130_fd_sc_hd__buf_2 output341 (.A(net341),
    .X(o[60]));
 sky130_fd_sc_hd__buf_2 output342 (.A(net342),
    .X(o[61]));
 sky130_fd_sc_hd__buf_2 output343 (.A(net343),
    .X(o[62]));
 sky130_fd_sc_hd__buf_2 output344 (.A(net344),
    .X(o[63]));
 sky130_fd_sc_hd__buf_2 output345 (.A(net345),
    .X(o[64]));
 sky130_fd_sc_hd__buf_2 output346 (.A(net346),
    .X(o[65]));
 sky130_fd_sc_hd__buf_2 output347 (.A(net347),
    .X(o[66]));
 sky130_fd_sc_hd__buf_2 output348 (.A(net348),
    .X(o[67]));
 sky130_fd_sc_hd__buf_2 output349 (.A(net349),
    .X(o[68]));
 sky130_fd_sc_hd__buf_2 output350 (.A(net350),
    .X(o[69]));
 sky130_fd_sc_hd__buf_2 output351 (.A(net351),
    .X(o[6]));
 sky130_fd_sc_hd__buf_2 output352 (.A(net352),
    .X(o[70]));
 sky130_fd_sc_hd__buf_2 output353 (.A(net353),
    .X(o[71]));
 sky130_fd_sc_hd__buf_2 output354 (.A(net354),
    .X(o[72]));
 sky130_fd_sc_hd__buf_2 output355 (.A(net355),
    .X(o[73]));
 sky130_fd_sc_hd__buf_2 output356 (.A(net356),
    .X(o[74]));
 sky130_fd_sc_hd__buf_2 output357 (.A(net357),
    .X(o[75]));
 sky130_fd_sc_hd__buf_2 output358 (.A(net358),
    .X(o[76]));
 sky130_fd_sc_hd__buf_2 output359 (.A(net359),
    .X(o[77]));
 sky130_fd_sc_hd__buf_2 output360 (.A(net360),
    .X(o[78]));
 sky130_fd_sc_hd__buf_2 output361 (.A(net361),
    .X(o[79]));
 sky130_fd_sc_hd__buf_2 output362 (.A(net362),
    .X(o[7]));
 sky130_fd_sc_hd__buf_2 output363 (.A(net363),
    .X(o[80]));
 sky130_fd_sc_hd__buf_2 output364 (.A(net364),
    .X(o[81]));
 sky130_fd_sc_hd__buf_2 output365 (.A(net365),
    .X(o[82]));
 sky130_fd_sc_hd__buf_2 output366 (.A(net366),
    .X(o[83]));
 sky130_fd_sc_hd__buf_2 output367 (.A(net367),
    .X(o[84]));
 sky130_fd_sc_hd__buf_2 output368 (.A(net368),
    .X(o[85]));
 sky130_fd_sc_hd__buf_2 output369 (.A(net369),
    .X(o[86]));
 sky130_fd_sc_hd__buf_2 output370 (.A(net370),
    .X(o[87]));
 sky130_fd_sc_hd__buf_2 output371 (.A(net371),
    .X(o[88]));
 sky130_fd_sc_hd__buf_2 output372 (.A(net372),
    .X(o[89]));
 sky130_fd_sc_hd__buf_2 output373 (.A(net373),
    .X(o[8]));
 sky130_fd_sc_hd__buf_2 output374 (.A(net374),
    .X(o[90]));
 sky130_fd_sc_hd__buf_2 output375 (.A(net375),
    .X(o[91]));
 sky130_fd_sc_hd__buf_2 output376 (.A(net376),
    .X(o[92]));
 sky130_fd_sc_hd__buf_2 output377 (.A(net377),
    .X(o[93]));
 sky130_fd_sc_hd__buf_2 output378 (.A(net378),
    .X(o[94]));
 sky130_fd_sc_hd__buf_2 output379 (.A(net379),
    .X(o[95]));
 sky130_fd_sc_hd__buf_2 output380 (.A(net380),
    .X(o[96]));
 sky130_fd_sc_hd__buf_2 output381 (.A(net381),
    .X(o[97]));
 sky130_fd_sc_hd__buf_2 output382 (.A(net382),
    .X(o[98]));
 sky130_fd_sc_hd__buf_2 output383 (.A(net383),
    .X(o[99]));
 sky130_fd_sc_hd__buf_2 output384 (.A(net384),
    .X(o[9]));
 sky130_fd_sc_hd__buf_4 fanout385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__buf_4 fanout386 (.A(net392),
    .X(net386));
 sky130_fd_sc_hd__buf_4 fanout387 (.A(net389),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_4 fanout388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_4 fanout389 (.A(net392),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_8 fanout390 (.A(net391),
    .X(net390));
 sky130_fd_sc_hd__buf_6 fanout391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__buf_8 fanout392 (.A(\sel_0$4897 ),
    .X(net392));
 sky130_fd_sc_hd__buf_4 fanout393 (.A(net394),
    .X(net393));
 sky130_fd_sc_hd__buf_6 fanout394 (.A(net400),
    .X(net394));
 sky130_fd_sc_hd__buf_4 fanout395 (.A(net400),
    .X(net395));
 sky130_fd_sc_hd__buf_4 fanout396 (.A(net398),
    .X(net396));
 sky130_fd_sc_hd__buf_4 fanout397 (.A(net398),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_4 fanout398 (.A(net399),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_8 fanout399 (.A(net400),
    .X(net399));
 sky130_fd_sc_hd__buf_6 fanout400 (.A(\sel_0$4827 ),
    .X(net400));
 sky130_fd_sc_hd__buf_4 fanout401 (.A(net402),
    .X(net401));
 sky130_fd_sc_hd__buf_4 fanout402 (.A(net408),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_8 fanout403 (.A(net408),
    .X(net403));
 sky130_fd_sc_hd__buf_4 fanout404 (.A(net407),
    .X(net404));
 sky130_fd_sc_hd__buf_2 fanout405 (.A(net406),
    .X(net405));
 sky130_fd_sc_hd__buf_4 fanout406 (.A(net407),
    .X(net406));
 sky130_fd_sc_hd__buf_6 fanout407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__buf_6 fanout408 (.A(\sel_0$4757 ),
    .X(net408));
 sky130_fd_sc_hd__buf_4 fanout409 (.A(net412),
    .X(net409));
 sky130_fd_sc_hd__buf_4 fanout410 (.A(net412),
    .X(net410));
 sky130_fd_sc_hd__buf_4 fanout411 (.A(net412),
    .X(net411));
 sky130_fd_sc_hd__buf_4 fanout412 (.A(net417),
    .X(net412));
 sky130_fd_sc_hd__buf_4 fanout413 (.A(net414),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_4 fanout414 (.A(net415),
    .X(net414));
 sky130_fd_sc_hd__buf_4 fanout415 (.A(net417),
    .X(net415));
 sky130_fd_sc_hd__buf_4 fanout416 (.A(net417),
    .X(net416));
 sky130_fd_sc_hd__buf_6 fanout417 (.A(\sel_0$4687 ),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_8 fanout418 (.A(net421),
    .X(net418));
 sky130_fd_sc_hd__buf_4 fanout419 (.A(net421),
    .X(net419));
 sky130_fd_sc_hd__buf_4 fanout420 (.A(net421),
    .X(net420));
 sky130_fd_sc_hd__buf_6 fanout421 (.A(\sel_0$6577 ),
    .X(net421));
 sky130_fd_sc_hd__buf_4 fanout422 (.A(net425),
    .X(net422));
 sky130_fd_sc_hd__buf_4 fanout423 (.A(net425),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_4 fanout424 (.A(net425),
    .X(net424));
 sky130_fd_sc_hd__buf_4 fanout425 (.A(\sel_0$6577 ),
    .X(net425));
 sky130_fd_sc_hd__buf_4 fanout426 (.A(net427),
    .X(net426));
 sky130_fd_sc_hd__buf_6 fanout427 (.A(net428),
    .X(net427));
 sky130_fd_sc_hd__buf_6 fanout428 (.A(net433),
    .X(net428));
 sky130_fd_sc_hd__buf_4 fanout429 (.A(net430),
    .X(net429));
 sky130_fd_sc_hd__buf_4 fanout430 (.A(net431),
    .X(net430));
 sky130_fd_sc_hd__buf_4 fanout431 (.A(net433),
    .X(net431));
 sky130_fd_sc_hd__buf_6 fanout432 (.A(net433),
    .X(net432));
 sky130_fd_sc_hd__buf_6 fanout433 (.A(\sel_0$4617 ),
    .X(net433));
 sky130_fd_sc_hd__buf_4 fanout434 (.A(net437),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_4 fanout435 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__buf_4 fanout436 (.A(net437),
    .X(net436));
 sky130_fd_sc_hd__buf_4 fanout437 (.A(net441),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_4 fanout438 (.A(net441),
    .X(net438));
 sky130_fd_sc_hd__buf_4 fanout439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__buf_4 fanout440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_4 fanout441 (.A(\sel_0$6507 ),
    .X(net441));
 sky130_fd_sc_hd__buf_4 fanout442 (.A(net450),
    .X(net442));
 sky130_fd_sc_hd__buf_2 fanout443 (.A(net450),
    .X(net443));
 sky130_fd_sc_hd__buf_4 fanout444 (.A(net445),
    .X(net444));
 sky130_fd_sc_hd__buf_4 fanout445 (.A(net450),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_4 fanout446 (.A(net447),
    .X(net446));
 sky130_fd_sc_hd__buf_2 fanout447 (.A(net449),
    .X(net447));
 sky130_fd_sc_hd__buf_4 fanout448 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__buf_6 fanout449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__buf_6 fanout450 (.A(sel_0),
    .X(net450));
 sky130_fd_sc_hd__buf_4 fanout451 (.A(net459),
    .X(net451));
 sky130_fd_sc_hd__buf_2 fanout452 (.A(net459),
    .X(net452));
 sky130_fd_sc_hd__buf_4 fanout453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__buf_4 fanout454 (.A(net459),
    .X(net454));
 sky130_fd_sc_hd__buf_6 fanout455 (.A(net458),
    .X(net455));
 sky130_fd_sc_hd__buf_4 fanout456 (.A(net458),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_4 fanout457 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__buf_4 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_4 fanout459 (.A(\sel_0$6437 ),
    .X(net459));
 sky130_fd_sc_hd__buf_4 fanout460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_4 fanout461 (.A(\sel_0$6367 ),
    .X(net461));
 sky130_fd_sc_hd__buf_4 fanout462 (.A(net463),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_8 fanout463 (.A(\sel_0$6367 ),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_8 fanout464 (.A(net467),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_8 fanout465 (.A(net467),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_4 fanout466 (.A(net467),
    .X(net466));
 sky130_fd_sc_hd__buf_6 fanout467 (.A(\sel_0$6367 ),
    .X(net467));
 sky130_fd_sc_hd__buf_6 fanout468 (.A(net471),
    .X(net468));
 sky130_fd_sc_hd__buf_4 fanout469 (.A(net471),
    .X(net469));
 sky130_fd_sc_hd__clkbuf_4 fanout470 (.A(net471),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_4 fanout471 (.A(\sel_0$6297 ),
    .X(net471));
 sky130_fd_sc_hd__buf_6 fanout472 (.A(net475),
    .X(net472));
 sky130_fd_sc_hd__buf_4 fanout473 (.A(net475),
    .X(net473));
 sky130_fd_sc_hd__buf_4 fanout474 (.A(net475),
    .X(net474));
 sky130_fd_sc_hd__buf_6 fanout475 (.A(\sel_0$6297 ),
    .X(net475));
 sky130_fd_sc_hd__buf_6 fanout476 (.A(net479),
    .X(net476));
 sky130_fd_sc_hd__buf_4 fanout477 (.A(net479),
    .X(net477));
 sky130_fd_sc_hd__buf_2 fanout478 (.A(net479),
    .X(net478));
 sky130_fd_sc_hd__buf_4 fanout479 (.A(\sel_0$6227 ),
    .X(net479));
 sky130_fd_sc_hd__buf_4 fanout480 (.A(net481),
    .X(net480));
 sky130_fd_sc_hd__buf_4 fanout481 (.A(\sel_0$6227 ),
    .X(net481));
 sky130_fd_sc_hd__buf_4 fanout482 (.A(net483),
    .X(net482));
 sky130_fd_sc_hd__buf_4 fanout483 (.A(\sel_0$6227 ),
    .X(net483));
 sky130_fd_sc_hd__buf_4 fanout484 (.A(net487),
    .X(net484));
 sky130_fd_sc_hd__buf_4 fanout485 (.A(net487),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_4 fanout486 (.A(net487),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_8 fanout487 (.A(\sel_0$6157 ),
    .X(net487));
 sky130_fd_sc_hd__buf_4 fanout488 (.A(net492),
    .X(net488));
 sky130_fd_sc_hd__buf_4 fanout489 (.A(net491),
    .X(net489));
 sky130_fd_sc_hd__buf_4 fanout490 (.A(net491),
    .X(net490));
 sky130_fd_sc_hd__buf_2 fanout491 (.A(net492),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_8 fanout492 (.A(\sel_0$6157 ),
    .X(net492));
 sky130_fd_sc_hd__buf_4 fanout493 (.A(net496),
    .X(net493));
 sky130_fd_sc_hd__buf_4 fanout494 (.A(net495),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_8 fanout495 (.A(net496),
    .X(net495));
 sky130_fd_sc_hd__buf_4 fanout496 (.A(\sel_0$6087 ),
    .X(net496));
 sky130_fd_sc_hd__buf_4 fanout497 (.A(net500),
    .X(net497));
 sky130_fd_sc_hd__buf_4 fanout498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__buf_6 fanout499 (.A(net500),
    .X(net499));
 sky130_fd_sc_hd__buf_6 fanout500 (.A(\sel_0$6087 ),
    .X(net500));
 sky130_fd_sc_hd__buf_4 fanout501 (.A(net502),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_4 fanout502 (.A(net509),
    .X(net502));
 sky130_fd_sc_hd__buf_4 fanout503 (.A(net509),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_4 fanout504 (.A(net509),
    .X(net504));
 sky130_fd_sc_hd__buf_4 fanout505 (.A(net506),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_4 fanout506 (.A(net509),
    .X(net506));
 sky130_fd_sc_hd__buf_4 fanout507 (.A(net508),
    .X(net507));
 sky130_fd_sc_hd__buf_4 fanout508 (.A(net509),
    .X(net508));
 sky130_fd_sc_hd__buf_4 fanout509 (.A(\sel_0$6017 ),
    .X(net509));
 sky130_fd_sc_hd__buf_4 fanout510 (.A(net518),
    .X(net510));
 sky130_fd_sc_hd__buf_4 fanout511 (.A(net518),
    .X(net511));
 sky130_fd_sc_hd__buf_4 fanout512 (.A(net518),
    .X(net512));
 sky130_fd_sc_hd__buf_4 fanout513 (.A(net518),
    .X(net513));
 sky130_fd_sc_hd__buf_4 fanout514 (.A(net517),
    .X(net514));
 sky130_fd_sc_hd__buf_4 fanout515 (.A(net516),
    .X(net515));
 sky130_fd_sc_hd__buf_4 fanout516 (.A(net517),
    .X(net516));
 sky130_fd_sc_hd__clkbuf_8 fanout517 (.A(net518),
    .X(net517));
 sky130_fd_sc_hd__buf_4 fanout518 (.A(\sel_0$5947 ),
    .X(net518));
 sky130_fd_sc_hd__buf_4 fanout519 (.A(net520),
    .X(net519));
 sky130_fd_sc_hd__buf_4 fanout520 (.A(\sel_0$5877 ),
    .X(net520));
 sky130_fd_sc_hd__buf_4 fanout521 (.A(net522),
    .X(net521));
 sky130_fd_sc_hd__buf_6 fanout522 (.A(\sel_0$5877 ),
    .X(net522));
 sky130_fd_sc_hd__buf_4 fanout523 (.A(net526),
    .X(net523));
 sky130_fd_sc_hd__buf_6 fanout524 (.A(net525),
    .X(net524));
 sky130_fd_sc_hd__buf_4 fanout525 (.A(net526),
    .X(net525));
 sky130_fd_sc_hd__clkbuf_8 fanout526 (.A(\sel_0$5877 ),
    .X(net526));
 sky130_fd_sc_hd__buf_4 fanout527 (.A(net530),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_4 fanout528 (.A(net530),
    .X(net528));
 sky130_fd_sc_hd__buf_4 fanout529 (.A(net530),
    .X(net529));
 sky130_fd_sc_hd__buf_6 fanout530 (.A(\sel_0$4547 ),
    .X(net530));
 sky130_fd_sc_hd__buf_4 fanout531 (.A(net532),
    .X(net531));
 sky130_fd_sc_hd__buf_4 fanout532 (.A(net534),
    .X(net532));
 sky130_fd_sc_hd__buf_4 fanout533 (.A(net534),
    .X(net533));
 sky130_fd_sc_hd__buf_4 fanout534 (.A(\sel_0$4547 ),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_8 fanout535 (.A(net536),
    .X(net535));
 sky130_fd_sc_hd__buf_4 fanout536 (.A(net542),
    .X(net536));
 sky130_fd_sc_hd__clkbuf_8 fanout537 (.A(net538),
    .X(net537));
 sky130_fd_sc_hd__buf_4 fanout538 (.A(net542),
    .X(net538));
 sky130_fd_sc_hd__buf_4 fanout539 (.A(net542),
    .X(net539));
 sky130_fd_sc_hd__buf_4 fanout540 (.A(net541),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_4 fanout541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__buf_8 fanout542 (.A(\sel_0$5807 ),
    .X(net542));
 sky130_fd_sc_hd__buf_4 fanout543 (.A(net544),
    .X(net543));
 sky130_fd_sc_hd__buf_6 fanout544 (.A(net550),
    .X(net544));
 sky130_fd_sc_hd__buf_6 fanout545 (.A(net546),
    .X(net545));
 sky130_fd_sc_hd__buf_6 fanout546 (.A(net550),
    .X(net546));
 sky130_fd_sc_hd__buf_4 fanout547 (.A(net548),
    .X(net547));
 sky130_fd_sc_hd__buf_4 fanout548 (.A(net550),
    .X(net548));
 sky130_fd_sc_hd__buf_4 fanout549 (.A(net550),
    .X(net549));
 sky130_fd_sc_hd__buf_6 fanout550 (.A(\sel_0$5737 ),
    .X(net550));
 sky130_fd_sc_hd__buf_4 fanout551 (.A(net553),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_4 fanout552 (.A(net553),
    .X(net552));
 sky130_fd_sc_hd__buf_4 fanout553 (.A(net559),
    .X(net553));
 sky130_fd_sc_hd__buf_4 fanout554 (.A(net559),
    .X(net554));
 sky130_fd_sc_hd__buf_4 fanout555 (.A(net556),
    .X(net555));
 sky130_fd_sc_hd__buf_6 fanout556 (.A(net558),
    .X(net556));
 sky130_fd_sc_hd__buf_4 fanout557 (.A(net558),
    .X(net557));
 sky130_fd_sc_hd__buf_4 fanout558 (.A(net559),
    .X(net558));
 sky130_fd_sc_hd__buf_6 fanout559 (.A(\sel_0$5667 ),
    .X(net559));
 sky130_fd_sc_hd__buf_4 fanout560 (.A(net562),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_2 fanout561 (.A(net562),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_8 fanout562 (.A(net568),
    .X(net562));
 sky130_fd_sc_hd__buf_4 fanout563 (.A(net564),
    .X(net563));
 sky130_fd_sc_hd__buf_4 fanout564 (.A(net568),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_8 fanout565 (.A(net568),
    .X(net565));
 sky130_fd_sc_hd__buf_4 fanout566 (.A(net568),
    .X(net566));
 sky130_fd_sc_hd__clkbuf_8 fanout567 (.A(net568),
    .X(net567));
 sky130_fd_sc_hd__buf_8 fanout568 (.A(\sel_0$5597 ),
    .X(net568));
 sky130_fd_sc_hd__buf_6 fanout569 (.A(net570),
    .X(net569));
 sky130_fd_sc_hd__buf_8 fanout570 (.A(\sel_0$5527 ),
    .X(net570));
 sky130_fd_sc_hd__buf_4 fanout571 (.A(net572),
    .X(net571));
 sky130_fd_sc_hd__buf_6 fanout572 (.A(\sel_0$5527 ),
    .X(net572));
 sky130_fd_sc_hd__buf_4 fanout573 (.A(net574),
    .X(net573));
 sky130_fd_sc_hd__buf_4 fanout574 (.A(net575),
    .X(net574));
 sky130_fd_sc_hd__buf_6 fanout575 (.A(\sel_0$5527 ),
    .X(net575));
 sky130_fd_sc_hd__buf_4 fanout576 (.A(net583),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_4 fanout577 (.A(net583),
    .X(net577));
 sky130_fd_sc_hd__buf_4 fanout578 (.A(net579),
    .X(net578));
 sky130_fd_sc_hd__buf_6 fanout579 (.A(net583),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_4 fanout580 (.A(net581),
    .X(net580));
 sky130_fd_sc_hd__buf_6 fanout581 (.A(net582),
    .X(net581));
 sky130_fd_sc_hd__buf_6 fanout582 (.A(net583),
    .X(net582));
 sky130_fd_sc_hd__buf_6 fanout583 (.A(\sel_0$5457 ),
    .X(net583));
 sky130_fd_sc_hd__buf_4 fanout584 (.A(net586),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_4 fanout585 (.A(net586),
    .X(net585));
 sky130_fd_sc_hd__buf_4 fanout586 (.A(net592),
    .X(net586));
 sky130_fd_sc_hd__buf_4 fanout587 (.A(net588),
    .X(net587));
 sky130_fd_sc_hd__buf_6 fanout588 (.A(net592),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_8 fanout589 (.A(net592),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_4 fanout590 (.A(net592),
    .X(net590));
 sky130_fd_sc_hd__buf_4 fanout591 (.A(net592),
    .X(net591));
 sky130_fd_sc_hd__buf_6 fanout592 (.A(\sel_0$5387 ),
    .X(net592));
 sky130_fd_sc_hd__buf_4 fanout593 (.A(net595),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_2 fanout594 (.A(net595),
    .X(net594));
 sky130_fd_sc_hd__buf_2 fanout595 (.A(net601),
    .X(net595));
 sky130_fd_sc_hd__buf_4 fanout596 (.A(net597),
    .X(net596));
 sky130_fd_sc_hd__buf_6 fanout597 (.A(net601),
    .X(net597));
 sky130_fd_sc_hd__buf_4 fanout598 (.A(net600),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_4 fanout599 (.A(net600),
    .X(net599));
 sky130_fd_sc_hd__buf_6 fanout600 (.A(net601),
    .X(net600));
 sky130_fd_sc_hd__buf_6 fanout601 (.A(\sel_0$5317 ),
    .X(net601));
 sky130_fd_sc_hd__buf_4 fanout602 (.A(net604),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_4 fanout603 (.A(net604),
    .X(net603));
 sky130_fd_sc_hd__buf_4 fanout604 (.A(\sel_0$5247 ),
    .X(net604));
 sky130_fd_sc_hd__buf_4 fanout605 (.A(net606),
    .X(net605));
 sky130_fd_sc_hd__buf_6 fanout606 (.A(\sel_0$5247 ),
    .X(net606));
 sky130_fd_sc_hd__buf_6 fanout607 (.A(net609),
    .X(net607));
 sky130_fd_sc_hd__clkbuf_4 fanout608 (.A(net609),
    .X(net608));
 sky130_fd_sc_hd__buf_6 fanout609 (.A(\sel_0$5247 ),
    .X(net609));
 sky130_fd_sc_hd__buf_4 fanout610 (.A(net612),
    .X(net610));
 sky130_fd_sc_hd__buf_2 fanout611 (.A(net612),
    .X(net611));
 sky130_fd_sc_hd__buf_6 fanout612 (.A(\sel_0$5177 ),
    .X(net612));
 sky130_fd_sc_hd__buf_4 fanout613 (.A(net615),
    .X(net613));
 sky130_fd_sc_hd__buf_2 fanout614 (.A(net615),
    .X(net614));
 sky130_fd_sc_hd__buf_4 fanout615 (.A(\sel_0$5177 ),
    .X(net615));
 sky130_fd_sc_hd__buf_4 fanout616 (.A(net618),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_4 fanout617 (.A(net618),
    .X(net617));
 sky130_fd_sc_hd__buf_6 fanout618 (.A(\sel_0$5177 ),
    .X(net618));
 sky130_fd_sc_hd__buf_4 fanout619 (.A(net622),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_4 fanout620 (.A(net622),
    .X(net620));
 sky130_fd_sc_hd__buf_4 fanout621 (.A(net622),
    .X(net621));
 sky130_fd_sc_hd__clkbuf_8 fanout622 (.A(\sel_0$4477 ),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_4 fanout623 (.A(net625),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_4 fanout624 (.A(net625),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_4 fanout625 (.A(\sel_0$4477 ),
    .X(net625));
 sky130_fd_sc_hd__buf_4 fanout626 (.A(\sel_0$4477 ),
    .X(net626));
 sky130_fd_sc_hd__buf_4 fanout627 (.A(net628),
    .X(net627));
 sky130_fd_sc_hd__buf_6 fanout628 (.A(net631),
    .X(net628));
 sky130_fd_sc_hd__clkbuf_8 fanout629 (.A(net630),
    .X(net629));
 sky130_fd_sc_hd__buf_6 fanout630 (.A(net631),
    .X(net630));
 sky130_fd_sc_hd__buf_4 fanout631 (.A(\sel_0$5107 ),
    .X(net631));
 sky130_fd_sc_hd__buf_4 fanout632 (.A(net634),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_4 fanout633 (.A(net634),
    .X(net633));
 sky130_fd_sc_hd__buf_6 fanout634 (.A(\sel_0$5107 ),
    .X(net634));
 sky130_fd_sc_hd__buf_4 fanout635 (.A(net636),
    .X(net635));
 sky130_fd_sc_hd__buf_6 fanout636 (.A(net639),
    .X(net636));
 sky130_fd_sc_hd__buf_4 fanout637 (.A(net638),
    .X(net637));
 sky130_fd_sc_hd__buf_6 fanout638 (.A(net639),
    .X(net638));
 sky130_fd_sc_hd__buf_6 fanout639 (.A(\sel_0$5037 ),
    .X(net639));
 sky130_fd_sc_hd__buf_4 fanout640 (.A(net642),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_4 fanout641 (.A(net642),
    .X(net641));
 sky130_fd_sc_hd__buf_6 fanout642 (.A(\sel_0$5037 ),
    .X(net642));
 sky130_fd_sc_hd__buf_4 fanout643 (.A(net644),
    .X(net643));
 sky130_fd_sc_hd__buf_6 fanout644 (.A(net647),
    .X(net644));
 sky130_fd_sc_hd__clkbuf_8 fanout645 (.A(net646),
    .X(net645));
 sky130_fd_sc_hd__buf_6 fanout646 (.A(net647),
    .X(net646));
 sky130_fd_sc_hd__buf_4 fanout647 (.A(\sel_0$4967 ),
    .X(net647));
 sky130_fd_sc_hd__buf_6 fanout648 (.A(net650),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_4 fanout649 (.A(net650),
    .X(net649));
 sky130_fd_sc_hd__buf_6 fanout650 (.A(\sel_0$4967 ),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_4 fanout651 (.A(net652),
    .X(net651));
 sky130_fd_sc_hd__buf_4 fanout652 (.A(net658),
    .X(net652));
 sky130_fd_sc_hd__buf_4 fanout653 (.A(net655),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_4 fanout654 (.A(net655),
    .X(net654));
 sky130_fd_sc_hd__clkbuf_4 fanout655 (.A(net658),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_8 fanout656 (.A(net657),
    .X(net656));
 sky130_fd_sc_hd__buf_6 fanout657 (.A(net658),
    .X(net657));
 sky130_fd_sc_hd__buf_8 fanout658 (.A(\sel_1$4898 ),
    .X(net658));
 sky130_fd_sc_hd__buf_4 fanout659 (.A(net660),
    .X(net659));
 sky130_fd_sc_hd__buf_6 fanout660 (.A(net666),
    .X(net660));
 sky130_fd_sc_hd__buf_4 fanout661 (.A(net666),
    .X(net661));
 sky130_fd_sc_hd__buf_4 fanout662 (.A(net664),
    .X(net662));
 sky130_fd_sc_hd__buf_4 fanout663 (.A(net664),
    .X(net663));
 sky130_fd_sc_hd__clkbuf_4 fanout664 (.A(net665),
    .X(net664));
 sky130_fd_sc_hd__clkbuf_8 fanout665 (.A(net666),
    .X(net665));
 sky130_fd_sc_hd__buf_6 fanout666 (.A(\sel_1$4828 ),
    .X(net666));
 sky130_fd_sc_hd__buf_4 fanout667 (.A(net668),
    .X(net667));
 sky130_fd_sc_hd__buf_4 fanout668 (.A(net674),
    .X(net668));
 sky130_fd_sc_hd__buf_4 fanout669 (.A(net674),
    .X(net669));
 sky130_fd_sc_hd__buf_4 fanout670 (.A(net673),
    .X(net670));
 sky130_fd_sc_hd__buf_2 fanout671 (.A(net672),
    .X(net671));
 sky130_fd_sc_hd__buf_4 fanout672 (.A(net673),
    .X(net672));
 sky130_fd_sc_hd__buf_6 fanout673 (.A(net674),
    .X(net673));
 sky130_fd_sc_hd__buf_6 fanout674 (.A(\sel_1$4758 ),
    .X(net674));
 sky130_fd_sc_hd__buf_4 fanout675 (.A(net678),
    .X(net675));
 sky130_fd_sc_hd__buf_4 fanout676 (.A(net678),
    .X(net676));
 sky130_fd_sc_hd__buf_4 fanout677 (.A(net678),
    .X(net677));
 sky130_fd_sc_hd__buf_4 fanout678 (.A(net683),
    .X(net678));
 sky130_fd_sc_hd__buf_4 fanout679 (.A(net680),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_4 fanout680 (.A(net681),
    .X(net680));
 sky130_fd_sc_hd__buf_4 fanout681 (.A(net683),
    .X(net681));
 sky130_fd_sc_hd__buf_4 fanout682 (.A(net683),
    .X(net682));
 sky130_fd_sc_hd__buf_6 fanout683 (.A(\sel_1$4688 ),
    .X(net683));
 sky130_fd_sc_hd__buf_4 fanout684 (.A(net692),
    .X(net684));
 sky130_fd_sc_hd__buf_2 fanout685 (.A(net692),
    .X(net685));
 sky130_fd_sc_hd__buf_4 fanout686 (.A(net687),
    .X(net686));
 sky130_fd_sc_hd__buf_4 fanout687 (.A(net692),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_4 fanout688 (.A(net689),
    .X(net688));
 sky130_fd_sc_hd__buf_2 fanout689 (.A(net691),
    .X(net689));
 sky130_fd_sc_hd__buf_4 fanout690 (.A(net691),
    .X(net690));
 sky130_fd_sc_hd__buf_6 fanout691 (.A(net692),
    .X(net691));
 sky130_fd_sc_hd__buf_6 fanout692 (.A(sel_1),
    .X(net692));
 sky130_fd_sc_hd__clkbuf_4 fanout693 (.A(net694),
    .X(net693));
 sky130_fd_sc_hd__buf_4 fanout694 (.A(net695),
    .X(net694));
 sky130_fd_sc_hd__buf_4 fanout695 (.A(\sel_1$6648 ),
    .X(net695));
 sky130_fd_sc_hd__buf_4 fanout696 (.A(net699),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_4 fanout697 (.A(net699),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_4 fanout698 (.A(net699),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_8 fanout699 (.A(\sel_1$6648 ),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_8 fanout700 (.A(net703),
    .X(net700));
 sky130_fd_sc_hd__buf_4 fanout701 (.A(net703),
    .X(net701));
 sky130_fd_sc_hd__buf_4 fanout702 (.A(net703),
    .X(net702));
 sky130_fd_sc_hd__buf_6 fanout703 (.A(\sel_1$6578 ),
    .X(net703));
 sky130_fd_sc_hd__buf_4 fanout704 (.A(net707),
    .X(net704));
 sky130_fd_sc_hd__buf_4 fanout705 (.A(net707),
    .X(net705));
 sky130_fd_sc_hd__clkbuf_4 fanout706 (.A(net707),
    .X(net706));
 sky130_fd_sc_hd__buf_4 fanout707 (.A(\sel_1$6578 ),
    .X(net707));
 sky130_fd_sc_hd__buf_4 fanout708 (.A(net709),
    .X(net708));
 sky130_fd_sc_hd__buf_6 fanout709 (.A(net710),
    .X(net709));
 sky130_fd_sc_hd__buf_6 fanout710 (.A(net715),
    .X(net710));
 sky130_fd_sc_hd__buf_4 fanout711 (.A(net712),
    .X(net711));
 sky130_fd_sc_hd__buf_4 fanout712 (.A(net713),
    .X(net712));
 sky130_fd_sc_hd__buf_4 fanout713 (.A(net715),
    .X(net713));
 sky130_fd_sc_hd__buf_6 fanout714 (.A(net715),
    .X(net714));
 sky130_fd_sc_hd__buf_6 fanout715 (.A(\sel_1$4618 ),
    .X(net715));
 sky130_fd_sc_hd__buf_4 fanout716 (.A(net719),
    .X(net716));
 sky130_fd_sc_hd__clkbuf_4 fanout717 (.A(net718),
    .X(net717));
 sky130_fd_sc_hd__buf_4 fanout718 (.A(net719),
    .X(net718));
 sky130_fd_sc_hd__buf_4 fanout719 (.A(net723),
    .X(net719));
 sky130_fd_sc_hd__clkbuf_4 fanout720 (.A(net723),
    .X(net720));
 sky130_fd_sc_hd__buf_4 fanout721 (.A(net722),
    .X(net721));
 sky130_fd_sc_hd__buf_4 fanout722 (.A(net723),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_4 fanout723 (.A(\sel_1$6508 ),
    .X(net723));
 sky130_fd_sc_hd__buf_4 fanout724 (.A(net732),
    .X(net724));
 sky130_fd_sc_hd__buf_2 fanout725 (.A(net732),
    .X(net725));
 sky130_fd_sc_hd__buf_4 fanout726 (.A(net727),
    .X(net726));
 sky130_fd_sc_hd__buf_4 fanout727 (.A(net732),
    .X(net727));
 sky130_fd_sc_hd__buf_6 fanout728 (.A(net731),
    .X(net728));
 sky130_fd_sc_hd__buf_4 fanout729 (.A(net731),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_4 fanout730 (.A(net731),
    .X(net730));
 sky130_fd_sc_hd__buf_4 fanout731 (.A(net732),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_4 fanout732 (.A(\sel_1$6438 ),
    .X(net732));
 sky130_fd_sc_hd__buf_4 fanout733 (.A(net734),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_4 fanout734 (.A(\sel_1$6368 ),
    .X(net734));
 sky130_fd_sc_hd__buf_4 fanout735 (.A(net736),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_8 fanout736 (.A(\sel_1$6368 ),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_8 fanout737 (.A(net740),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_8 fanout738 (.A(net740),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_4 fanout739 (.A(net740),
    .X(net739));
 sky130_fd_sc_hd__buf_6 fanout740 (.A(\sel_1$6368 ),
    .X(net740));
 sky130_fd_sc_hd__buf_6 fanout741 (.A(net744),
    .X(net741));
 sky130_fd_sc_hd__buf_4 fanout742 (.A(net744),
    .X(net742));
 sky130_fd_sc_hd__clkbuf_4 fanout743 (.A(net744),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_4 fanout744 (.A(\sel_1$6298 ),
    .X(net744));
 sky130_fd_sc_hd__buf_6 fanout745 (.A(net748),
    .X(net745));
 sky130_fd_sc_hd__buf_4 fanout746 (.A(net748),
    .X(net746));
 sky130_fd_sc_hd__buf_4 fanout747 (.A(net748),
    .X(net747));
 sky130_fd_sc_hd__buf_6 fanout748 (.A(\sel_1$6298 ),
    .X(net748));
 sky130_fd_sc_hd__buf_6 fanout749 (.A(net752),
    .X(net749));
 sky130_fd_sc_hd__buf_4 fanout750 (.A(net752),
    .X(net750));
 sky130_fd_sc_hd__buf_2 fanout751 (.A(net752),
    .X(net751));
 sky130_fd_sc_hd__buf_4 fanout752 (.A(\sel_1$6228 ),
    .X(net752));
 sky130_fd_sc_hd__buf_4 fanout753 (.A(net754),
    .X(net753));
 sky130_fd_sc_hd__buf_4 fanout754 (.A(\sel_1$6228 ),
    .X(net754));
 sky130_fd_sc_hd__buf_4 fanout755 (.A(net756),
    .X(net755));
 sky130_fd_sc_hd__buf_4 fanout756 (.A(\sel_1$6228 ),
    .X(net756));
 sky130_fd_sc_hd__buf_4 fanout757 (.A(net760),
    .X(net757));
 sky130_fd_sc_hd__buf_4 fanout758 (.A(net760),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_4 fanout759 (.A(net760),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_8 fanout760 (.A(\sel_1$6158 ),
    .X(net760));
 sky130_fd_sc_hd__buf_4 fanout761 (.A(net765),
    .X(net761));
 sky130_fd_sc_hd__buf_4 fanout762 (.A(net764),
    .X(net762));
 sky130_fd_sc_hd__buf_4 fanout763 (.A(net764),
    .X(net763));
 sky130_fd_sc_hd__buf_2 fanout764 (.A(net765),
    .X(net764));
 sky130_fd_sc_hd__clkbuf_8 fanout765 (.A(\sel_1$6158 ),
    .X(net765));
 sky130_fd_sc_hd__buf_4 fanout766 (.A(net769),
    .X(net766));
 sky130_fd_sc_hd__buf_4 fanout767 (.A(net768),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_8 fanout768 (.A(net769),
    .X(net768));
 sky130_fd_sc_hd__buf_4 fanout769 (.A(\sel_1$6088 ),
    .X(net769));
 sky130_fd_sc_hd__buf_4 fanout770 (.A(net773),
    .X(net770));
 sky130_fd_sc_hd__buf_4 fanout771 (.A(net772),
    .X(net771));
 sky130_fd_sc_hd__buf_6 fanout772 (.A(net773),
    .X(net772));
 sky130_fd_sc_hd__buf_6 fanout773 (.A(\sel_1$6088 ),
    .X(net773));
 sky130_fd_sc_hd__buf_4 fanout774 (.A(net775),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_4 fanout775 (.A(net782),
    .X(net775));
 sky130_fd_sc_hd__buf_4 fanout776 (.A(net782),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_4 fanout777 (.A(net782),
    .X(net777));
 sky130_fd_sc_hd__buf_4 fanout778 (.A(net779),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_4 fanout779 (.A(net782),
    .X(net779));
 sky130_fd_sc_hd__buf_4 fanout780 (.A(net781),
    .X(net780));
 sky130_fd_sc_hd__buf_4 fanout781 (.A(net782),
    .X(net781));
 sky130_fd_sc_hd__clkbuf_8 fanout782 (.A(\sel_1$6018 ),
    .X(net782));
 sky130_fd_sc_hd__buf_4 fanout783 (.A(net791),
    .X(net783));
 sky130_fd_sc_hd__buf_4 fanout784 (.A(net791),
    .X(net784));
 sky130_fd_sc_hd__buf_4 fanout785 (.A(net791),
    .X(net785));
 sky130_fd_sc_hd__buf_4 fanout786 (.A(net791),
    .X(net786));
 sky130_fd_sc_hd__buf_4 fanout787 (.A(net790),
    .X(net787));
 sky130_fd_sc_hd__buf_4 fanout788 (.A(net789),
    .X(net788));
 sky130_fd_sc_hd__buf_4 fanout789 (.A(net790),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_8 fanout790 (.A(net791),
    .X(net790));
 sky130_fd_sc_hd__buf_4 fanout791 (.A(\sel_1$5948 ),
    .X(net791));
 sky130_fd_sc_hd__buf_4 fanout792 (.A(net793),
    .X(net792));
 sky130_fd_sc_hd__buf_4 fanout793 (.A(\sel_1$5878 ),
    .X(net793));
 sky130_fd_sc_hd__buf_4 fanout794 (.A(net795),
    .X(net794));
 sky130_fd_sc_hd__buf_6 fanout795 (.A(\sel_1$5878 ),
    .X(net795));
 sky130_fd_sc_hd__buf_4 fanout796 (.A(net799),
    .X(net796));
 sky130_fd_sc_hd__buf_6 fanout797 (.A(net798),
    .X(net797));
 sky130_fd_sc_hd__buf_4 fanout798 (.A(net799),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_8 fanout799 (.A(\sel_1$5878 ),
    .X(net799));
 sky130_fd_sc_hd__buf_4 fanout800 (.A(net803),
    .X(net800));
 sky130_fd_sc_hd__buf_2 fanout801 (.A(net803),
    .X(net801));
 sky130_fd_sc_hd__buf_4 fanout802 (.A(net803),
    .X(net802));
 sky130_fd_sc_hd__buf_6 fanout803 (.A(\sel_1$4548 ),
    .X(net803));
 sky130_fd_sc_hd__buf_4 fanout804 (.A(net805),
    .X(net804));
 sky130_fd_sc_hd__buf_4 fanout805 (.A(net807),
    .X(net805));
 sky130_fd_sc_hd__buf_4 fanout806 (.A(net807),
    .X(net806));
 sky130_fd_sc_hd__buf_4 fanout807 (.A(\sel_1$4548 ),
    .X(net807));
 sky130_fd_sc_hd__buf_4 fanout808 (.A(net809),
    .X(net808));
 sky130_fd_sc_hd__buf_4 fanout809 (.A(net815),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_8 fanout810 (.A(net811),
    .X(net810));
 sky130_fd_sc_hd__buf_4 fanout811 (.A(net815),
    .X(net811));
 sky130_fd_sc_hd__buf_4 fanout812 (.A(net815),
    .X(net812));
 sky130_fd_sc_hd__buf_4 fanout813 (.A(net814),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_4 fanout814 (.A(net815),
    .X(net814));
 sky130_fd_sc_hd__buf_8 fanout815 (.A(\sel_1$5808 ),
    .X(net815));
 sky130_fd_sc_hd__buf_4 fanout816 (.A(net817),
    .X(net816));
 sky130_fd_sc_hd__buf_6 fanout817 (.A(net823),
    .X(net817));
 sky130_fd_sc_hd__buf_6 fanout818 (.A(net819),
    .X(net818));
 sky130_fd_sc_hd__buf_6 fanout819 (.A(net823),
    .X(net819));
 sky130_fd_sc_hd__buf_4 fanout820 (.A(net821),
    .X(net820));
 sky130_fd_sc_hd__buf_4 fanout821 (.A(net823),
    .X(net821));
 sky130_fd_sc_hd__buf_4 fanout822 (.A(net823),
    .X(net822));
 sky130_fd_sc_hd__buf_6 fanout823 (.A(\sel_1$5738 ),
    .X(net823));
 sky130_fd_sc_hd__buf_4 fanout824 (.A(net826),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_4 fanout825 (.A(net826),
    .X(net825));
 sky130_fd_sc_hd__buf_4 fanout826 (.A(net832),
    .X(net826));
 sky130_fd_sc_hd__buf_4 fanout827 (.A(net832),
    .X(net827));
 sky130_fd_sc_hd__buf_4 fanout828 (.A(net829),
    .X(net828));
 sky130_fd_sc_hd__buf_6 fanout829 (.A(net831),
    .X(net829));
 sky130_fd_sc_hd__buf_4 fanout830 (.A(net831),
    .X(net830));
 sky130_fd_sc_hd__buf_4 fanout831 (.A(net832),
    .X(net831));
 sky130_fd_sc_hd__buf_4 fanout832 (.A(\sel_1$5668 ),
    .X(net832));
 sky130_fd_sc_hd__buf_4 fanout833 (.A(net835),
    .X(net833));
 sky130_fd_sc_hd__clkbuf_2 fanout834 (.A(net835),
    .X(net834));
 sky130_fd_sc_hd__buf_4 fanout835 (.A(net841),
    .X(net835));
 sky130_fd_sc_hd__buf_4 fanout836 (.A(net837),
    .X(net836));
 sky130_fd_sc_hd__buf_4 fanout837 (.A(net841),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_8 fanout838 (.A(net841),
    .X(net838));
 sky130_fd_sc_hd__buf_4 fanout839 (.A(net841),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_8 fanout840 (.A(net841),
    .X(net840));
 sky130_fd_sc_hd__buf_8 fanout841 (.A(\sel_1$5598 ),
    .X(net841));
 sky130_fd_sc_hd__buf_6 fanout842 (.A(net843),
    .X(net842));
 sky130_fd_sc_hd__buf_8 fanout843 (.A(\sel_1$5528 ),
    .X(net843));
 sky130_fd_sc_hd__buf_4 fanout844 (.A(net845),
    .X(net844));
 sky130_fd_sc_hd__buf_6 fanout845 (.A(\sel_1$5528 ),
    .X(net845));
 sky130_fd_sc_hd__buf_4 fanout846 (.A(net847),
    .X(net846));
 sky130_fd_sc_hd__buf_4 fanout847 (.A(net848),
    .X(net847));
 sky130_fd_sc_hd__buf_6 fanout848 (.A(\sel_1$5528 ),
    .X(net848));
 sky130_fd_sc_hd__buf_4 fanout849 (.A(net856),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_4 fanout850 (.A(net856),
    .X(net850));
 sky130_fd_sc_hd__buf_4 fanout851 (.A(net852),
    .X(net851));
 sky130_fd_sc_hd__buf_6 fanout852 (.A(net856),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_4 fanout853 (.A(net854),
    .X(net853));
 sky130_fd_sc_hd__buf_6 fanout854 (.A(net855),
    .X(net854));
 sky130_fd_sc_hd__buf_6 fanout855 (.A(net856),
    .X(net855));
 sky130_fd_sc_hd__buf_6 fanout856 (.A(\sel_1$5458 ),
    .X(net856));
 sky130_fd_sc_hd__buf_4 fanout857 (.A(net859),
    .X(net857));
 sky130_fd_sc_hd__clkbuf_4 fanout858 (.A(net859),
    .X(net858));
 sky130_fd_sc_hd__buf_4 fanout859 (.A(net865),
    .X(net859));
 sky130_fd_sc_hd__buf_4 fanout860 (.A(net861),
    .X(net860));
 sky130_fd_sc_hd__buf_6 fanout861 (.A(net865),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_8 fanout862 (.A(net865),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_4 fanout863 (.A(net865),
    .X(net863));
 sky130_fd_sc_hd__buf_4 fanout864 (.A(net865),
    .X(net864));
 sky130_fd_sc_hd__buf_6 fanout865 (.A(\sel_1$5388 ),
    .X(net865));
 sky130_fd_sc_hd__buf_4 fanout866 (.A(net868),
    .X(net866));
 sky130_fd_sc_hd__clkbuf_2 fanout867 (.A(net868),
    .X(net867));
 sky130_fd_sc_hd__buf_2 fanout868 (.A(net874),
    .X(net868));
 sky130_fd_sc_hd__buf_4 fanout869 (.A(net870),
    .X(net869));
 sky130_fd_sc_hd__buf_6 fanout870 (.A(net874),
    .X(net870));
 sky130_fd_sc_hd__buf_4 fanout871 (.A(net873),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_4 fanout872 (.A(net873),
    .X(net872));
 sky130_fd_sc_hd__buf_6 fanout873 (.A(net874),
    .X(net873));
 sky130_fd_sc_hd__buf_6 fanout874 (.A(\sel_1$5318 ),
    .X(net874));
 sky130_fd_sc_hd__buf_4 fanout875 (.A(net877),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_4 fanout876 (.A(net877),
    .X(net876));
 sky130_fd_sc_hd__buf_4 fanout877 (.A(\sel_1$5248 ),
    .X(net877));
 sky130_fd_sc_hd__buf_4 fanout878 (.A(net879),
    .X(net878));
 sky130_fd_sc_hd__buf_6 fanout879 (.A(\sel_1$5248 ),
    .X(net879));
 sky130_fd_sc_hd__buf_6 fanout880 (.A(net882),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_4 fanout881 (.A(net882),
    .X(net881));
 sky130_fd_sc_hd__buf_6 fanout882 (.A(\sel_1$5248 ),
    .X(net882));
 sky130_fd_sc_hd__buf_4 fanout883 (.A(net885),
    .X(net883));
 sky130_fd_sc_hd__buf_2 fanout884 (.A(net885),
    .X(net884));
 sky130_fd_sc_hd__buf_6 fanout885 (.A(\sel_1$5178 ),
    .X(net885));
 sky130_fd_sc_hd__buf_4 fanout886 (.A(net888),
    .X(net886));
 sky130_fd_sc_hd__buf_2 fanout887 (.A(net888),
    .X(net887));
 sky130_fd_sc_hd__buf_4 fanout888 (.A(\sel_1$5178 ),
    .X(net888));
 sky130_fd_sc_hd__buf_4 fanout889 (.A(net891),
    .X(net889));
 sky130_fd_sc_hd__clkbuf_4 fanout890 (.A(net891),
    .X(net890));
 sky130_fd_sc_hd__buf_6 fanout891 (.A(\sel_1$5178 ),
    .X(net891));
 sky130_fd_sc_hd__buf_4 fanout892 (.A(net895),
    .X(net892));
 sky130_fd_sc_hd__clkbuf_4 fanout893 (.A(net895),
    .X(net893));
 sky130_fd_sc_hd__buf_4 fanout894 (.A(net895),
    .X(net894));
 sky130_fd_sc_hd__clkbuf_8 fanout895 (.A(\sel_1$4478 ),
    .X(net895));
 sky130_fd_sc_hd__clkbuf_4 fanout896 (.A(net898),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_4 fanout897 (.A(net898),
    .X(net897));
 sky130_fd_sc_hd__clkbuf_4 fanout898 (.A(\sel_1$4478 ),
    .X(net898));
 sky130_fd_sc_hd__buf_4 fanout899 (.A(\sel_1$4478 ),
    .X(net899));
 sky130_fd_sc_hd__buf_4 fanout900 (.A(net901),
    .X(net900));
 sky130_fd_sc_hd__buf_6 fanout901 (.A(net904),
    .X(net901));
 sky130_fd_sc_hd__clkbuf_8 fanout902 (.A(net903),
    .X(net902));
 sky130_fd_sc_hd__buf_6 fanout903 (.A(net904),
    .X(net903));
 sky130_fd_sc_hd__buf_4 fanout904 (.A(\sel_1$5108 ),
    .X(net904));
 sky130_fd_sc_hd__buf_4 fanout905 (.A(net907),
    .X(net905));
 sky130_fd_sc_hd__clkbuf_4 fanout906 (.A(net907),
    .X(net906));
 sky130_fd_sc_hd__buf_6 fanout907 (.A(\sel_1$5108 ),
    .X(net907));
 sky130_fd_sc_hd__buf_4 fanout908 (.A(net909),
    .X(net908));
 sky130_fd_sc_hd__buf_6 fanout909 (.A(net912),
    .X(net909));
 sky130_fd_sc_hd__buf_4 fanout910 (.A(net911),
    .X(net910));
 sky130_fd_sc_hd__buf_6 fanout911 (.A(net912),
    .X(net911));
 sky130_fd_sc_hd__buf_6 fanout912 (.A(\sel_1$5038 ),
    .X(net912));
 sky130_fd_sc_hd__buf_4 fanout913 (.A(net915),
    .X(net913));
 sky130_fd_sc_hd__clkbuf_4 fanout914 (.A(net915),
    .X(net914));
 sky130_fd_sc_hd__buf_6 fanout915 (.A(\sel_1$5038 ),
    .X(net915));
 sky130_fd_sc_hd__buf_4 fanout916 (.A(net917),
    .X(net916));
 sky130_fd_sc_hd__buf_6 fanout917 (.A(net920),
    .X(net917));
 sky130_fd_sc_hd__clkbuf_8 fanout918 (.A(net919),
    .X(net918));
 sky130_fd_sc_hd__buf_6 fanout919 (.A(net920),
    .X(net919));
 sky130_fd_sc_hd__buf_4 fanout920 (.A(\sel_1$4968 ),
    .X(net920));
 sky130_fd_sc_hd__buf_6 fanout921 (.A(net923),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_4 fanout922 (.A(net923),
    .X(net922));
 sky130_fd_sc_hd__buf_6 fanout923 (.A(\sel_1$4968 ),
    .X(net923));
 sky130_fd_sc_hd__buf_4 fanout924 (.A(net925),
    .X(net924));
 sky130_fd_sc_hd__buf_6 fanout925 (.A(net931),
    .X(net925));
 sky130_fd_sc_hd__clkbuf_8 fanout926 (.A(net931),
    .X(net926));
 sky130_fd_sc_hd__buf_4 fanout927 (.A(net931),
    .X(net927));
 sky130_fd_sc_hd__buf_6 fanout928 (.A(net931),
    .X(net928));
 sky130_fd_sc_hd__clkbuf_8 fanout929 (.A(net930),
    .X(net929));
 sky130_fd_sc_hd__buf_4 fanout930 (.A(net931),
    .X(net930));
 sky130_fd_sc_hd__buf_12 fanout931 (.A(net99),
    .X(net931));
 sky130_fd_sc_hd__clkbuf_4 fanout932 (.A(net934),
    .X(net932));
 sky130_fd_sc_hd__buf_4 fanout933 (.A(net934),
    .X(net933));
 sky130_fd_sc_hd__clkbuf_4 fanout934 (.A(net935),
    .X(net934));
 sky130_fd_sc_hd__buf_6 fanout935 (.A(net98),
    .X(net935));
 sky130_fd_sc_hd__buf_4 fanout936 (.A(net939),
    .X(net936));
 sky130_fd_sc_hd__clkbuf_4 fanout937 (.A(net939),
    .X(net937));
 sky130_fd_sc_hd__buf_4 fanout938 (.A(net939),
    .X(net938));
 sky130_fd_sc_hd__clkbuf_8 fanout939 (.A(net98),
    .X(net939));
 sky130_fd_sc_hd__buf_4 fanout940 (.A(net941),
    .X(net940));
 sky130_fd_sc_hd__buf_6 fanout941 (.A(net947),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_8 fanout942 (.A(net947),
    .X(net942));
 sky130_fd_sc_hd__buf_4 fanout943 (.A(net947),
    .X(net943));
 sky130_fd_sc_hd__buf_4 fanout944 (.A(net947),
    .X(net944));
 sky130_fd_sc_hd__buf_4 fanout945 (.A(net946),
    .X(net945));
 sky130_fd_sc_hd__buf_4 fanout946 (.A(net947),
    .X(net946));
 sky130_fd_sc_hd__buf_12 fanout947 (.A(net97),
    .X(net947));
 sky130_fd_sc_hd__buf_4 fanout948 (.A(net949),
    .X(net948));
 sky130_fd_sc_hd__buf_6 fanout949 (.A(net952),
    .X(net949));
 sky130_fd_sc_hd__buf_6 fanout950 (.A(net952),
    .X(net950));
 sky130_fd_sc_hd__buf_4 fanout951 (.A(net952),
    .X(net951));
 sky130_fd_sc_hd__buf_6 fanout952 (.A(net96),
    .X(net952));
 sky130_fd_sc_hd__buf_6 fanout953 (.A(net954),
    .X(net953));
 sky130_fd_sc_hd__buf_4 fanout954 (.A(net96),
    .X(net954));
 sky130_fd_sc_hd__buf_4 fanout955 (.A(net96),
    .X(net955));
 sky130_fd_sc_hd__buf_4 fanout956 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__buf_6 fanout957 (.A(net960),
    .X(net957));
 sky130_fd_sc_hd__buf_6 fanout958 (.A(net959),
    .X(net958));
 sky130_fd_sc_hd__buf_6 fanout959 (.A(net960),
    .X(net959));
 sky130_fd_sc_hd__buf_4 fanout960 (.A(net95),
    .X(net960));
 sky130_fd_sc_hd__buf_4 fanout961 (.A(net963),
    .X(net961));
 sky130_fd_sc_hd__buf_6 fanout962 (.A(net963),
    .X(net962));
 sky130_fd_sc_hd__buf_4 fanout963 (.A(net95),
    .X(net963));
 sky130_fd_sc_hd__buf_4 fanout964 (.A(net965),
    .X(net964));
 sky130_fd_sc_hd__buf_6 fanout965 (.A(net968),
    .X(net965));
 sky130_fd_sc_hd__buf_4 fanout966 (.A(net968),
    .X(net966));
 sky130_fd_sc_hd__buf_4 fanout967 (.A(net968),
    .X(net967));
 sky130_fd_sc_hd__buf_6 fanout968 (.A(net94),
    .X(net968));
 sky130_fd_sc_hd__buf_4 fanout969 (.A(net972),
    .X(net969));
 sky130_fd_sc_hd__buf_6 fanout970 (.A(net972),
    .X(net970));
 sky130_fd_sc_hd__buf_2 fanout971 (.A(net972),
    .X(net971));
 sky130_fd_sc_hd__buf_6 fanout972 (.A(net94),
    .X(net972));
 sky130_fd_sc_hd__buf_4 fanout973 (.A(net974),
    .X(net973));
 sky130_fd_sc_hd__buf_6 fanout974 (.A(net981),
    .X(net974));
 sky130_fd_sc_hd__buf_4 fanout975 (.A(net981),
    .X(net975));
 sky130_fd_sc_hd__buf_4 fanout976 (.A(net981),
    .X(net976));
 sky130_fd_sc_hd__buf_6 fanout977 (.A(net980),
    .X(net977));
 sky130_fd_sc_hd__buf_2 fanout978 (.A(net980),
    .X(net978));
 sky130_fd_sc_hd__buf_6 fanout979 (.A(net980),
    .X(net979));
 sky130_fd_sc_hd__buf_4 fanout980 (.A(net981),
    .X(net980));
 sky130_fd_sc_hd__buf_8 fanout981 (.A(net93),
    .X(net981));
 sky130_fd_sc_hd__buf_4 fanout982 (.A(net983),
    .X(net982));
 sky130_fd_sc_hd__buf_6 fanout983 (.A(net986),
    .X(net983));
 sky130_fd_sc_hd__buf_4 fanout984 (.A(net986),
    .X(net984));
 sky130_fd_sc_hd__buf_4 fanout985 (.A(net986),
    .X(net985));
 sky130_fd_sc_hd__buf_6 fanout986 (.A(net92),
    .X(net986));
 sky130_fd_sc_hd__buf_4 fanout987 (.A(net989),
    .X(net987));
 sky130_fd_sc_hd__buf_6 fanout988 (.A(net989),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_8 fanout989 (.A(net92),
    .X(net989));
 sky130_fd_sc_hd__buf_4 fanout990 (.A(net991),
    .X(net990));
 sky130_fd_sc_hd__buf_6 fanout991 (.A(net91),
    .X(net991));
 sky130_fd_sc_hd__buf_4 fanout992 (.A(net993),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_4 fanout993 (.A(net91),
    .X(net993));
 sky130_fd_sc_hd__buf_6 fanout994 (.A(net997),
    .X(net994));
 sky130_fd_sc_hd__buf_4 fanout995 (.A(net997),
    .X(net995));
 sky130_fd_sc_hd__buf_4 fanout996 (.A(net997),
    .X(net996));
 sky130_fd_sc_hd__clkbuf_8 fanout997 (.A(net91),
    .X(net997));
 sky130_fd_sc_hd__buf_4 fanout998 (.A(net999),
    .X(net998));
 sky130_fd_sc_hd__buf_6 fanout999 (.A(net1005),
    .X(net999));
 sky130_fd_sc_hd__buf_4 fanout1000 (.A(net1001),
    .X(net1000));
 sky130_fd_sc_hd__buf_4 fanout1001 (.A(net1005),
    .X(net1001));
 sky130_fd_sc_hd__buf_6 fanout1002 (.A(net1004),
    .X(net1002));
 sky130_fd_sc_hd__buf_4 fanout1003 (.A(net1004),
    .X(net1003));
 sky130_fd_sc_hd__buf_6 fanout1004 (.A(net1005),
    .X(net1004));
 sky130_fd_sc_hd__buf_6 fanout1005 (.A(net90),
    .X(net1005));
 sky130_fd_sc_hd__buf_6 fanout1006 (.A(net1008),
    .X(net1006));
 sky130_fd_sc_hd__buf_6 fanout1007 (.A(net1008),
    .X(net1007));
 sky130_fd_sc_hd__buf_6 fanout1008 (.A(net1011),
    .X(net1008));
 sky130_fd_sc_hd__buf_6 fanout1009 (.A(net1010),
    .X(net1009));
 sky130_fd_sc_hd__buf_6 fanout1010 (.A(net1011),
    .X(net1010));
 sky130_fd_sc_hd__buf_6 fanout1011 (.A(net9),
    .X(net1011));
 sky130_fd_sc_hd__buf_6 fanout1012 (.A(net1014),
    .X(net1012));
 sky130_fd_sc_hd__buf_4 fanout1013 (.A(net1014),
    .X(net1013));
 sky130_fd_sc_hd__buf_6 fanout1014 (.A(net9),
    .X(net1014));
 sky130_fd_sc_hd__buf_4 fanout1015 (.A(net1016),
    .X(net1015));
 sky130_fd_sc_hd__buf_6 fanout1016 (.A(net1022),
    .X(net1016));
 sky130_fd_sc_hd__buf_4 fanout1017 (.A(net1018),
    .X(net1017));
 sky130_fd_sc_hd__buf_6 fanout1018 (.A(net1022),
    .X(net1018));
 sky130_fd_sc_hd__buf_6 fanout1019 (.A(net1021),
    .X(net1019));
 sky130_fd_sc_hd__buf_4 fanout1020 (.A(net1021),
    .X(net1020));
 sky130_fd_sc_hd__buf_6 fanout1021 (.A(net1022),
    .X(net1021));
 sky130_fd_sc_hd__buf_8 fanout1022 (.A(net89),
    .X(net1022));
 sky130_fd_sc_hd__buf_4 fanout1023 (.A(net1024),
    .X(net1023));
 sky130_fd_sc_hd__buf_6 fanout1024 (.A(net1030),
    .X(net1024));
 sky130_fd_sc_hd__buf_4 fanout1025 (.A(net1026),
    .X(net1025));
 sky130_fd_sc_hd__buf_6 fanout1026 (.A(net1030),
    .X(net1026));
 sky130_fd_sc_hd__buf_4 fanout1027 (.A(net1029),
    .X(net1027));
 sky130_fd_sc_hd__buf_4 fanout1028 (.A(net1029),
    .X(net1028));
 sky130_fd_sc_hd__buf_6 fanout1029 (.A(net1030),
    .X(net1029));
 sky130_fd_sc_hd__buf_6 fanout1030 (.A(net88),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_4 fanout1031 (.A(net1033),
    .X(net1031));
 sky130_fd_sc_hd__buf_4 fanout1032 (.A(net1033),
    .X(net1032));
 sky130_fd_sc_hd__buf_2 fanout1033 (.A(net1034),
    .X(net1033));
 sky130_fd_sc_hd__buf_6 fanout1034 (.A(net87),
    .X(net1034));
 sky130_fd_sc_hd__clkbuf_4 fanout1035 (.A(net1038),
    .X(net1035));
 sky130_fd_sc_hd__buf_4 fanout1036 (.A(net1038),
    .X(net1036));
 sky130_fd_sc_hd__buf_4 fanout1037 (.A(net1038),
    .X(net1037));
 sky130_fd_sc_hd__buf_4 fanout1038 (.A(net87),
    .X(net1038));
 sky130_fd_sc_hd__clkbuf_8 fanout1039 (.A(net1040),
    .X(net1039));
 sky130_fd_sc_hd__buf_6 fanout1040 (.A(net1046),
    .X(net1040));
 sky130_fd_sc_hd__buf_4 fanout1041 (.A(net1042),
    .X(net1041));
 sky130_fd_sc_hd__buf_6 fanout1042 (.A(net1046),
    .X(net1042));
 sky130_fd_sc_hd__buf_4 fanout1043 (.A(net1045),
    .X(net1043));
 sky130_fd_sc_hd__buf_2 fanout1044 (.A(net1045),
    .X(net1044));
 sky130_fd_sc_hd__buf_6 fanout1045 (.A(net1046),
    .X(net1045));
 sky130_fd_sc_hd__buf_6 fanout1046 (.A(net86),
    .X(net1046));
 sky130_fd_sc_hd__clkbuf_8 fanout1047 (.A(net1048),
    .X(net1047));
 sky130_fd_sc_hd__buf_6 fanout1048 (.A(net1054),
    .X(net1048));
 sky130_fd_sc_hd__buf_4 fanout1049 (.A(net1050),
    .X(net1049));
 sky130_fd_sc_hd__buf_6 fanout1050 (.A(net1054),
    .X(net1050));
 sky130_fd_sc_hd__buf_4 fanout1051 (.A(net1053),
    .X(net1051));
 sky130_fd_sc_hd__buf_2 fanout1052 (.A(net1053),
    .X(net1052));
 sky130_fd_sc_hd__buf_6 fanout1053 (.A(net1054),
    .X(net1053));
 sky130_fd_sc_hd__buf_6 fanout1054 (.A(net85),
    .X(net1054));
 sky130_fd_sc_hd__buf_4 fanout1055 (.A(net1056),
    .X(net1055));
 sky130_fd_sc_hd__buf_6 fanout1056 (.A(net1059),
    .X(net1056));
 sky130_fd_sc_hd__buf_4 fanout1057 (.A(net1058),
    .X(net1057));
 sky130_fd_sc_hd__buf_6 fanout1058 (.A(net1059),
    .X(net1058));
 sky130_fd_sc_hd__buf_4 fanout1059 (.A(net84),
    .X(net1059));
 sky130_fd_sc_hd__buf_4 fanout1060 (.A(net1062),
    .X(net1060));
 sky130_fd_sc_hd__buf_2 fanout1061 (.A(net1062),
    .X(net1061));
 sky130_fd_sc_hd__buf_6 fanout1062 (.A(net84),
    .X(net1062));
 sky130_fd_sc_hd__buf_4 fanout1063 (.A(net1064),
    .X(net1063));
 sky130_fd_sc_hd__buf_4 fanout1064 (.A(net83),
    .X(net1064));
 sky130_fd_sc_hd__buf_2 fanout1065 (.A(net83),
    .X(net1065));
 sky130_fd_sc_hd__buf_4 fanout1066 (.A(net1067),
    .X(net1066));
 sky130_fd_sc_hd__buf_4 fanout1067 (.A(net83),
    .X(net1067));
 sky130_fd_sc_hd__clkbuf_8 fanout1068 (.A(net1070),
    .X(net1068));
 sky130_fd_sc_hd__clkbuf_4 fanout1069 (.A(net1070),
    .X(net1069));
 sky130_fd_sc_hd__buf_6 fanout1070 (.A(net83),
    .X(net1070));
 sky130_fd_sc_hd__buf_4 fanout1071 (.A(net1072),
    .X(net1071));
 sky130_fd_sc_hd__clkbuf_4 fanout1072 (.A(net1079),
    .X(net1072));
 sky130_fd_sc_hd__buf_4 fanout1073 (.A(net1079),
    .X(net1073));
 sky130_fd_sc_hd__buf_4 fanout1074 (.A(net1075),
    .X(net1074));
 sky130_fd_sc_hd__buf_4 fanout1075 (.A(net1079),
    .X(net1075));
 sky130_fd_sc_hd__buf_4 fanout1076 (.A(net1078),
    .X(net1076));
 sky130_fd_sc_hd__clkbuf_4 fanout1077 (.A(net1078),
    .X(net1077));
 sky130_fd_sc_hd__buf_6 fanout1078 (.A(net1079),
    .X(net1078));
 sky130_fd_sc_hd__buf_4 fanout1079 (.A(net82),
    .X(net1079));
 sky130_fd_sc_hd__buf_4 fanout1080 (.A(net1081),
    .X(net1080));
 sky130_fd_sc_hd__buf_4 fanout1081 (.A(net1082),
    .X(net1081));
 sky130_fd_sc_hd__buf_6 fanout1082 (.A(net81),
    .X(net1082));
 sky130_fd_sc_hd__buf_4 fanout1083 (.A(net1084),
    .X(net1083));
 sky130_fd_sc_hd__clkbuf_8 fanout1084 (.A(net81),
    .X(net1084));
 sky130_fd_sc_hd__buf_4 fanout1085 (.A(net1086),
    .X(net1085));
 sky130_fd_sc_hd__buf_4 fanout1086 (.A(net1087),
    .X(net1086));
 sky130_fd_sc_hd__buf_4 fanout1087 (.A(net81),
    .X(net1087));
 sky130_fd_sc_hd__buf_4 fanout1088 (.A(net1093),
    .X(net1088));
 sky130_fd_sc_hd__buf_2 fanout1089 (.A(net1093),
    .X(net1089));
 sky130_fd_sc_hd__buf_6 fanout1090 (.A(net1093),
    .X(net1090));
 sky130_fd_sc_hd__clkbuf_8 fanout1091 (.A(net1092),
    .X(net1091));
 sky130_fd_sc_hd__clkbuf_8 fanout1092 (.A(net1093),
    .X(net1092));
 sky130_fd_sc_hd__buf_4 fanout1093 (.A(net80),
    .X(net1093));
 sky130_fd_sc_hd__clkbuf_8 fanout1094 (.A(net1096),
    .X(net1094));
 sky130_fd_sc_hd__buf_4 fanout1095 (.A(net1096),
    .X(net1095));
 sky130_fd_sc_hd__clkbuf_8 fanout1096 (.A(net80),
    .X(net1096));
 sky130_fd_sc_hd__buf_4 fanout1097 (.A(net1099),
    .X(net1097));
 sky130_fd_sc_hd__clkbuf_8 fanout1098 (.A(net1099),
    .X(net1098));
 sky130_fd_sc_hd__buf_4 fanout1099 (.A(net79),
    .X(net1099));
 sky130_fd_sc_hd__clkbuf_8 fanout1100 (.A(net1101),
    .X(net1100));
 sky130_fd_sc_hd__buf_6 fanout1101 (.A(net79),
    .X(net1101));
 sky130_fd_sc_hd__clkbuf_8 fanout1102 (.A(net1104),
    .X(net1102));
 sky130_fd_sc_hd__buf_4 fanout1103 (.A(net1104),
    .X(net1103));
 sky130_fd_sc_hd__buf_4 fanout1104 (.A(net79),
    .X(net1104));
 sky130_fd_sc_hd__buf_4 fanout1105 (.A(net1110),
    .X(net1105));
 sky130_fd_sc_hd__clkbuf_4 fanout1106 (.A(net1110),
    .X(net1106));
 sky130_fd_sc_hd__clkbuf_8 fanout1107 (.A(net1110),
    .X(net1107));
 sky130_fd_sc_hd__buf_4 fanout1108 (.A(net1110),
    .X(net1108));
 sky130_fd_sc_hd__buf_4 fanout1109 (.A(net1110),
    .X(net1109));
 sky130_fd_sc_hd__buf_6 fanout1110 (.A(net78),
    .X(net1110));
 sky130_fd_sc_hd__buf_4 fanout1111 (.A(net1113),
    .X(net1111));
 sky130_fd_sc_hd__buf_4 fanout1112 (.A(net1113),
    .X(net1112));
 sky130_fd_sc_hd__buf_4 fanout1113 (.A(net78),
    .X(net1113));
 sky130_fd_sc_hd__buf_4 fanout1114 (.A(net1116),
    .X(net1114));
 sky130_fd_sc_hd__buf_2 fanout1115 (.A(net1116),
    .X(net1115));
 sky130_fd_sc_hd__buf_6 fanout1116 (.A(net77),
    .X(net1116));
 sky130_fd_sc_hd__buf_4 fanout1117 (.A(net1118),
    .X(net1117));
 sky130_fd_sc_hd__buf_4 fanout1118 (.A(net77),
    .X(net1118));
 sky130_fd_sc_hd__buf_6 fanout1119 (.A(net1120),
    .X(net1119));
 sky130_fd_sc_hd__buf_6 fanout1120 (.A(net1121),
    .X(net1120));
 sky130_fd_sc_hd__buf_4 fanout1121 (.A(net77),
    .X(net1121));
 sky130_fd_sc_hd__buf_4 fanout1122 (.A(net1124),
    .X(net1122));
 sky130_fd_sc_hd__buf_4 fanout1123 (.A(net1124),
    .X(net1123));
 sky130_fd_sc_hd__buf_2 fanout1124 (.A(net1125),
    .X(net1124));
 sky130_fd_sc_hd__buf_4 fanout1125 (.A(net76),
    .X(net1125));
 sky130_fd_sc_hd__buf_4 fanout1126 (.A(net1128),
    .X(net1126));
 sky130_fd_sc_hd__clkbuf_4 fanout1127 (.A(net1128),
    .X(net1127));
 sky130_fd_sc_hd__clkbuf_4 fanout1128 (.A(net76),
    .X(net1128));
 sky130_fd_sc_hd__buf_4 fanout1129 (.A(net76),
    .X(net1129));
 sky130_fd_sc_hd__buf_4 fanout1130 (.A(net1132),
    .X(net1130));
 sky130_fd_sc_hd__buf_2 fanout1131 (.A(net1132),
    .X(net1131));
 sky130_fd_sc_hd__buf_6 fanout1132 (.A(net75),
    .X(net1132));
 sky130_fd_sc_hd__buf_4 fanout1133 (.A(net1134),
    .X(net1133));
 sky130_fd_sc_hd__buf_4 fanout1134 (.A(net75),
    .X(net1134));
 sky130_fd_sc_hd__buf_6 fanout1135 (.A(net1136),
    .X(net1135));
 sky130_fd_sc_hd__buf_6 fanout1136 (.A(net1137),
    .X(net1136));
 sky130_fd_sc_hd__clkbuf_8 fanout1137 (.A(net75),
    .X(net1137));
 sky130_fd_sc_hd__buf_4 fanout1138 (.A(net1140),
    .X(net1138));
 sky130_fd_sc_hd__buf_4 fanout1139 (.A(net1140),
    .X(net1139));
 sky130_fd_sc_hd__clkbuf_4 fanout1140 (.A(net74),
    .X(net1140));
 sky130_fd_sc_hd__buf_4 fanout1141 (.A(net74),
    .X(net1141));
 sky130_fd_sc_hd__clkbuf_4 fanout1142 (.A(net74),
    .X(net1142));
 sky130_fd_sc_hd__buf_4 fanout1143 (.A(net1145),
    .X(net1143));
 sky130_fd_sc_hd__clkbuf_4 fanout1144 (.A(net1145),
    .X(net1144));
 sky130_fd_sc_hd__buf_4 fanout1145 (.A(net74),
    .X(net1145));
 sky130_fd_sc_hd__buf_4 fanout1146 (.A(net1147),
    .X(net1146));
 sky130_fd_sc_hd__buf_4 fanout1147 (.A(net1154),
    .X(net1147));
 sky130_fd_sc_hd__clkbuf_4 fanout1148 (.A(net1154),
    .X(net1148));
 sky130_fd_sc_hd__clkbuf_8 fanout1149 (.A(net1154),
    .X(net1149));
 sky130_fd_sc_hd__buf_4 fanout1150 (.A(net1154),
    .X(net1150));
 sky130_fd_sc_hd__buf_4 fanout1151 (.A(net1153),
    .X(net1151));
 sky130_fd_sc_hd__buf_4 fanout1152 (.A(net1153),
    .X(net1152));
 sky130_fd_sc_hd__clkbuf_8 fanout1153 (.A(net1154),
    .X(net1153));
 sky130_fd_sc_hd__buf_4 fanout1154 (.A(net73),
    .X(net1154));
 sky130_fd_sc_hd__buf_4 fanout1155 (.A(net1158),
    .X(net1155));
 sky130_fd_sc_hd__buf_2 fanout1156 (.A(net1158),
    .X(net1156));
 sky130_fd_sc_hd__buf_4 fanout1157 (.A(net1158),
    .X(net1157));
 sky130_fd_sc_hd__buf_4 fanout1158 (.A(net72),
    .X(net1158));
 sky130_fd_sc_hd__buf_6 fanout1159 (.A(net72),
    .X(net1159));
 sky130_fd_sc_hd__buf_2 fanout1160 (.A(net72),
    .X(net1160));
 sky130_fd_sc_hd__clkbuf_8 fanout1161 (.A(net1163),
    .X(net1161));
 sky130_fd_sc_hd__clkbuf_2 fanout1162 (.A(net1163),
    .X(net1162));
 sky130_fd_sc_hd__buf_4 fanout1163 (.A(net72),
    .X(net1163));
 sky130_fd_sc_hd__buf_4 fanout1164 (.A(net1167),
    .X(net1164));
 sky130_fd_sc_hd__buf_2 fanout1165 (.A(net1167),
    .X(net1165));
 sky130_fd_sc_hd__buf_4 fanout1166 (.A(net1167),
    .X(net1166));
 sky130_fd_sc_hd__buf_4 fanout1167 (.A(net71),
    .X(net1167));
 sky130_fd_sc_hd__clkbuf_8 fanout1168 (.A(net71),
    .X(net1168));
 sky130_fd_sc_hd__clkbuf_2 fanout1169 (.A(net71),
    .X(net1169));
 sky130_fd_sc_hd__buf_6 fanout1170 (.A(net1172),
    .X(net1170));
 sky130_fd_sc_hd__clkbuf_4 fanout1171 (.A(net1172),
    .X(net1171));
 sky130_fd_sc_hd__clkbuf_8 fanout1172 (.A(net71),
    .X(net1172));
 sky130_fd_sc_hd__buf_4 fanout1173 (.A(net1174),
    .X(net1173));
 sky130_fd_sc_hd__clkbuf_4 fanout1174 (.A(net1176),
    .X(net1174));
 sky130_fd_sc_hd__buf_4 fanout1175 (.A(net1176),
    .X(net1175));
 sky130_fd_sc_hd__clkbuf_4 fanout1176 (.A(net1182),
    .X(net1176));
 sky130_fd_sc_hd__buf_4 fanout1177 (.A(net1182),
    .X(net1177));
 sky130_fd_sc_hd__clkbuf_4 fanout1178 (.A(net1182),
    .X(net1178));
 sky130_fd_sc_hd__buf_6 fanout1179 (.A(net1181),
    .X(net1179));
 sky130_fd_sc_hd__clkbuf_4 fanout1180 (.A(net1181),
    .X(net1180));
 sky130_fd_sc_hd__buf_4 fanout1181 (.A(net1182),
    .X(net1181));
 sky130_fd_sc_hd__clkbuf_8 fanout1182 (.A(net70),
    .X(net1182));
 sky130_fd_sc_hd__buf_6 fanout1183 (.A(net1184),
    .X(net1183));
 sky130_fd_sc_hd__buf_8 fanout1184 (.A(net7),
    .X(net1184));
 sky130_fd_sc_hd__buf_6 fanout1185 (.A(net1187),
    .X(net1185));
 sky130_fd_sc_hd__clkbuf_8 fanout1186 (.A(net1187),
    .X(net1186));
 sky130_fd_sc_hd__buf_6 fanout1187 (.A(net7),
    .X(net1187));
 sky130_fd_sc_hd__buf_6 fanout1188 (.A(net1189),
    .X(net1188));
 sky130_fd_sc_hd__clkbuf_4 fanout1189 (.A(net1190),
    .X(net1189));
 sky130_fd_sc_hd__buf_4 fanout1190 (.A(net1191),
    .X(net1190));
 sky130_fd_sc_hd__buf_6 fanout1191 (.A(net7),
    .X(net1191));
 sky130_fd_sc_hd__buf_4 fanout1192 (.A(net1193),
    .X(net1192));
 sky130_fd_sc_hd__buf_4 fanout1193 (.A(net1195),
    .X(net1193));
 sky130_fd_sc_hd__buf_4 fanout1194 (.A(net1195),
    .X(net1194));
 sky130_fd_sc_hd__clkbuf_4 fanout1195 (.A(net1197),
    .X(net1195));
 sky130_fd_sc_hd__clkbuf_8 fanout1196 (.A(net1197),
    .X(net1196));
 sky130_fd_sc_hd__clkbuf_4 fanout1197 (.A(net69),
    .X(net1197));
 sky130_fd_sc_hd__buf_6 fanout1198 (.A(net1200),
    .X(net1198));
 sky130_fd_sc_hd__clkbuf_4 fanout1199 (.A(net1200),
    .X(net1199));
 sky130_fd_sc_hd__buf_4 fanout1200 (.A(net69),
    .X(net1200));
 sky130_fd_sc_hd__buf_4 fanout1201 (.A(net1202),
    .X(net1201));
 sky130_fd_sc_hd__buf_4 fanout1202 (.A(net1209),
    .X(net1202));
 sky130_fd_sc_hd__buf_4 fanout1203 (.A(net1204),
    .X(net1203));
 sky130_fd_sc_hd__clkbuf_4 fanout1204 (.A(net1209),
    .X(net1204));
 sky130_fd_sc_hd__buf_6 fanout1205 (.A(net1209),
    .X(net1205));
 sky130_fd_sc_hd__buf_6 fanout1206 (.A(net1208),
    .X(net1206));
 sky130_fd_sc_hd__clkbuf_4 fanout1207 (.A(net1208),
    .X(net1207));
 sky130_fd_sc_hd__buf_4 fanout1208 (.A(net1209),
    .X(net1208));
 sky130_fd_sc_hd__buf_6 fanout1209 (.A(net68),
    .X(net1209));
 sky130_fd_sc_hd__buf_4 fanout1210 (.A(net1213),
    .X(net1210));
 sky130_fd_sc_hd__buf_4 fanout1211 (.A(net1212),
    .X(net1211));
 sky130_fd_sc_hd__clkbuf_4 fanout1212 (.A(net1213),
    .X(net1212));
 sky130_fd_sc_hd__clkbuf_4 fanout1213 (.A(net1215),
    .X(net1213));
 sky130_fd_sc_hd__buf_6 fanout1214 (.A(net1215),
    .X(net1214));
 sky130_fd_sc_hd__clkbuf_4 fanout1215 (.A(net67),
    .X(net1215));
 sky130_fd_sc_hd__clkbuf_8 fanout1216 (.A(net1218),
    .X(net1216));
 sky130_fd_sc_hd__buf_4 fanout1217 (.A(net1218),
    .X(net1217));
 sky130_fd_sc_hd__buf_6 fanout1218 (.A(net67),
    .X(net1218));
 sky130_fd_sc_hd__buf_4 fanout1219 (.A(net1220),
    .X(net1219));
 sky130_fd_sc_hd__buf_4 fanout1220 (.A(net1223),
    .X(net1220));
 sky130_fd_sc_hd__buf_4 fanout1221 (.A(net1223),
    .X(net1221));
 sky130_fd_sc_hd__buf_6 fanout1222 (.A(net1223),
    .X(net1222));
 sky130_fd_sc_hd__clkbuf_8 fanout1223 (.A(net66),
    .X(net1223));
 sky130_fd_sc_hd__buf_4 fanout1224 (.A(net1226),
    .X(net1224));
 sky130_fd_sc_hd__buf_2 fanout1225 (.A(net1226),
    .X(net1225));
 sky130_fd_sc_hd__buf_6 fanout1226 (.A(net66),
    .X(net1226));
 sky130_fd_sc_hd__buf_4 fanout1227 (.A(net1229),
    .X(net1227));
 sky130_fd_sc_hd__buf_4 fanout1228 (.A(net1229),
    .X(net1228));
 sky130_fd_sc_hd__buf_4 fanout1229 (.A(net1234),
    .X(net1229));
 sky130_fd_sc_hd__clkbuf_4 fanout1230 (.A(net1232),
    .X(net1230));
 sky130_fd_sc_hd__clkbuf_4 fanout1231 (.A(net1232),
    .X(net1231));
 sky130_fd_sc_hd__buf_4 fanout1232 (.A(net1234),
    .X(net1232));
 sky130_fd_sc_hd__buf_6 fanout1233 (.A(net1234),
    .X(net1233));
 sky130_fd_sc_hd__clkbuf_8 fanout1234 (.A(net65),
    .X(net1234));
 sky130_fd_sc_hd__buf_6 fanout1235 (.A(net64),
    .X(net1235));
 sky130_fd_sc_hd__clkbuf_8 fanout1236 (.A(net64),
    .X(net1236));
 sky130_fd_sc_hd__buf_6 fanout1237 (.A(net1238),
    .X(net1237));
 sky130_fd_sc_hd__buf_4 fanout1238 (.A(net64),
    .X(net1238));
 sky130_fd_sc_hd__buf_6 fanout1239 (.A(net1243),
    .X(net1239));
 sky130_fd_sc_hd__buf_2 fanout1240 (.A(net1243),
    .X(net1240));
 sky130_fd_sc_hd__buf_8 fanout1241 (.A(net1243),
    .X(net1241));
 sky130_fd_sc_hd__buf_6 fanout1242 (.A(net1243),
    .X(net1242));
 sky130_fd_sc_hd__buf_6 fanout1243 (.A(net64),
    .X(net1243));
 sky130_fd_sc_hd__buf_6 fanout1244 (.A(net1245),
    .X(net1244));
 sky130_fd_sc_hd__buf_6 fanout1245 (.A(net1253),
    .X(net1245));
 sky130_fd_sc_hd__buf_4 fanout1246 (.A(net1247),
    .X(net1246));
 sky130_fd_sc_hd__buf_4 fanout1247 (.A(net1253),
    .X(net1247));
 sky130_fd_sc_hd__buf_4 fanout1248 (.A(net1249),
    .X(net1248));
 sky130_fd_sc_hd__clkbuf_4 fanout1249 (.A(net1252),
    .X(net1249));
 sky130_fd_sc_hd__buf_6 fanout1250 (.A(net1252),
    .X(net1250));
 sky130_fd_sc_hd__buf_6 fanout1251 (.A(net1252),
    .X(net1251));
 sky130_fd_sc_hd__clkbuf_8 fanout1252 (.A(net1253),
    .X(net1252));
 sky130_fd_sc_hd__buf_6 fanout1253 (.A(net62),
    .X(net1253));
 sky130_fd_sc_hd__buf_6 fanout1254 (.A(net1258),
    .X(net1254));
 sky130_fd_sc_hd__clkbuf_8 fanout1255 (.A(net1257),
    .X(net1255));
 sky130_fd_sc_hd__buf_6 fanout1256 (.A(net1257),
    .X(net1256));
 sky130_fd_sc_hd__buf_4 fanout1257 (.A(net1258),
    .X(net1257));
 sky130_fd_sc_hd__buf_4 fanout1258 (.A(net60),
    .X(net1258));
 sky130_fd_sc_hd__buf_6 fanout1259 (.A(net1262),
    .X(net1259));
 sky130_fd_sc_hd__buf_6 fanout1260 (.A(net1261),
    .X(net1260));
 sky130_fd_sc_hd__buf_6 fanout1261 (.A(net1262),
    .X(net1261));
 sky130_fd_sc_hd__buf_6 fanout1262 (.A(net60),
    .X(net1262));
 sky130_fd_sc_hd__buf_6 fanout1263 (.A(net58),
    .X(net1263));
 sky130_fd_sc_hd__clkbuf_4 fanout1264 (.A(net58),
    .X(net1264));
 sky130_fd_sc_hd__buf_4 fanout1265 (.A(net1266),
    .X(net1265));
 sky130_fd_sc_hd__buf_2 fanout1266 (.A(net1267),
    .X(net1266));
 sky130_fd_sc_hd__buf_4 fanout1267 (.A(net1268),
    .X(net1267));
 sky130_fd_sc_hd__buf_4 fanout1268 (.A(net58),
    .X(net1268));
 sky130_fd_sc_hd__buf_6 fanout1269 (.A(net1272),
    .X(net1269));
 sky130_fd_sc_hd__buf_6 fanout1270 (.A(net1271),
    .X(net1270));
 sky130_fd_sc_hd__buf_6 fanout1271 (.A(net1272),
    .X(net1271));
 sky130_fd_sc_hd__buf_4 fanout1272 (.A(net58),
    .X(net1272));
 sky130_fd_sc_hd__buf_6 fanout1273 (.A(net1274),
    .X(net1273));
 sky130_fd_sc_hd__buf_6 fanout1274 (.A(net1276),
    .X(net1274));
 sky130_fd_sc_hd__buf_4 fanout1275 (.A(net1276),
    .X(net1275));
 sky130_fd_sc_hd__buf_8 fanout1276 (.A(net1281),
    .X(net1276));
 sky130_fd_sc_hd__buf_6 fanout1277 (.A(net1278),
    .X(net1277));
 sky130_fd_sc_hd__buf_4 fanout1278 (.A(net1281),
    .X(net1278));
 sky130_fd_sc_hd__buf_6 fanout1279 (.A(net1281),
    .X(net1279));
 sky130_fd_sc_hd__buf_6 fanout1280 (.A(net1281),
    .X(net1280));
 sky130_fd_sc_hd__buf_6 fanout1281 (.A(net56),
    .X(net1281));
 sky130_fd_sc_hd__buf_6 fanout1282 (.A(net55),
    .X(net1282));
 sky130_fd_sc_hd__clkbuf_4 fanout1283 (.A(net55),
    .X(net1283));
 sky130_fd_sc_hd__clkbuf_4 fanout1284 (.A(net1285),
    .X(net1284));
 sky130_fd_sc_hd__buf_4 fanout1285 (.A(net1286),
    .X(net1285));
 sky130_fd_sc_hd__buf_6 fanout1286 (.A(net55),
    .X(net1286));
 sky130_fd_sc_hd__buf_6 fanout1287 (.A(net1290),
    .X(net1287));
 sky130_fd_sc_hd__buf_6 fanout1288 (.A(net1290),
    .X(net1288));
 sky130_fd_sc_hd__buf_6 fanout1289 (.A(net1290),
    .X(net1289));
 sky130_fd_sc_hd__buf_6 fanout1290 (.A(net55),
    .X(net1290));
 sky130_fd_sc_hd__buf_6 fanout1291 (.A(net1295),
    .X(net1291));
 sky130_fd_sc_hd__buf_4 fanout1292 (.A(net1293),
    .X(net1292));
 sky130_fd_sc_hd__buf_6 fanout1293 (.A(net1294),
    .X(net1293));
 sky130_fd_sc_hd__buf_6 fanout1294 (.A(net1295),
    .X(net1294));
 sky130_fd_sc_hd__buf_4 fanout1295 (.A(net53),
    .X(net1295));
 sky130_fd_sc_hd__buf_6 fanout1296 (.A(net1299),
    .X(net1296));
 sky130_fd_sc_hd__buf_6 fanout1297 (.A(net1299),
    .X(net1297));
 sky130_fd_sc_hd__buf_4 fanout1298 (.A(net1299),
    .X(net1298));
 sky130_fd_sc_hd__buf_6 fanout1299 (.A(net53),
    .X(net1299));
 sky130_fd_sc_hd__buf_8 fanout1300 (.A(net1309),
    .X(net1300));
 sky130_fd_sc_hd__buf_6 fanout1301 (.A(net1303),
    .X(net1301));
 sky130_fd_sc_hd__clkbuf_4 fanout1302 (.A(net1303),
    .X(net1302));
 sky130_fd_sc_hd__buf_6 fanout1303 (.A(net1309),
    .X(net1303));
 sky130_fd_sc_hd__clkbuf_8 fanout1304 (.A(net1305),
    .X(net1304));
 sky130_fd_sc_hd__buf_4 fanout1305 (.A(net1308),
    .X(net1305));
 sky130_fd_sc_hd__buf_6 fanout1306 (.A(net1308),
    .X(net1306));
 sky130_fd_sc_hd__buf_6 fanout1307 (.A(net1308),
    .X(net1307));
 sky130_fd_sc_hd__buf_4 fanout1308 (.A(net1309),
    .X(net1308));
 sky130_fd_sc_hd__buf_4 fanout1309 (.A(net51),
    .X(net1309));
 sky130_fd_sc_hd__buf_6 fanout1310 (.A(net1311),
    .X(net1310));
 sky130_fd_sc_hd__buf_6 fanout1311 (.A(net5),
    .X(net1311));
 sky130_fd_sc_hd__buf_6 fanout1312 (.A(net1315),
    .X(net1312));
 sky130_fd_sc_hd__clkbuf_4 fanout1313 (.A(net1315),
    .X(net1313));
 sky130_fd_sc_hd__buf_6 fanout1314 (.A(net1315),
    .X(net1314));
 sky130_fd_sc_hd__buf_4 fanout1315 (.A(net5),
    .X(net1315));
 sky130_fd_sc_hd__buf_4 fanout1316 (.A(net1317),
    .X(net1316));
 sky130_fd_sc_hd__buf_6 fanout1317 (.A(net1318),
    .X(net1317));
 sky130_fd_sc_hd__buf_8 fanout1318 (.A(net5),
    .X(net1318));
 sky130_fd_sc_hd__buf_6 fanout1319 (.A(net1328),
    .X(net1319));
 sky130_fd_sc_hd__clkbuf_4 fanout1320 (.A(net1328),
    .X(net1320));
 sky130_fd_sc_hd__clkbuf_8 fanout1321 (.A(net1322),
    .X(net1321));
 sky130_fd_sc_hd__buf_4 fanout1322 (.A(net1323),
    .X(net1322));
 sky130_fd_sc_hd__buf_4 fanout1323 (.A(net1328),
    .X(net1323));
 sky130_fd_sc_hd__buf_6 fanout1324 (.A(net1325),
    .X(net1324));
 sky130_fd_sc_hd__buf_4 fanout1325 (.A(net1328),
    .X(net1325));
 sky130_fd_sc_hd__buf_6 fanout1326 (.A(net1327),
    .X(net1326));
 sky130_fd_sc_hd__buf_8 fanout1327 (.A(net1328),
    .X(net1327));
 sky130_fd_sc_hd__buf_6 fanout1328 (.A(net49),
    .X(net1328));
 sky130_fd_sc_hd__buf_6 fanout1329 (.A(net1332),
    .X(net1329));
 sky130_fd_sc_hd__buf_6 fanout1330 (.A(net1332),
    .X(net1330));
 sky130_fd_sc_hd__buf_6 fanout1331 (.A(net1332),
    .X(net1331));
 sky130_fd_sc_hd__buf_8 fanout1332 (.A(net47),
    .X(net1332));
 sky130_fd_sc_hd__buf_6 fanout1333 (.A(net1337),
    .X(net1333));
 sky130_fd_sc_hd__buf_6 fanout1334 (.A(net1336),
    .X(net1334));
 sky130_fd_sc_hd__buf_6 fanout1335 (.A(net1336),
    .X(net1335));
 sky130_fd_sc_hd__clkbuf_4 fanout1336 (.A(net1337),
    .X(net1336));
 sky130_fd_sc_hd__buf_6 fanout1337 (.A(net47),
    .X(net1337));
 sky130_fd_sc_hd__buf_6 fanout1338 (.A(net1347),
    .X(net1338));
 sky130_fd_sc_hd__clkbuf_4 fanout1339 (.A(net1347),
    .X(net1339));
 sky130_fd_sc_hd__buf_6 fanout1340 (.A(net1342),
    .X(net1340));
 sky130_fd_sc_hd__buf_6 fanout1341 (.A(net1347),
    .X(net1341));
 sky130_fd_sc_hd__clkbuf_4 fanout1342 (.A(net1347),
    .X(net1342));
 sky130_fd_sc_hd__clkbuf_8 fanout1343 (.A(net1346),
    .X(net1343));
 sky130_fd_sc_hd__buf_6 fanout1344 (.A(net1345),
    .X(net1344));
 sky130_fd_sc_hd__buf_6 fanout1345 (.A(net1346),
    .X(net1345));
 sky130_fd_sc_hd__buf_6 fanout1346 (.A(net1347),
    .X(net1346));
 sky130_fd_sc_hd__buf_4 fanout1347 (.A(net44),
    .X(net1347));
 sky130_fd_sc_hd__buf_6 fanout1348 (.A(net1349),
    .X(net1348));
 sky130_fd_sc_hd__clkbuf_8 fanout1349 (.A(net1352),
    .X(net1349));
 sky130_fd_sc_hd__buf_6 fanout1350 (.A(net1352),
    .X(net1350));
 sky130_fd_sc_hd__buf_6 fanout1351 (.A(net1352),
    .X(net1351));
 sky130_fd_sc_hd__buf_4 fanout1352 (.A(net42),
    .X(net1352));
 sky130_fd_sc_hd__buf_6 fanout1353 (.A(net1354),
    .X(net1353));
 sky130_fd_sc_hd__buf_4 fanout1354 (.A(net42),
    .X(net1354));
 sky130_fd_sc_hd__buf_6 fanout1355 (.A(net1356),
    .X(net1355));
 sky130_fd_sc_hd__buf_6 fanout1356 (.A(net42),
    .X(net1356));
 sky130_fd_sc_hd__buf_6 fanout1357 (.A(net1366),
    .X(net1357));
 sky130_fd_sc_hd__buf_6 fanout1358 (.A(net1366),
    .X(net1358));
 sky130_fd_sc_hd__buf_6 fanout1359 (.A(net1361),
    .X(net1359));
 sky130_fd_sc_hd__buf_6 fanout1360 (.A(net1361),
    .X(net1360));
 sky130_fd_sc_hd__clkbuf_4 fanout1361 (.A(net1366),
    .X(net1361));
 sky130_fd_sc_hd__buf_6 fanout1362 (.A(net1363),
    .X(net1362));
 sky130_fd_sc_hd__buf_4 fanout1363 (.A(net1366),
    .X(net1363));
 sky130_fd_sc_hd__buf_6 fanout1364 (.A(net1365),
    .X(net1364));
 sky130_fd_sc_hd__buf_4 fanout1365 (.A(net1366),
    .X(net1365));
 sky130_fd_sc_hd__buf_6 fanout1366 (.A(net40),
    .X(net1366));
 sky130_fd_sc_hd__buf_6 fanout1367 (.A(net1368),
    .X(net1367));
 sky130_fd_sc_hd__buf_6 fanout1368 (.A(net38),
    .X(net1368));
 sky130_fd_sc_hd__buf_4 fanout1369 (.A(net1370),
    .X(net1369));
 sky130_fd_sc_hd__buf_4 fanout1370 (.A(net1371),
    .X(net1370));
 sky130_fd_sc_hd__buf_6 fanout1371 (.A(net38),
    .X(net1371));
 sky130_fd_sc_hd__buf_6 fanout1372 (.A(net1375),
    .X(net1372));
 sky130_fd_sc_hd__buf_6 fanout1373 (.A(net1374),
    .X(net1373));
 sky130_fd_sc_hd__buf_4 fanout1374 (.A(net1375),
    .X(net1374));
 sky130_fd_sc_hd__buf_6 fanout1375 (.A(net38),
    .X(net1375));
 sky130_fd_sc_hd__buf_6 fanout1376 (.A(net1377),
    .X(net1376));
 sky130_fd_sc_hd__buf_6 fanout1377 (.A(net1384),
    .X(net1377));
 sky130_fd_sc_hd__buf_6 fanout1378 (.A(net1380),
    .X(net1378));
 sky130_fd_sc_hd__buf_4 fanout1379 (.A(net1380),
    .X(net1379));
 sky130_fd_sc_hd__buf_6 fanout1380 (.A(net1384),
    .X(net1380));
 sky130_fd_sc_hd__buf_6 fanout1381 (.A(net1384),
    .X(net1381));
 sky130_fd_sc_hd__buf_6 fanout1382 (.A(net1383),
    .X(net1382));
 sky130_fd_sc_hd__buf_4 fanout1383 (.A(net1384),
    .X(net1383));
 sky130_fd_sc_hd__clkbuf_16 fanout1384 (.A(net36),
    .X(net1384));
 sky130_fd_sc_hd__buf_6 fanout1385 (.A(net1386),
    .X(net1385));
 sky130_fd_sc_hd__buf_6 fanout1386 (.A(net1393),
    .X(net1386));
 sky130_fd_sc_hd__buf_6 fanout1387 (.A(net1388),
    .X(net1387));
 sky130_fd_sc_hd__buf_6 fanout1388 (.A(net1393),
    .X(net1388));
 sky130_fd_sc_hd__buf_6 fanout1389 (.A(net1391),
    .X(net1389));
 sky130_fd_sc_hd__clkbuf_8 fanout1390 (.A(net1391),
    .X(net1390));
 sky130_fd_sc_hd__buf_4 fanout1391 (.A(net1393),
    .X(net1391));
 sky130_fd_sc_hd__buf_6 fanout1392 (.A(net1393),
    .X(net1392));
 sky130_fd_sc_hd__buf_6 fanout1393 (.A(net34),
    .X(net1393));
 sky130_fd_sc_hd__buf_6 fanout1394 (.A(net33),
    .X(net1394));
 sky130_fd_sc_hd__buf_6 fanout1395 (.A(net33),
    .X(net1395));
 sky130_fd_sc_hd__buf_8 fanout1396 (.A(net1398),
    .X(net1396));
 sky130_fd_sc_hd__buf_6 fanout1397 (.A(net1398),
    .X(net1397));
 sky130_fd_sc_hd__clkbuf_4 fanout1398 (.A(net33),
    .X(net1398));
 sky130_fd_sc_hd__buf_6 fanout1399 (.A(net1402),
    .X(net1399));
 sky130_fd_sc_hd__buf_6 fanout1400 (.A(net1401),
    .X(net1400));
 sky130_fd_sc_hd__buf_4 fanout1401 (.A(net1402),
    .X(net1401));
 sky130_fd_sc_hd__buf_6 fanout1402 (.A(net33),
    .X(net1402));
 sky130_fd_sc_hd__buf_6 fanout1403 (.A(net1405),
    .X(net1403));
 sky130_fd_sc_hd__buf_4 fanout1404 (.A(net1405),
    .X(net1404));
 sky130_fd_sc_hd__buf_6 fanout1405 (.A(net1407),
    .X(net1405));
 sky130_fd_sc_hd__buf_6 fanout1406 (.A(net1407),
    .X(net1406));
 sky130_fd_sc_hd__clkbuf_4 fanout1407 (.A(net31),
    .X(net1407));
 sky130_fd_sc_hd__clkbuf_8 fanout1408 (.A(net1411),
    .X(net1408));
 sky130_fd_sc_hd__buf_6 fanout1409 (.A(net1411),
    .X(net1409));
 sky130_fd_sc_hd__buf_6 fanout1410 (.A(net1411),
    .X(net1410));
 sky130_fd_sc_hd__clkbuf_16 fanout1411 (.A(net31),
    .X(net1411));
 sky130_fd_sc_hd__buf_6 fanout1412 (.A(net3),
    .X(net1412));
 sky130_fd_sc_hd__buf_4 fanout1413 (.A(net3),
    .X(net1413));
 sky130_fd_sc_hd__clkbuf_8 fanout1414 (.A(net1415),
    .X(net1414));
 sky130_fd_sc_hd__buf_6 fanout1415 (.A(net1416),
    .X(net1415));
 sky130_fd_sc_hd__buf_6 fanout1416 (.A(net3),
    .X(net1416));
 sky130_fd_sc_hd__buf_4 fanout1417 (.A(net1418),
    .X(net1417));
 sky130_fd_sc_hd__buf_6 fanout1418 (.A(net1419),
    .X(net1418));
 sky130_fd_sc_hd__clkbuf_16 fanout1419 (.A(net3),
    .X(net1419));
 sky130_fd_sc_hd__buf_6 fanout1420 (.A(net1422),
    .X(net1420));
 sky130_fd_sc_hd__buf_4 fanout1421 (.A(net1422),
    .X(net1421));
 sky130_fd_sc_hd__buf_6 fanout1422 (.A(net1429),
    .X(net1422));
 sky130_fd_sc_hd__buf_6 fanout1423 (.A(net1424),
    .X(net1423));
 sky130_fd_sc_hd__buf_4 fanout1424 (.A(net1429),
    .X(net1424));
 sky130_fd_sc_hd__buf_6 fanout1425 (.A(net1427),
    .X(net1425));
 sky130_fd_sc_hd__buf_4 fanout1426 (.A(net1427),
    .X(net1426));
 sky130_fd_sc_hd__buf_6 fanout1427 (.A(net1429),
    .X(net1427));
 sky130_fd_sc_hd__buf_6 fanout1428 (.A(net1429),
    .X(net1428));
 sky130_fd_sc_hd__buf_8 fanout1429 (.A(net29),
    .X(net1429));
 sky130_fd_sc_hd__buf_6 fanout1430 (.A(net1431),
    .X(net1430));
 sky130_fd_sc_hd__buf_8 fanout1431 (.A(net1438),
    .X(net1431));
 sky130_fd_sc_hd__buf_6 fanout1432 (.A(net1433),
    .X(net1432));
 sky130_fd_sc_hd__buf_8 fanout1433 (.A(net1438),
    .X(net1433));
 sky130_fd_sc_hd__buf_6 fanout1434 (.A(net1436),
    .X(net1434));
 sky130_fd_sc_hd__buf_6 fanout1435 (.A(net1436),
    .X(net1435));
 sky130_fd_sc_hd__buf_4 fanout1436 (.A(net1437),
    .X(net1436));
 sky130_fd_sc_hd__clkbuf_16 fanout1437 (.A(net1438),
    .X(net1437));
 sky130_fd_sc_hd__buf_8 fanout1438 (.A(net27),
    .X(net1438));
 sky130_fd_sc_hd__buf_6 fanout1439 (.A(net1440),
    .X(net1439));
 sky130_fd_sc_hd__buf_8 fanout1440 (.A(net1443),
    .X(net1440));
 sky130_fd_sc_hd__buf_6 fanout1441 (.A(net1442),
    .X(net1441));
 sky130_fd_sc_hd__buf_8 fanout1442 (.A(net1443),
    .X(net1442));
 sky130_fd_sc_hd__buf_6 fanout1443 (.A(net1447),
    .X(net1443));
 sky130_fd_sc_hd__buf_6 fanout1444 (.A(net1445),
    .X(net1444));
 sky130_fd_sc_hd__buf_8 fanout1445 (.A(net1446),
    .X(net1445));
 sky130_fd_sc_hd__buf_8 fanout1446 (.A(net1447),
    .X(net1446));
 sky130_fd_sc_hd__buf_8 fanout1447 (.A(net25),
    .X(net1447));
 sky130_fd_sc_hd__buf_6 fanout1448 (.A(net1450),
    .X(net1448));
 sky130_fd_sc_hd__buf_4 fanout1449 (.A(net1450),
    .X(net1449));
 sky130_fd_sc_hd__buf_6 fanout1450 (.A(net1456),
    .X(net1450));
 sky130_fd_sc_hd__buf_6 fanout1451 (.A(net1452),
    .X(net1451));
 sky130_fd_sc_hd__buf_8 fanout1452 (.A(net1456),
    .X(net1452));
 sky130_fd_sc_hd__buf_6 fanout1453 (.A(net1454),
    .X(net1453));
 sky130_fd_sc_hd__buf_6 fanout1454 (.A(net1456),
    .X(net1454));
 sky130_fd_sc_hd__buf_6 fanout1455 (.A(net1456),
    .X(net1455));
 sky130_fd_sc_hd__buf_6 fanout1456 (.A(net22),
    .X(net1456));
 sky130_fd_sc_hd__buf_6 fanout1457 (.A(net1459),
    .X(net1457));
 sky130_fd_sc_hd__clkbuf_4 fanout1458 (.A(net1459),
    .X(net1458));
 sky130_fd_sc_hd__buf_6 fanout1459 (.A(net20),
    .X(net1459));
 sky130_fd_sc_hd__buf_6 fanout1460 (.A(net1462),
    .X(net1460));
 sky130_fd_sc_hd__buf_2 fanout1461 (.A(net1462),
    .X(net1461));
 sky130_fd_sc_hd__buf_6 fanout1462 (.A(net20),
    .X(net1462));
 sky130_fd_sc_hd__clkbuf_8 fanout1463 (.A(net1465),
    .X(net1463));
 sky130_fd_sc_hd__buf_8 fanout1464 (.A(net1465),
    .X(net1464));
 sky130_fd_sc_hd__buf_8 fanout1465 (.A(net20),
    .X(net1465));
 sky130_fd_sc_hd__buf_6 fanout1466 (.A(net1468),
    .X(net1466));
 sky130_fd_sc_hd__buf_4 fanout1467 (.A(net1468),
    .X(net1467));
 sky130_fd_sc_hd__buf_6 fanout1468 (.A(net18),
    .X(net1468));
 sky130_fd_sc_hd__buf_6 fanout1469 (.A(net1470),
    .X(net1469));
 sky130_fd_sc_hd__buf_6 fanout1470 (.A(net18),
    .X(net1470));
 sky130_fd_sc_hd__buf_4 fanout1471 (.A(net1472),
    .X(net1471));
 sky130_fd_sc_hd__clkbuf_4 fanout1472 (.A(net1473),
    .X(net1472));
 sky130_fd_sc_hd__buf_6 fanout1473 (.A(net1474),
    .X(net1473));
 sky130_fd_sc_hd__buf_8 fanout1474 (.A(net18),
    .X(net1474));
 sky130_fd_sc_hd__buf_6 fanout1475 (.A(net1477),
    .X(net1475));
 sky130_fd_sc_hd__clkbuf_4 fanout1476 (.A(net1477),
    .X(net1476));
 sky130_fd_sc_hd__buf_6 fanout1477 (.A(net16),
    .X(net1477));
 sky130_fd_sc_hd__buf_6 fanout1478 (.A(net1480),
    .X(net1478));
 sky130_fd_sc_hd__clkbuf_4 fanout1479 (.A(net1480),
    .X(net1479));
 sky130_fd_sc_hd__buf_6 fanout1480 (.A(net16),
    .X(net1480));
 sky130_fd_sc_hd__buf_4 fanout1481 (.A(net1482),
    .X(net1481));
 sky130_fd_sc_hd__buf_4 fanout1482 (.A(net1483),
    .X(net1482));
 sky130_fd_sc_hd__buf_8 fanout1483 (.A(net1484),
    .X(net1483));
 sky130_fd_sc_hd__buf_6 fanout1484 (.A(net16),
    .X(net1484));
 sky130_fd_sc_hd__buf_6 fanout1485 (.A(net1486),
    .X(net1485));
 sky130_fd_sc_hd__buf_6 fanout1486 (.A(net1490),
    .X(net1486));
 sky130_fd_sc_hd__buf_6 fanout1487 (.A(net1489),
    .X(net1487));
 sky130_fd_sc_hd__clkbuf_4 fanout1488 (.A(net1489),
    .X(net1488));
 sky130_fd_sc_hd__buf_6 fanout1489 (.A(net1490),
    .X(net1489));
 sky130_fd_sc_hd__buf_4 fanout1490 (.A(net14),
    .X(net1490));
 sky130_fd_sc_hd__clkbuf_8 fanout1491 (.A(net1492),
    .X(net1491));
 sky130_fd_sc_hd__buf_6 fanout1492 (.A(net1493),
    .X(net1492));
 sky130_fd_sc_hd__buf_8 fanout1493 (.A(net14),
    .X(net1493));
 sky130_fd_sc_hd__buf_4 fanout1494 (.A(net1495),
    .X(net1494));
 sky130_fd_sc_hd__buf_2 fanout1495 (.A(net1498),
    .X(net1495));
 sky130_fd_sc_hd__buf_4 fanout1496 (.A(net1498),
    .X(net1496));
 sky130_fd_sc_hd__buf_2 fanout1497 (.A(net1498),
    .X(net1497));
 sky130_fd_sc_hd__buf_6 fanout1498 (.A(net1502),
    .X(net1498));
 sky130_fd_sc_hd__buf_4 fanout1499 (.A(net1501),
    .X(net1499));
 sky130_fd_sc_hd__clkbuf_4 fanout1500 (.A(net1501),
    .X(net1500));
 sky130_fd_sc_hd__clkbuf_8 fanout1501 (.A(net1502),
    .X(net1501));
 sky130_fd_sc_hd__buf_6 fanout1502 (.A(net128),
    .X(net1502));
 sky130_fd_sc_hd__buf_4 fanout1503 (.A(net1506),
    .X(net1503));
 sky130_fd_sc_hd__buf_2 fanout1504 (.A(net1506),
    .X(net1504));
 sky130_fd_sc_hd__buf_4 fanout1505 (.A(net1506),
    .X(net1505));
 sky130_fd_sc_hd__clkbuf_4 fanout1506 (.A(net1507),
    .X(net1506));
 sky130_fd_sc_hd__buf_6 fanout1507 (.A(net127),
    .X(net1507));
 sky130_fd_sc_hd__buf_4 fanout1508 (.A(net1510),
    .X(net1508));
 sky130_fd_sc_hd__buf_4 fanout1509 (.A(net1510),
    .X(net1509));
 sky130_fd_sc_hd__buf_6 fanout1510 (.A(net127),
    .X(net1510));
 sky130_fd_sc_hd__buf_4 fanout1511 (.A(net1514),
    .X(net1511));
 sky130_fd_sc_hd__clkbuf_2 fanout1512 (.A(net1514),
    .X(net1512));
 sky130_fd_sc_hd__buf_4 fanout1513 (.A(net1514),
    .X(net1513));
 sky130_fd_sc_hd__buf_6 fanout1514 (.A(net1518),
    .X(net1514));
 sky130_fd_sc_hd__buf_4 fanout1515 (.A(net1516),
    .X(net1515));
 sky130_fd_sc_hd__buf_4 fanout1516 (.A(net1518),
    .X(net1516));
 sky130_fd_sc_hd__buf_4 fanout1517 (.A(net1518),
    .X(net1517));
 sky130_fd_sc_hd__buf_8 fanout1518 (.A(net126),
    .X(net1518));
 sky130_fd_sc_hd__buf_4 fanout1519 (.A(net1521),
    .X(net1519));
 sky130_fd_sc_hd__buf_2 fanout1520 (.A(net1521),
    .X(net1520));
 sky130_fd_sc_hd__buf_4 fanout1521 (.A(net1522),
    .X(net1521));
 sky130_fd_sc_hd__buf_6 fanout1522 (.A(net125),
    .X(net1522));
 sky130_fd_sc_hd__buf_4 fanout1523 (.A(net1524),
    .X(net1523));
 sky130_fd_sc_hd__buf_4 fanout1524 (.A(net1526),
    .X(net1524));
 sky130_fd_sc_hd__buf_4 fanout1525 (.A(net1526),
    .X(net1525));
 sky130_fd_sc_hd__buf_4 fanout1526 (.A(net125),
    .X(net1526));
 sky130_fd_sc_hd__buf_4 fanout1527 (.A(net1530),
    .X(net1527));
 sky130_fd_sc_hd__buf_4 fanout1528 (.A(net1530),
    .X(net1528));
 sky130_fd_sc_hd__buf_2 fanout1529 (.A(net1530),
    .X(net1529));
 sky130_fd_sc_hd__buf_4 fanout1530 (.A(net124),
    .X(net1530));
 sky130_fd_sc_hd__buf_4 fanout1531 (.A(net124),
    .X(net1531));
 sky130_fd_sc_hd__buf_4 fanout1532 (.A(net1534),
    .X(net1532));
 sky130_fd_sc_hd__buf_2 fanout1533 (.A(net1534),
    .X(net1533));
 sky130_fd_sc_hd__buf_4 fanout1534 (.A(net124),
    .X(net1534));
 sky130_fd_sc_hd__buf_4 fanout1535 (.A(net1538),
    .X(net1535));
 sky130_fd_sc_hd__buf_4 fanout1536 (.A(net1538),
    .X(net1536));
 sky130_fd_sc_hd__buf_2 fanout1537 (.A(net1538),
    .X(net1537));
 sky130_fd_sc_hd__buf_6 fanout1538 (.A(net123),
    .X(net1538));
 sky130_fd_sc_hd__buf_4 fanout1539 (.A(net123),
    .X(net1539));
 sky130_fd_sc_hd__buf_4 fanout1540 (.A(net1542),
    .X(net1540));
 sky130_fd_sc_hd__clkbuf_4 fanout1541 (.A(net1542),
    .X(net1541));
 sky130_fd_sc_hd__buf_4 fanout1542 (.A(net123),
    .X(net1542));
 sky130_fd_sc_hd__buf_4 fanout1543 (.A(net1546),
    .X(net1543));
 sky130_fd_sc_hd__buf_4 fanout1544 (.A(net1546),
    .X(net1544));
 sky130_fd_sc_hd__buf_2 fanout1545 (.A(net1546),
    .X(net1545));
 sky130_fd_sc_hd__buf_4 fanout1546 (.A(net122),
    .X(net1546));
 sky130_fd_sc_hd__buf_4 fanout1547 (.A(net122),
    .X(net1547));
 sky130_fd_sc_hd__buf_4 fanout1548 (.A(net1550),
    .X(net1548));
 sky130_fd_sc_hd__clkbuf_4 fanout1549 (.A(net1550),
    .X(net1549));
 sky130_fd_sc_hd__buf_4 fanout1550 (.A(net122),
    .X(net1550));
 sky130_fd_sc_hd__buf_4 fanout1551 (.A(net1552),
    .X(net1551));
 sky130_fd_sc_hd__clkbuf_4 fanout1552 (.A(net1559),
    .X(net1552));
 sky130_fd_sc_hd__buf_4 fanout1553 (.A(net1559),
    .X(net1553));
 sky130_fd_sc_hd__buf_2 fanout1554 (.A(net1559),
    .X(net1554));
 sky130_fd_sc_hd__buf_6 fanout1555 (.A(net1559),
    .X(net1555));
 sky130_fd_sc_hd__buf_4 fanout1556 (.A(net1557),
    .X(net1556));
 sky130_fd_sc_hd__clkbuf_8 fanout1557 (.A(net1559),
    .X(net1557));
 sky130_fd_sc_hd__buf_2 fanout1558 (.A(net1559),
    .X(net1558));
 sky130_fd_sc_hd__buf_8 fanout1559 (.A(net121),
    .X(net1559));
 sky130_fd_sc_hd__clkbuf_4 fanout1560 (.A(net1562),
    .X(net1560));
 sky130_fd_sc_hd__buf_4 fanout1561 (.A(net1562),
    .X(net1561));
 sky130_fd_sc_hd__buf_4 fanout1562 (.A(net1563),
    .X(net1562));
 sky130_fd_sc_hd__clkbuf_8 fanout1563 (.A(net120),
    .X(net1563));
 sky130_fd_sc_hd__buf_4 fanout1564 (.A(net1565),
    .X(net1564));
 sky130_fd_sc_hd__clkbuf_8 fanout1565 (.A(net1567),
    .X(net1565));
 sky130_fd_sc_hd__buf_6 fanout1566 (.A(net1567),
    .X(net1566));
 sky130_fd_sc_hd__buf_6 fanout1567 (.A(net120),
    .X(net1567));
 sky130_fd_sc_hd__buf_6 fanout1568 (.A(net1577),
    .X(net1568));
 sky130_fd_sc_hd__clkbuf_4 fanout1569 (.A(net1577),
    .X(net1569));
 sky130_fd_sc_hd__buf_6 fanout1570 (.A(net1572),
    .X(net1570));
 sky130_fd_sc_hd__buf_2 fanout1571 (.A(net1572),
    .X(net1571));
 sky130_fd_sc_hd__buf_4 fanout1572 (.A(net1577),
    .X(net1572));
 sky130_fd_sc_hd__buf_4 fanout1573 (.A(net1574),
    .X(net1573));
 sky130_fd_sc_hd__buf_4 fanout1574 (.A(net1575),
    .X(net1574));
 sky130_fd_sc_hd__buf_6 fanout1575 (.A(net1576),
    .X(net1575));
 sky130_fd_sc_hd__buf_6 fanout1576 (.A(net1577),
    .X(net1576));
 sky130_fd_sc_hd__buf_6 fanout1577 (.A(net12),
    .X(net1577));
 sky130_fd_sc_hd__buf_4 fanout1578 (.A(net1581),
    .X(net1578));
 sky130_fd_sc_hd__buf_4 fanout1579 (.A(net1581),
    .X(net1579));
 sky130_fd_sc_hd__clkbuf_4 fanout1580 (.A(net1581),
    .X(net1580));
 sky130_fd_sc_hd__buf_4 fanout1581 (.A(net119),
    .X(net1581));
 sky130_fd_sc_hd__clkbuf_8 fanout1582 (.A(net1585),
    .X(net1582));
 sky130_fd_sc_hd__buf_4 fanout1583 (.A(net1584),
    .X(net1583));
 sky130_fd_sc_hd__buf_4 fanout1584 (.A(net1585),
    .X(net1584));
 sky130_fd_sc_hd__buf_4 fanout1585 (.A(net119),
    .X(net1585));
 sky130_fd_sc_hd__buf_4 fanout1586 (.A(net1594),
    .X(net1586));
 sky130_fd_sc_hd__buf_2 fanout1587 (.A(net1594),
    .X(net1587));
 sky130_fd_sc_hd__buf_4 fanout1588 (.A(net1594),
    .X(net1588));
 sky130_fd_sc_hd__buf_2 fanout1589 (.A(net1594),
    .X(net1589));
 sky130_fd_sc_hd__buf_6 fanout1590 (.A(net1593),
    .X(net1590));
 sky130_fd_sc_hd__buf_4 fanout1591 (.A(net1592),
    .X(net1591));
 sky130_fd_sc_hd__clkbuf_8 fanout1592 (.A(net1593),
    .X(net1592));
 sky130_fd_sc_hd__buf_4 fanout1593 (.A(net1594),
    .X(net1593));
 sky130_fd_sc_hd__buf_6 fanout1594 (.A(net118),
    .X(net1594));
 sky130_fd_sc_hd__buf_4 fanout1595 (.A(net1598),
    .X(net1595));
 sky130_fd_sc_hd__buf_2 fanout1596 (.A(net1598),
    .X(net1596));
 sky130_fd_sc_hd__buf_4 fanout1597 (.A(net1598),
    .X(net1597));
 sky130_fd_sc_hd__buf_4 fanout1598 (.A(net117),
    .X(net1598));
 sky130_fd_sc_hd__clkbuf_8 fanout1599 (.A(net1603),
    .X(net1599));
 sky130_fd_sc_hd__buf_4 fanout1600 (.A(net1602),
    .X(net1600));
 sky130_fd_sc_hd__buf_2 fanout1601 (.A(net1602),
    .X(net1601));
 sky130_fd_sc_hd__buf_4 fanout1602 (.A(net1603),
    .X(net1602));
 sky130_fd_sc_hd__clkbuf_4 fanout1603 (.A(net117),
    .X(net1603));
 sky130_fd_sc_hd__buf_4 fanout1604 (.A(net1606),
    .X(net1604));
 sky130_fd_sc_hd__buf_4 fanout1605 (.A(net1606),
    .X(net1605));
 sky130_fd_sc_hd__buf_6 fanout1606 (.A(net116),
    .X(net1606));
 sky130_fd_sc_hd__buf_4 fanout1607 (.A(net1611),
    .X(net1607));
 sky130_fd_sc_hd__buf_4 fanout1608 (.A(net1610),
    .X(net1608));
 sky130_fd_sc_hd__buf_4 fanout1609 (.A(net1610),
    .X(net1609));
 sky130_fd_sc_hd__clkbuf_4 fanout1610 (.A(net1611),
    .X(net1610));
 sky130_fd_sc_hd__clkbuf_4 fanout1611 (.A(net116),
    .X(net1611));
 sky130_fd_sc_hd__buf_4 fanout1612 (.A(net1614),
    .X(net1612));
 sky130_fd_sc_hd__clkbuf_8 fanout1613 (.A(net1614),
    .X(net1613));
 sky130_fd_sc_hd__buf_4 fanout1614 (.A(net115),
    .X(net1614));
 sky130_fd_sc_hd__buf_4 fanout1615 (.A(net1619),
    .X(net1615));
 sky130_fd_sc_hd__buf_4 fanout1616 (.A(net1619),
    .X(net1616));
 sky130_fd_sc_hd__clkbuf_2 fanout1617 (.A(net1619),
    .X(net1617));
 sky130_fd_sc_hd__buf_4 fanout1618 (.A(net1619),
    .X(net1618));
 sky130_fd_sc_hd__buf_6 fanout1619 (.A(net115),
    .X(net1619));
 sky130_fd_sc_hd__buf_4 fanout1620 (.A(net1621),
    .X(net1620));
 sky130_fd_sc_hd__buf_4 fanout1621 (.A(net1628),
    .X(net1621));
 sky130_fd_sc_hd__clkbuf_8 fanout1622 (.A(net1628),
    .X(net1622));
 sky130_fd_sc_hd__buf_4 fanout1623 (.A(net1627),
    .X(net1623));
 sky130_fd_sc_hd__buf_4 fanout1624 (.A(net1626),
    .X(net1624));
 sky130_fd_sc_hd__buf_2 fanout1625 (.A(net1626),
    .X(net1625));
 sky130_fd_sc_hd__buf_4 fanout1626 (.A(net1627),
    .X(net1626));
 sky130_fd_sc_hd__buf_4 fanout1627 (.A(net1628),
    .X(net1627));
 sky130_fd_sc_hd__buf_4 fanout1628 (.A(net114),
    .X(net1628));
 sky130_fd_sc_hd__buf_4 fanout1629 (.A(net1630),
    .X(net1629));
 sky130_fd_sc_hd__buf_4 fanout1630 (.A(net1632),
    .X(net1630));
 sky130_fd_sc_hd__buf_6 fanout1631 (.A(net1632),
    .X(net1631));
 sky130_fd_sc_hd__clkbuf_4 fanout1632 (.A(net113),
    .X(net1632));
 sky130_fd_sc_hd__clkbuf_8 fanout1633 (.A(net1637),
    .X(net1633));
 sky130_fd_sc_hd__buf_4 fanout1634 (.A(net1636),
    .X(net1634));
 sky130_fd_sc_hd__buf_4 fanout1635 (.A(net1636),
    .X(net1635));
 sky130_fd_sc_hd__clkbuf_4 fanout1636 (.A(net1637),
    .X(net1636));
 sky130_fd_sc_hd__buf_4 fanout1637 (.A(net113),
    .X(net1637));
 sky130_fd_sc_hd__buf_6 fanout1638 (.A(net1640),
    .X(net1638));
 sky130_fd_sc_hd__buf_6 fanout1639 (.A(net1640),
    .X(net1639));
 sky130_fd_sc_hd__buf_6 fanout1640 (.A(net112),
    .X(net1640));
 sky130_fd_sc_hd__buf_4 fanout1641 (.A(net112),
    .X(net1641));
 sky130_fd_sc_hd__clkbuf_4 fanout1642 (.A(net112),
    .X(net1642));
 sky130_fd_sc_hd__buf_4 fanout1643 (.A(net1645),
    .X(net1643));
 sky130_fd_sc_hd__buf_4 fanout1644 (.A(net1645),
    .X(net1644));
 sky130_fd_sc_hd__buf_2 fanout1645 (.A(net112),
    .X(net1645));
 sky130_fd_sc_hd__clkbuf_8 fanout1646 (.A(net1648),
    .X(net1646));
 sky130_fd_sc_hd__buf_6 fanout1647 (.A(net1648),
    .X(net1647));
 sky130_fd_sc_hd__buf_6 fanout1648 (.A(net111),
    .X(net1648));
 sky130_fd_sc_hd__clkbuf_8 fanout1649 (.A(net111),
    .X(net1649));
 sky130_fd_sc_hd__clkbuf_4 fanout1650 (.A(net111),
    .X(net1650));
 sky130_fd_sc_hd__buf_4 fanout1651 (.A(net1653),
    .X(net1651));
 sky130_fd_sc_hd__buf_4 fanout1652 (.A(net1653),
    .X(net1652));
 sky130_fd_sc_hd__clkbuf_4 fanout1653 (.A(net111),
    .X(net1653));
 sky130_fd_sc_hd__buf_4 fanout1654 (.A(net1656),
    .X(net1654));
 sky130_fd_sc_hd__clkbuf_8 fanout1655 (.A(net1656),
    .X(net1655));
 sky130_fd_sc_hd__clkbuf_8 fanout1656 (.A(net110),
    .X(net1656));
 sky130_fd_sc_hd__buf_4 fanout1657 (.A(net110),
    .X(net1657));
 sky130_fd_sc_hd__buf_2 fanout1658 (.A(net110),
    .X(net1658));
 sky130_fd_sc_hd__clkbuf_8 fanout1659 (.A(net1661),
    .X(net1659));
 sky130_fd_sc_hd__buf_4 fanout1660 (.A(net1661),
    .X(net1660));
 sky130_fd_sc_hd__clkbuf_4 fanout1661 (.A(net110),
    .X(net1661));
 sky130_fd_sc_hd__buf_6 fanout1662 (.A(net1667),
    .X(net1662));
 sky130_fd_sc_hd__buf_6 fanout1663 (.A(net1667),
    .X(net1663));
 sky130_fd_sc_hd__buf_6 fanout1664 (.A(net1666),
    .X(net1664));
 sky130_fd_sc_hd__clkbuf_4 fanout1665 (.A(net1666),
    .X(net1665));
 sky130_fd_sc_hd__buf_6 fanout1666 (.A(net1667),
    .X(net1666));
 sky130_fd_sc_hd__buf_6 fanout1667 (.A(net11),
    .X(net1667));
 sky130_fd_sc_hd__buf_6 fanout1668 (.A(net1669),
    .X(net1668));
 sky130_fd_sc_hd__buf_8 fanout1669 (.A(net1670),
    .X(net1669));
 sky130_fd_sc_hd__buf_6 fanout1670 (.A(net11),
    .X(net1670));
 sky130_fd_sc_hd__buf_4 fanout1671 (.A(net1673),
    .X(net1671));
 sky130_fd_sc_hd__buf_4 fanout1672 (.A(net1673),
    .X(net1672));
 sky130_fd_sc_hd__clkbuf_4 fanout1673 (.A(net1674),
    .X(net1673));
 sky130_fd_sc_hd__buf_4 fanout1674 (.A(net109),
    .X(net1674));
 sky130_fd_sc_hd__clkbuf_4 fanout1675 (.A(net1678),
    .X(net1675));
 sky130_fd_sc_hd__buf_4 fanout1676 (.A(net1678),
    .X(net1676));
 sky130_fd_sc_hd__buf_6 fanout1677 (.A(net1678),
    .X(net1677));
 sky130_fd_sc_hd__buf_6 fanout1678 (.A(net109),
    .X(net1678));
 sky130_fd_sc_hd__buf_4 fanout1679 (.A(net1681),
    .X(net1679));
 sky130_fd_sc_hd__buf_6 fanout1680 (.A(net1681),
    .X(net1680));
 sky130_fd_sc_hd__buf_6 fanout1681 (.A(net108),
    .X(net1681));
 sky130_fd_sc_hd__buf_4 fanout1682 (.A(net1683),
    .X(net1682));
 sky130_fd_sc_hd__buf_4 fanout1683 (.A(net108),
    .X(net1683));
 sky130_fd_sc_hd__buf_4 fanout1684 (.A(net1686),
    .X(net1684));
 sky130_fd_sc_hd__buf_4 fanout1685 (.A(net108),
    .X(net1685));
 sky130_fd_sc_hd__buf_2 fanout1686 (.A(net108),
    .X(net1686));
 sky130_fd_sc_hd__buf_4 fanout1687 (.A(net1689),
    .X(net1687));
 sky130_fd_sc_hd__buf_6 fanout1688 (.A(net1689),
    .X(net1688));
 sky130_fd_sc_hd__buf_4 fanout1689 (.A(net107),
    .X(net1689));
 sky130_fd_sc_hd__buf_4 fanout1690 (.A(net107),
    .X(net1690));
 sky130_fd_sc_hd__clkbuf_4 fanout1691 (.A(net107),
    .X(net1691));
 sky130_fd_sc_hd__buf_6 fanout1692 (.A(net1694),
    .X(net1692));
 sky130_fd_sc_hd__buf_4 fanout1693 (.A(net1694),
    .X(net1693));
 sky130_fd_sc_hd__clkbuf_4 fanout1694 (.A(net107),
    .X(net1694));
 sky130_fd_sc_hd__buf_6 fanout1695 (.A(net1697),
    .X(net1695));
 sky130_fd_sc_hd__buf_4 fanout1696 (.A(net1697),
    .X(net1696));
 sky130_fd_sc_hd__buf_6 fanout1697 (.A(net106),
    .X(net1697));
 sky130_fd_sc_hd__buf_6 fanout1698 (.A(net106),
    .X(net1698));
 sky130_fd_sc_hd__clkbuf_2 fanout1699 (.A(net106),
    .X(net1699));
 sky130_fd_sc_hd__buf_4 fanout1700 (.A(net1702),
    .X(net1700));
 sky130_fd_sc_hd__clkbuf_2 fanout1701 (.A(net1702),
    .X(net1701));
 sky130_fd_sc_hd__buf_6 fanout1702 (.A(net106),
    .X(net1702));
 sky130_fd_sc_hd__buf_4 fanout1703 (.A(net1705),
    .X(net1703));
 sky130_fd_sc_hd__buf_4 fanout1704 (.A(net1705),
    .X(net1704));
 sky130_fd_sc_hd__buf_6 fanout1705 (.A(net105),
    .X(net1705));
 sky130_fd_sc_hd__buf_8 fanout1706 (.A(net105),
    .X(net1706));
 sky130_fd_sc_hd__clkbuf_2 fanout1707 (.A(net105),
    .X(net1707));
 sky130_fd_sc_hd__buf_4 fanout1708 (.A(net1710),
    .X(net1708));
 sky130_fd_sc_hd__clkbuf_2 fanout1709 (.A(net1710),
    .X(net1709));
 sky130_fd_sc_hd__buf_6 fanout1710 (.A(net105),
    .X(net1710));
 sky130_fd_sc_hd__buf_4 fanout1711 (.A(net1714),
    .X(net1711));
 sky130_fd_sc_hd__clkbuf_4 fanout1712 (.A(net1714),
    .X(net1712));
 sky130_fd_sc_hd__buf_4 fanout1713 (.A(net1714),
    .X(net1713));
 sky130_fd_sc_hd__buf_4 fanout1714 (.A(net104),
    .X(net1714));
 sky130_fd_sc_hd__buf_6 fanout1715 (.A(net104),
    .X(net1715));
 sky130_fd_sc_hd__clkbuf_2 fanout1716 (.A(net104),
    .X(net1716));
 sky130_fd_sc_hd__buf_4 fanout1717 (.A(net1719),
    .X(net1717));
 sky130_fd_sc_hd__clkbuf_2 fanout1718 (.A(net1719),
    .X(net1718));
 sky130_fd_sc_hd__buf_6 fanout1719 (.A(net104),
    .X(net1719));
 sky130_fd_sc_hd__buf_4 fanout1720 (.A(net1723),
    .X(net1720));
 sky130_fd_sc_hd__clkbuf_4 fanout1721 (.A(net1723),
    .X(net1721));
 sky130_fd_sc_hd__buf_4 fanout1722 (.A(net1723),
    .X(net1722));
 sky130_fd_sc_hd__buf_4 fanout1723 (.A(net103),
    .X(net1723));
 sky130_fd_sc_hd__buf_4 fanout1724 (.A(net1728),
    .X(net1724));
 sky130_fd_sc_hd__clkbuf_4 fanout1725 (.A(net1728),
    .X(net1725));
 sky130_fd_sc_hd__buf_4 fanout1726 (.A(net1727),
    .X(net1726));
 sky130_fd_sc_hd__buf_6 fanout1727 (.A(net1728),
    .X(net1727));
 sky130_fd_sc_hd__buf_4 fanout1728 (.A(net103),
    .X(net1728));
 sky130_fd_sc_hd__buf_4 fanout1729 (.A(net1732),
    .X(net1729));
 sky130_fd_sc_hd__clkbuf_4 fanout1730 (.A(net1732),
    .X(net1730));
 sky130_fd_sc_hd__buf_4 fanout1731 (.A(net1732),
    .X(net1731));
 sky130_fd_sc_hd__buf_4 fanout1732 (.A(net102),
    .X(net1732));
 sky130_fd_sc_hd__buf_6 fanout1733 (.A(net1736),
    .X(net1733));
 sky130_fd_sc_hd__buf_4 fanout1734 (.A(net1735),
    .X(net1734));
 sky130_fd_sc_hd__buf_6 fanout1735 (.A(net1736),
    .X(net1735));
 sky130_fd_sc_hd__buf_6 fanout1736 (.A(net102),
    .X(net1736));
 sky130_fd_sc_hd__buf_4 fanout1737 (.A(net1738),
    .X(net1737));
 sky130_fd_sc_hd__buf_6 fanout1738 (.A(net101),
    .X(net1738));
 sky130_fd_sc_hd__buf_6 fanout1739 (.A(net101),
    .X(net1739));
 sky130_fd_sc_hd__clkbuf_4 fanout1740 (.A(net101),
    .X(net1740));
 sky130_fd_sc_hd__buf_6 fanout1741 (.A(net1744),
    .X(net1741));
 sky130_fd_sc_hd__buf_4 fanout1742 (.A(net1743),
    .X(net1742));
 sky130_fd_sc_hd__buf_4 fanout1743 (.A(net1744),
    .X(net1743));
 sky130_fd_sc_hd__buf_4 fanout1744 (.A(net101),
    .X(net1744));
 sky130_fd_sc_hd__clkbuf_4 fanout1745 (.A(net1746),
    .X(net1745));
 sky130_fd_sc_hd__buf_6 fanout1746 (.A(net1752),
    .X(net1746));
 sky130_fd_sc_hd__buf_6 fanout1747 (.A(net1752),
    .X(net1747));
 sky130_fd_sc_hd__clkbuf_4 fanout1748 (.A(net1752),
    .X(net1748));
 sky130_fd_sc_hd__buf_6 fanout1749 (.A(net1752),
    .X(net1749));
 sky130_fd_sc_hd__buf_4 fanout1750 (.A(net1751),
    .X(net1750));
 sky130_fd_sc_hd__buf_4 fanout1751 (.A(net1752),
    .X(net1751));
 sky130_fd_sc_hd__buf_12 fanout1752 (.A(net100),
    .X(net1752));
 sky130_fd_sc_hd__conb_1 \U$$0_1753  (.LO(net1753));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_199_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_201_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_202_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_206_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_207_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_210_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_212_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_214_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_215_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_216_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_217_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_218_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_219_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_220_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_222_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_223_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_224_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_226_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_227_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_228_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_229_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_230_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_231_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_232_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_233_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_234_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_235_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_236_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_237_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_238_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_239_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_240_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_241_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_242_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_243_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_244_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_245_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_246_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_247_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_248_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_249_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_250_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_251_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_0__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_1__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_2__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_3__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_4__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_5__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_6__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_7__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_8__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_8__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_9__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_9__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_10__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_10__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_11__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_11__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_12__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_12__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_13__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_14__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_14__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_15__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_15__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_16__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_16__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_17__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_17__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_18__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_18__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_19__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_19__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_20__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_20__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_21__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_21__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_22__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_22__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_23__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_23__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_24__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_24__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_25__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_25__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_26__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_26__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_27__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_28__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_28__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_29__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_29__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_30__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_30__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_31__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_31__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\c$1338 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\c$1388 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\c$4184 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\c$4188 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\c$4238 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\c$4240 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\c$628 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\final_adder.g_new$855 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\final_adder.g_new$967 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\final_adder.g_new$987 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\final_adder.p_new$734 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(pp_row54_29));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(pp_row55_28));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\s$4323 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\s$4405 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\sel_0$4477 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\sel_0$5107 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\sel_0$5177 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\sel_0$5247 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\sel_0$6227 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\sel_1$4478 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(net891));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(net1234));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(net1234));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(net1252));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(net1253));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(net1290));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(net1309));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(net1366));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(net1384));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(net1384));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(net1429));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(net1447));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(net1487));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(net1506));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(net1522));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(net1522));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(net1567));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(net1567));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(net1594));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(net1594));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(net1594));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(net1594));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(net1619));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(net1619));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(net1619));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(net1619));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(net1640));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(net1667));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(net1674));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(net1723));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(net1723));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(net1723));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(net1723));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(net1728));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(net1728));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(net1728));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(net1732));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(net1741));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(net1744));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(net1752));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(net1752));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(net1752));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(\c$1412 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(\c$4206 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(\c$4210 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(\c$4212 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(\c$4242 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(\c$580 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(\final_adder.p_new$604 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(\final_adder.p_new$840 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(pp_row46_25));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(\s$4213 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(\s$4217 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(\sel_1$4968 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(\sel_1$5038 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(\sel_1$5248 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(\sel_1$6228 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_328 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_329 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_330 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_331 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_332 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA_333 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_334 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_335 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_336 (.DIODE(net740));
 sky130_fd_sc_hd__diode_2 ANTENNA_337 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA_338 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA_339 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_340 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_341 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_342 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_343 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_344 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_345 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_346 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_347 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_348 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_349 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_350 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_351 (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_352 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_353 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_354 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_355 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_356 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_357 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_358 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_359 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_360 (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_361 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_362 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_363 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_364 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_365 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_366 (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_367 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_368 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_369 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_370 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_371 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_372 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA_373 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA_374 (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA_375 (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA_376 (.DIODE(net1184));
 sky130_fd_sc_hd__diode_2 ANTENNA_377 (.DIODE(net1195));
 sky130_fd_sc_hd__diode_2 ANTENNA_378 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA_379 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA_380 (.DIODE(net1299));
 sky130_fd_sc_hd__diode_2 ANTENNA_381 (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA_382 (.DIODE(net1393));
 sky130_fd_sc_hd__diode_2 ANTENNA_383 (.DIODE(net1429));
 sky130_fd_sc_hd__diode_2 ANTENNA_384 (.DIODE(net1462));
 sky130_fd_sc_hd__diode_2 ANTENNA_385 (.DIODE(net1464));
 sky130_fd_sc_hd__diode_2 ANTENNA_386 (.DIODE(net1470));
 sky130_fd_sc_hd__diode_2 ANTENNA_387 (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA_388 (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA_389 (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA_390 (.DIODE(net1518));
 sky130_fd_sc_hd__diode_2 ANTENNA_391 (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA_392 (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA_393 (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA_394 (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA_395 (.DIODE(net1546));
 sky130_fd_sc_hd__diode_2 ANTENNA_396 (.DIODE(net1552));
 sky130_fd_sc_hd__diode_2 ANTENNA_397 (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA_398 (.DIODE(net1627));
 sky130_fd_sc_hd__diode_2 ANTENNA_399 (.DIODE(net1627));
 sky130_fd_sc_hd__diode_2 ANTENNA_400 (.DIODE(net1631));
 sky130_fd_sc_hd__diode_2 ANTENNA_401 (.DIODE(net1639));
 sky130_fd_sc_hd__diode_2 ANTENNA_402 (.DIODE(net1650));
 sky130_fd_sc_hd__diode_2 ANTENNA_403 (.DIODE(net1667));
 sky130_fd_sc_hd__diode_2 ANTENNA_404 (.DIODE(net1683));
 sky130_fd_sc_hd__diode_2 ANTENNA_405 (.DIODE(net1714));
 sky130_fd_sc_hd__diode_2 ANTENNA_406 (.DIODE(net1714));
 sky130_fd_sc_hd__diode_2 ANTENNA_407 (.DIODE(net1714));
 sky130_fd_sc_hd__diode_2 ANTENNA_408 (.DIODE(net1714));
 sky130_fd_sc_hd__diode_2 ANTENNA_409 (.DIODE(net1732));
 sky130_fd_sc_hd__diode_2 ANTENNA_410 (.DIODE(net1732));
 sky130_fd_sc_hd__diode_2 ANTENNA_411 (.DIODE(net1752));
 sky130_fd_sc_hd__diode_2 ANTENNA_412 (.DIODE(net1752));
 sky130_fd_sc_hd__diode_2 ANTENNA_413 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_414 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_415 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_416 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_417 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_418 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_419 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA_420 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_421 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_422 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_423 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA_424 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_425 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_426 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_427 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_428 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_429 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA_430 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_431 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_432 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_433 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_434 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_435 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_436 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_437 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_438 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_439 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_440 (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_441 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_442 (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_443 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_444 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_445 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_446 (.DIODE(net1480));
 sky130_fd_sc_hd__diode_2 ANTENNA_447 (.DIODE(net1502));
 sky130_fd_sc_hd__diode_2 ANTENNA_448 (.DIODE(net1502));
 sky130_fd_sc_hd__diode_2 ANTENNA_449 (.DIODE(net1506));
 sky130_fd_sc_hd__diode_2 ANTENNA_450 (.DIODE(net1506));
 sky130_fd_sc_hd__diode_2 ANTENNA_451 (.DIODE(net1518));
 sky130_fd_sc_hd__diode_2 ANTENNA_452 (.DIODE(net1563));
 sky130_fd_sc_hd__diode_2 ANTENNA_453 (.DIODE(net1563));
 sky130_fd_sc_hd__diode_2 ANTENNA_454 (.DIODE(net1563));
 sky130_fd_sc_hd__diode_2 ANTENNA_455 (.DIODE(net1588));
 sky130_fd_sc_hd__diode_2 ANTENNA_456 (.DIODE(net1614));
 sky130_fd_sc_hd__diode_2 ANTENNA_457 (.DIODE(net1619));
 sky130_fd_sc_hd__diode_2 ANTENNA_458 (.DIODE(net1640));
 sky130_fd_sc_hd__diode_2 ANTENNA_459 (.DIODE(net1640));
 sky130_fd_sc_hd__diode_2 ANTENNA_460 (.DIODE(net1674));
 sky130_fd_sc_hd__diode_2 ANTENNA_461 (.DIODE(net1683));
 sky130_fd_sc_hd__diode_2 ANTENNA_462 (.DIODE(net1706));
 sky130_fd_sc_hd__diode_2 ANTENNA_463 (.DIODE(net1751));
 sky130_fd_sc_hd__diode_2 ANTENNA_464 (.DIODE(net1752));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_843 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1092 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1151 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1095 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1122 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1064 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_927 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1095 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1148 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1092 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_843 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1161 ();
endmodule

