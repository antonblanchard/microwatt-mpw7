* NGSPICE file created from Microwatt_FP_DFFRFile.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

.subckt Microwatt_FP_DFFRFile CLK D1[0] D1[10] D1[11] D1[12] D1[13] D1[14] D1[15]
+ D1[16] D1[17] D1[18] D1[19] D1[1] D1[20] D1[21] D1[22] D1[23] D1[24] D1[25] D1[26]
+ D1[27] D1[28] D1[29] D1[2] D1[30] D1[31] D1[32] D1[33] D1[34] D1[35] D1[36] D1[37]
+ D1[38] D1[39] D1[3] D1[40] D1[41] D1[42] D1[43] D1[44] D1[45] D1[46] D1[47] D1[48]
+ D1[49] D1[4] D1[50] D1[51] D1[52] D1[53] D1[54] D1[55] D1[56] D1[57] D1[58] D1[59]
+ D1[5] D1[60] D1[61] D1[62] D1[63] D1[6] D1[7] D1[8] D1[9] D2[0] D2[10] D2[11] D2[12]
+ D2[13] D2[14] D2[15] D2[16] D2[17] D2[18] D2[19] D2[1] D2[20] D2[21] D2[22] D2[23]
+ D2[24] D2[25] D2[26] D2[27] D2[28] D2[29] D2[2] D2[30] D2[31] D2[32] D2[33] D2[34]
+ D2[35] D2[36] D2[37] D2[38] D2[39] D2[3] D2[40] D2[41] D2[42] D2[43] D2[44] D2[45]
+ D2[46] D2[47] D2[48] D2[49] D2[4] D2[50] D2[51] D2[52] D2[53] D2[54] D2[55] D2[56]
+ D2[57] D2[58] D2[59] D2[5] D2[60] D2[61] D2[62] D2[63] D2[6] D2[7] D2[8] D2[9] D3[0]
+ D3[10] D3[11] D3[12] D3[13] D3[14] D3[15] D3[16] D3[17] D3[18] D3[19] D3[1] D3[20]
+ D3[21] D3[22] D3[23] D3[24] D3[25] D3[26] D3[27] D3[28] D3[29] D3[2] D3[30] D3[31]
+ D3[32] D3[33] D3[34] D3[35] D3[36] D3[37] D3[38] D3[39] D3[3] D3[40] D3[41] D3[42]
+ D3[43] D3[44] D3[45] D3[46] D3[47] D3[48] D3[49] D3[4] D3[50] D3[51] D3[52] D3[53]
+ D3[54] D3[55] D3[56] D3[57] D3[58] D3[59] D3[5] D3[60] D3[61] D3[62] D3[63] D3[6]
+ D3[7] D3[8] D3[9] DW[0] DW[10] DW[11] DW[12] DW[13] DW[14] DW[15] DW[16] DW[17]
+ DW[18] DW[19] DW[1] DW[20] DW[21] DW[22] DW[23] DW[24] DW[25] DW[26] DW[27] DW[28]
+ DW[29] DW[2] DW[30] DW[31] DW[32] DW[33] DW[34] DW[35] DW[36] DW[37] DW[38] DW[39]
+ DW[3] DW[40] DW[41] DW[42] DW[43] DW[44] DW[45] DW[46] DW[47] DW[48] DW[49] DW[4]
+ DW[50] DW[51] DW[52] DW[53] DW[54] DW[55] DW[56] DW[57] DW[58] DW[59] DW[5] DW[60]
+ DW[61] DW[62] DW[63] DW[6] DW[7] DW[8] DW[9] R1[0] R1[1] R1[2] R1[3] R1[4] R1[5]
+ R2[0] R2[1] R2[2] R2[3] R2[4] R2[5] R3[0] R3[1] R3[2] R3[3] R3[4] R3[5] RW[0] RW[1]
+ RW[2] RW[3] RW[4] RW[5] VGND VPWR WE
XFILLER_228_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34984_ _34987_/CLK _34984_/D VGND VGND VPWR VPWR _34984_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1360 _23105_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1371 _24407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1382 _28776_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33935_ _34262_/CLK _33935_/D VGND VGND VPWR VPWR _33935_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1393 _16623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18869_ _18649_/X _18867_/X _18868_/X _18655_/X VGND VGND VPWR VPWR _18869_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20900_ _22312_/A VGND VGND VPWR VPWR _20900_/X sky130_fd_sc_hd__buf_6
X_21880_ _21875_/X _21879_/X _21736_/X _21737_/X VGND VGND VPWR VPWR _21897_/B sky130_fd_sc_hd__o211a_1
X_33866_ _35852_/CLK _33866_/D VGND VGND VPWR VPWR _33866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20831_ _34770_/Q _34706_/Q _34642_/Q _34578_/Q _20829_/X _20830_/X VGND VGND VPWR
+ VPWR _20831_/X sky130_fd_sc_hd__mux4_1
X_35605_ _35669_/CLK _35605_/D VGND VGND VPWR VPWR _35605_/Q sky130_fd_sc_hd__dfxtp_1
X_32817_ _33009_/CLK _32817_/D VGND VGND VPWR VPWR _32817_/Q sky130_fd_sc_hd__dfxtp_1
X_33797_ _34309_/CLK _33797_/D VGND VGND VPWR VPWR _33797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23550_ _23550_/A VGND VGND VPWR VPWR _32328_/D sky130_fd_sc_hd__clkbuf_1
X_20762_ _20758_/X _20761_/X _20671_/X VGND VGND VPWR VPWR _20772_/C sky130_fd_sc_hd__o21ba_1
X_35536_ _35793_/CLK _35536_/D VGND VGND VPWR VPWR _35536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32748_ _36076_/CLK _32748_/D VGND VGND VPWR VPWR _32748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22501_ _22501_/A VGND VGND VPWR VPWR _22501_/X sky130_fd_sc_hd__buf_4
XFILLER_168_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23481_ _23481_/A VGND VGND VPWR VPWR _32295_/D sky130_fd_sc_hd__clkbuf_1
X_35467_ _35978_/CLK _35467_/D VGND VGND VPWR VPWR _35467_/Q sky130_fd_sc_hd__dfxtp_1
X_32679_ _33255_/CLK _32679_/D VGND VGND VPWR VPWR _32679_/Q sky130_fd_sc_hd__dfxtp_1
X_20693_ _22370_/A VGND VGND VPWR VPWR _21757_/A sky130_fd_sc_hd__buf_12
X_22432_ _34048_/Q _33984_/Q _33920_/Q _32256_/Q _22326_/X _22327_/X VGND VGND VPWR
+ VPWR _22432_/X sky130_fd_sc_hd__mux4_1
X_25220_ _25035_/X _33052_/Q _25230_/S VGND VGND VPWR VPWR _25221_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34418_ _34866_/CLK _34418_/D VGND VGND VPWR VPWR _34418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35398_ _35975_/CLK _35398_/D VGND VGND VPWR VPWR _35398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25151_ _25150_/X _33025_/Q _25175_/S VGND VGND VPWR VPWR _25152_/A sky130_fd_sc_hd__mux2_1
X_22363_ _32766_/Q _32702_/Q _32638_/Q _36094_/Q _22225_/X _22362_/X VGND VGND VPWR
+ VPWR _22363_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34349_ _35307_/CLK _34349_/D VGND VGND VPWR VPWR _34349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24102_ _23068_/X _32587_/Q _24106_/S VGND VGND VPWR VPWR _24103_/A sky130_fd_sc_hd__mux2_1
X_21314_ _22511_/A VGND VGND VPWR VPWR _21314_/X sky130_fd_sc_hd__clkbuf_4
X_25082_ _25081_/X _33003_/Q _25082_/S VGND VGND VPWR VPWR _25083_/A sky130_fd_sc_hd__mux2_1
X_22294_ _32508_/Q _32380_/Q _32060_/Q _36028_/Q _22229_/X _22017_/X VGND VGND VPWR
+ VPWR _22294_/X sky130_fd_sc_hd__mux4_1
XFILLER_102_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28910_ _28910_/A VGND VGND VPWR VPWR _34764_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24033_ _22966_/X _32554_/Q _24035_/S VGND VGND VPWR VPWR _24034_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21245_ _21241_/X _21242_/X _21243_/X _21244_/X VGND VGND VPWR VPWR _21245_/X sky130_fd_sc_hd__a22o_1
X_36019_ _36019_/CLK _36019_/D VGND VGND VPWR VPWR _36019_/Q sky130_fd_sc_hd__dfxtp_1
X_29890_ _29890_/A VGND VGND VPWR VPWR _35197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28841_ _28841_/A VGND VGND VPWR VPWR _34731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21176_ _35740_/Q _35100_/Q _34460_/Q _33820_/Q _21034_/X _21035_/X VGND VGND VPWR
+ VPWR _21176_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20127_ _34304_/Q _34240_/Q _34176_/Q _34112_/Q _20095_/X _20096_/X VGND VGND VPWR
+ VPWR _20127_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28772_ _27011_/X _34699_/Q _28776_/S VGND VGND VPWR VPWR _28773_/A sky130_fd_sc_hd__mux2_1
X_25984_ _25984_/A VGND VGND VPWR VPWR _33409_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27723_ _34201_/Q _24280_/X _27739_/S VGND VGND VPWR VPWR _27724_/A sky130_fd_sc_hd__mux2_1
X_20058_ _34046_/Q _33982_/Q _33918_/Q _32254_/Q _20026_/X _20027_/X VGND VGND VPWR
+ VPWR _20058_/X sky130_fd_sc_hd__mux4_1
X_24935_ _22997_/X _32948_/Q _24937_/S VGND VGND VPWR VPWR _24936_/A sky130_fd_sc_hd__mux2_1
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27654_ _27654_/A VGND VGND VPWR VPWR _34168_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24866_ _22895_/X _32915_/Q _24874_/S VGND VGND VPWR VPWR _24867_/A sky130_fd_sc_hd__mux2_1
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_202 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26605_ _26605_/A VGND VGND VPWR VPWR _33703_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_213 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23817_ _23817_/A VGND VGND VPWR VPWR _32452_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_224 _32136_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27585_ _27696_/S VGND VGND VPWR VPWR _27604_/S sky130_fd_sc_hd__buf_4
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_235 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24797_ _24797_/A VGND VGND VPWR VPWR _32882_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_246 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_257 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29324_ _23253_/X _34929_/Q _29332_/S VGND VGND VPWR VPWR _29325_/A sky130_fd_sc_hd__mux2_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26536_ _26536_/A VGND VGND VPWR VPWR _33671_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_268 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23748_ _23748_/A VGND VGND VPWR VPWR _32419_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_279 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29255_ _23093_/X _34896_/Q _29269_/S VGND VGND VPWR VPWR _29256_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26467_ _26467_/A VGND VGND VPWR VPWR _33638_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23679_ _23679_/A VGND VGND VPWR VPWR _32388_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28206_ _28206_/A VGND VGND VPWR VPWR _34430_/D sky130_fd_sc_hd__clkbuf_1
X_16220_ _16026_/X _16218_/X _16219_/X _16037_/X VGND VGND VPWR VPWR _16220_/X sky130_fd_sc_hd__a22o_1
X_25418_ _25418_/A VGND VGND VPWR VPWR _33145_/D sky130_fd_sc_hd__clkbuf_1
X_29186_ _34873_/Q _29185_/X _29204_/S VGND VGND VPWR VPWR _29187_/A sky130_fd_sc_hd__mux2_1
X_26398_ _25165_/X _33606_/Q _26404_/S VGND VGND VPWR VPWR _26399_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16151_ _16014_/X _16149_/X _16150_/X _16023_/X VGND VGND VPWR VPWR _16151_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28137_ _28137_/A VGND VGND VPWR VPWR _34397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25349_ _25349_/A VGND VGND VPWR VPWR _33112_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_867 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16082_ _35278_/Q _35214_/Q _35150_/Q _32270_/Q _16079_/X _16081_/X VGND VGND VPWR
+ VPWR _16082_/X sky130_fd_sc_hd__mux4_1
X_28068_ _26968_/X _34365_/Q _28072_/S VGND VGND VPWR VPWR _28069_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27019_ _27019_/A VGND VGND VPWR VPWR _33869_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19910_ _35321_/Q _35257_/Q _35193_/Q _32313_/Q _19659_/X _19660_/X VGND VGND VPWR
+ VPWR _19910_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30030_ _30057_/S VGND VGND VPWR VPWR _30049_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_194_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19841_ _19802_/X _19839_/X _19840_/X _19805_/X VGND VGND VPWR VPWR _19841_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19772_ _19772_/A VGND VGND VPWR VPWR _32117_/D sky130_fd_sc_hd__buf_2
XFILLER_96_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16984_ _16980_/X _16983_/X _16775_/X VGND VGND VPWR VPWR _17014_/A sky130_fd_sc_hd__o21ba_1
XFILLER_122_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18723_ _18716_/X _18721_/X _18722_/X VGND VGND VPWR VPWR _18757_/A sky130_fd_sc_hd__o21ba_1
XTAP_5160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31981_ _35166_/CLK _31981_/D VGND VGND VPWR VPWR _31981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18654_ _33238_/Q _36118_/Q _33110_/Q _33046_/Q _18652_/X _18653_/X VGND VGND VPWR
+ VPWR _18654_/X sky130_fd_sc_hd__mux4_1
X_33720_ _34297_/CLK _33720_/D VGND VGND VPWR VPWR _33720_/Q sky130_fd_sc_hd__dfxtp_1
X_30932_ _35691_/Q _29141_/X _30932_/S VGND VGND VPWR VPWR _30933_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _35034_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17605_ _35577_/Q _35513_/Q _35449_/Q _35385_/Q _17603_/X _17604_/X VGND VGND VPWR
+ VPWR _17605_/X sky130_fd_sc_hd__mux4_2
XFILLER_91_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30863_ _30863_/A VGND VGND VPWR VPWR _35658_/D sky130_fd_sc_hd__clkbuf_1
X_18585_ _32980_/Q _32916_/Q _32852_/Q _32788_/Q _18583_/X _18584_/X VGND VGND VPWR
+ VPWR _18585_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33651_ _34227_/CLK _33651_/D VGND VGND VPWR VPWR _33651_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17536_ _33207_/Q _32567_/Q _35959_/Q _35895_/Q _17427_/X _17428_/X VGND VGND VPWR
+ VPWR _17536_/X sky130_fd_sc_hd__mux4_1
X_32602_ _32666_/CLK _32602_/D VGND VGND VPWR VPWR _32602_/Q sky130_fd_sc_hd__dfxtp_1
X_33582_ _34288_/CLK _33582_/D VGND VGND VPWR VPWR _33582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30794_ _30794_/A VGND VGND VPWR VPWR _35625_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_780 _22604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_791 _22693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32533_ _35925_/CLK _32533_/D VGND VGND VPWR VPWR _32533_/Q sky130_fd_sc_hd__dfxtp_1
X_35321_ _35577_/CLK _35321_/D VGND VGND VPWR VPWR _35321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17467_ _34549_/Q _32437_/Q _34421_/Q _34357_/Q _17225_/X _17226_/X VGND VGND VPWR
+ VPWR _17467_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16418_ _17796_/A VGND VGND VPWR VPWR _16418_/X sky130_fd_sc_hd__buf_4
X_19206_ _34533_/Q _32421_/Q _34405_/Q _34341_/Q _19172_/X _19173_/X VGND VGND VPWR
+ VPWR _19206_/X sky130_fd_sc_hd__mux4_1
X_32464_ _36049_/CLK _32464_/D VGND VGND VPWR VPWR _32464_/Q sky130_fd_sc_hd__dfxtp_1
X_35252_ _35252_/CLK _35252_/D VGND VGND VPWR VPWR _35252_/Q sky130_fd_sc_hd__dfxtp_1
X_17398_ _17394_/X _17397_/X _17161_/X VGND VGND VPWR VPWR _17399_/D sky130_fd_sc_hd__o21ba_1
XFILLER_158_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31415_ _31415_/A VGND VGND VPWR VPWR _35919_/D sky130_fd_sc_hd__clkbuf_1
X_34203_ _34267_/CLK _34203_/D VGND VGND VPWR VPWR _34203_/Q sky130_fd_sc_hd__dfxtp_1
X_19137_ _35043_/Q _34979_/Q _34915_/Q _34851_/Q _19103_/X _19104_/X VGND VGND VPWR
+ VPWR _19137_/X sky130_fd_sc_hd__mux4_1
X_16349_ _17901_/A VGND VGND VPWR VPWR _16349_/X sky130_fd_sc_hd__clkbuf_4
X_35183_ _35564_/CLK _35183_/D VGND VGND VPWR VPWR _35183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32395_ _36172_/CLK _32395_/D VGND VGND VPWR VPWR _32395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34134_ _34197_/CLK _34134_/D VGND VGND VPWR VPWR _34134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31346_ _35887_/Q input27/X _31358_/S VGND VGND VPWR VPWR _31347_/A sky130_fd_sc_hd__mux2_1
X_19068_ _34274_/Q _34210_/Q _34146_/Q _34082_/Q _19036_/X _19037_/X VGND VGND VPWR
+ VPWR _19068_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18019_ _35845_/Q _32224_/Q _35717_/Q _35653_/Q _15989_/X _15991_/X VGND VGND VPWR
+ VPWR _18019_/X sky130_fd_sc_hd__mux4_1
X_34065_ _34262_/CLK _34065_/D VGND VGND VPWR VPWR _34065_/Q sky130_fd_sc_hd__dfxtp_1
X_31277_ _35854_/Q input1/X _31295_/S VGND VGND VPWR VPWR _31278_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33016_ _36089_/CLK _33016_/D VGND VGND VPWR VPWR _33016_/Q sky130_fd_sc_hd__dfxtp_1
X_21030_ _22442_/A VGND VGND VPWR VPWR _21030_/X sky130_fd_sc_hd__clkbuf_4
X_30228_ _30228_/A VGND VGND VPWR VPWR _35357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30159_ _35325_/Q _29197_/X _30163_/S VGND VGND VPWR VPWR _30160_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34967_ _34967_/CLK _34967_/D VGND VGND VPWR VPWR _34967_/Q sky130_fd_sc_hd__dfxtp_1
X_22981_ _22981_/A VGND VGND VPWR VPWR _32046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1190 _23075_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24720_ _24852_/S VGND VGND VPWR VPWR _24739_/S sky130_fd_sc_hd__buf_4
XFILLER_83_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33918_ _34046_/CLK _33918_/D VGND VGND VPWR VPWR _33918_/Q sky130_fd_sc_hd__dfxtp_1
X_21932_ _34290_/Q _34226_/Q _34162_/Q _34098_/Q _21689_/X _21690_/X VGND VGND VPWR
+ VPWR _21932_/X sky130_fd_sc_hd__mux4_1
XFILLER_243_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34898_ _35026_/CLK _34898_/D VGND VGND VPWR VPWR _34898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24651_ _22979_/X _32814_/Q _24665_/S VGND VGND VPWR VPWR _24652_/A sky130_fd_sc_hd__mux2_1
X_33849_ _35771_/CLK _33849_/D VGND VGND VPWR VPWR _33849_/Q sky130_fd_sc_hd__dfxtp_1
X_21863_ _21863_/A _21863_/B _21863_/C _21863_/D VGND VGND VPWR VPWR _21864_/A sky130_fd_sc_hd__or4_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23602_ _32352_/Q _23142_/X _23604_/S VGND VGND VPWR VPWR _23603_/A sky130_fd_sc_hd__mux2_1
XFILLER_247_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20814_ _32722_/Q _32658_/Q _32594_/Q _36050_/Q _20813_/X _22313_/A VGND VGND VPWR
+ VPWR _20814_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27370_ _34035_/Q _24360_/X _27374_/S VGND VGND VPWR VPWR _27371_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24582_ _27968_/A _31815_/B VGND VGND VPWR VPWR _24715_/S sky130_fd_sc_hd__nand2_8
X_21794_ _21794_/A VGND VGND VPWR VPWR _36205_/D sky130_fd_sc_hd__buf_6
XFILLER_93_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26321_ _26321_/A VGND VGND VPWR VPWR _33569_/D sky130_fd_sc_hd__clkbuf_1
X_23533_ _23034_/X _32320_/Q _23551_/S VGND VGND VPWR VPWR _23534_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35519_ _35583_/CLK _35519_/D VGND VGND VPWR VPWR _35519_/Q sky130_fd_sc_hd__dfxtp_1
X_20745_ _34000_/Q _33936_/Q _33872_/Q _32144_/Q _20708_/X _20709_/X VGND VGND VPWR
+ VPWR _20745_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29040_ _34826_/Q _24431_/X _29046_/S VGND VGND VPWR VPWR _29041_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26252_ _26252_/A VGND VGND VPWR VPWR _33536_/D sky130_fd_sc_hd__clkbuf_1
X_20676_ _22532_/A VGND VGND VPWR VPWR _20676_/X sky130_fd_sc_hd__buf_4
X_23464_ _23464_/A VGND VGND VPWR VPWR _32287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25203_ _25010_/X _33044_/Q _25209_/S VGND VGND VPWR VPWR _25204_/A sky130_fd_sc_hd__mux2_1
X_22415_ _22305_/X _22413_/X _22414_/X _22308_/X VGND VGND VPWR VPWR _22415_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26183_ _25047_/X _33504_/Q _26185_/S VGND VGND VPWR VPWR _26184_/A sky130_fd_sc_hd__mux2_1
X_23395_ _32256_/Q _23303_/X _23413_/S VGND VGND VPWR VPWR _23396_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25134_ input41/X VGND VGND VPWR VPWR _25134_/X sky130_fd_sc_hd__buf_2
XFILLER_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22346_ _35325_/Q _35261_/Q _35197_/Q _32317_/Q _22312_/X _22313_/X VGND VGND VPWR
+ VPWR _22346_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29942_ _35222_/Q _29076_/X _29944_/S VGND VGND VPWR VPWR _29943_/A sky130_fd_sc_hd__mux2_1
X_22277_ _22102_/X _22275_/X _22276_/X _22105_/X VGND VGND VPWR VPWR _22277_/X sky130_fd_sc_hd__a22o_1
X_25065_ _25065_/A VGND VGND VPWR VPWR _32997_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24016_ _24106_/S VGND VGND VPWR VPWR _24035_/S sky130_fd_sc_hd__buf_4
X_21228_ _33502_/Q _33438_/Q _33374_/Q _33310_/Q _21017_/X _21018_/X VGND VGND VPWR
+ VPWR _21228_/X sky130_fd_sc_hd__mux4_1
X_29873_ _29873_/A VGND VGND VPWR VPWR _35189_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28824_ _26888_/X _34723_/Q _28840_/S VGND VGND VPWR VPWR _28825_/A sky130_fd_sc_hd__mux2_1
X_21159_ _33756_/Q _33692_/Q _33628_/Q _33564_/Q _21090_/X _21091_/X VGND VGND VPWR
+ VPWR _21159_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28755_ _28755_/A VGND VGND VPWR VPWR _34690_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25967_ _25967_/A VGND VGND VPWR VPWR _33401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27706_ _34193_/Q _24255_/X _27718_/S VGND VGND VPWR VPWR _27707_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24918_ _24987_/S VGND VGND VPWR VPWR _24937_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_18_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28686_ _28776_/S VGND VGND VPWR VPWR _28705_/S sky130_fd_sc_hd__buf_4
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25898_ _25898_/A VGND VGND VPWR VPWR _33368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27637_ _27637_/A VGND VGND VPWR VPWR _34160_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24849_ _24849_/A VGND VGND VPWR VPWR _32907_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ input81/X input82/X VGND VGND VPWR VPWR _20153_/A sky130_fd_sc_hd__or2_4
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27568_ _27568_/A VGND VGND VPWR VPWR _34127_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _17317_/X _17320_/X _17147_/X VGND VGND VPWR VPWR _17329_/C sky130_fd_sc_hd__o21ba_1
X_29307_ _23228_/X _34921_/Q _29311_/S VGND VGND VPWR VPWR _29308_/A sky130_fd_sc_hd__mux2_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26519_ _26519_/A VGND VGND VPWR VPWR _33663_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27499_ _26928_/X _34096_/Q _27509_/S VGND VGND VPWR VPWR _27500_/A sky130_fd_sc_hd__mux2_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1056 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29238_ _34890_/Q _29237_/X _29247_/S VGND VGND VPWR VPWR _29239_/A sky130_fd_sc_hd__mux2_1
X_17252_ _35567_/Q _35503_/Q _35439_/Q _35375_/Q _17250_/X _17251_/X VGND VGND VPWR
+ VPWR _17252_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16203_ _16199_/X _16202_/X _16100_/X VGND VGND VPWR VPWR _16204_/D sky130_fd_sc_hd__o21ba_1
XFILLER_168_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17183_ _33197_/Q _32557_/Q _35949_/Q _35885_/Q _17074_/X _17075_/X VGND VGND VPWR
+ VPWR _17183_/X sky130_fd_sc_hd__mux4_1
X_29169_ input32/X VGND VGND VPWR VPWR _29169_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_127_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31200_ _35818_/Q input21/X _31202_/S VGND VGND VPWR VPWR _31201_/A sky130_fd_sc_hd__mux2_1
X_16134_ _16134_/A _16134_/B _16134_/C _16134_/D VGND VGND VPWR VPWR _16135_/A sky130_fd_sc_hd__or4_4
XFILLER_183_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32180_ _35744_/CLK _32180_/D VGND VGND VPWR VPWR _32180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31131_ _31131_/A VGND VGND VPWR VPWR _35785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16065_ _17932_/A VGND VGND VPWR VPWR _16065_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_185_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31062_ _31062_/A VGND VGND VPWR VPWR _35752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30013_ _30013_/A VGND VGND VPWR VPWR _35255_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19824_ _19820_/X _19823_/X _19781_/X VGND VGND VPWR VPWR _19846_/A sky130_fd_sc_hd__o21ba_1
X_35870_ _35935_/CLK _35870_/D VGND VGND VPWR VPWR _35870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34821_ _35333_/CLK _34821_/D VGND VGND VPWR VPWR _34821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19755_ _19716_/X _19753_/X _19754_/X _19720_/X VGND VGND VPWR VPWR _19755_/X sky130_fd_sc_hd__a22o_1
XFILLER_110_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16967_ _16646_/X _16965_/X _16966_/X _16649_/X VGND VGND VPWR VPWR _16967_/X sky130_fd_sc_hd__a22o_1
X_18706_ _35287_/Q _35223_/Q _35159_/Q _32279_/Q _18600_/X _18601_/X VGND VGND VPWR
+ VPWR _18706_/X sky130_fd_sc_hd__mux4_1
X_34752_ _34752_/CLK _34752_/D VGND VGND VPWR VPWR _34752_/Q sky130_fd_sc_hd__dfxtp_1
X_31964_ _35166_/CLK _31964_/D VGND VGND VPWR VPWR _31964_/Q sky130_fd_sc_hd__dfxtp_1
X_16898_ _17957_/A VGND VGND VPWR VPWR _16898_/X sky130_fd_sc_hd__buf_4
X_19686_ _35763_/Q _35123_/Q _34483_/Q _33843_/Q _19440_/X _19441_/X VGND VGND VPWR
+ VPWR _19686_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33703_ _34278_/CLK _33703_/D VGND VGND VPWR VPWR _33703_/Q sky130_fd_sc_hd__dfxtp_1
X_18637_ _35029_/Q _34965_/Q _34901_/Q _34837_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _18637_/X sky130_fd_sc_hd__mux4_1
X_30915_ _30915_/A VGND VGND VPWR VPWR _35682_/D sky130_fd_sc_hd__clkbuf_1
X_34683_ _34811_/CLK _34683_/D VGND VGND VPWR VPWR _34683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31895_ _31895_/A VGND VGND VPWR VPWR _36147_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30846_ _23310_/X _35650_/Q _30860_/S VGND VGND VPWR VPWR _30847_/A sky130_fd_sc_hd__mux2_1
X_33634_ _33635_/CLK _33634_/D VGND VGND VPWR VPWR _33634_/Q sky130_fd_sc_hd__dfxtp_1
X_18568_ _18387_/X _18566_/X _18567_/X _18397_/X VGND VGND VPWR VPWR _18568_/X sky130_fd_sc_hd__a22o_1
XFILLER_240_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17519_ _34295_/Q _34231_/Q _34167_/Q _34103_/Q _17442_/X _17443_/X VGND VGND VPWR
+ VPWR _17519_/X sky130_fd_sc_hd__mux4_1
X_18499_ _18374_/X _18497_/X _18498_/X _18384_/X VGND VGND VPWR VPWR _18499_/X sky130_fd_sc_hd__a22o_1
X_30777_ _30777_/A VGND VGND VPWR VPWR _35617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33565_ _34010_/CLK _33565_/D VGND VGND VPWR VPWR _33565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20530_ _35788_/Q _35148_/Q _34508_/Q _33868_/Q _18408_/X _18409_/X VGND VGND VPWR
+ VPWR _20530_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_1156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35304_ _35304_/CLK _35304_/D VGND VGND VPWR VPWR _35304_/Q sky130_fd_sc_hd__dfxtp_1
X_32516_ _32901_/CLK _32516_/D VGND VGND VPWR VPWR _32516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33496_ _34267_/CLK _33496_/D VGND VGND VPWR VPWR _33496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20461_ _20457_/X _20460_/X _20134_/A VGND VGND VPWR VPWR _20483_/A sky130_fd_sc_hd__o21ba_1
X_32447_ _35966_/CLK _32447_/D VGND VGND VPWR VPWR _32447_/Q sky130_fd_sc_hd__dfxtp_1
X_35235_ _35299_/CLK _35235_/D VGND VGND VPWR VPWR _35235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22200_ _35833_/Q _32211_/Q _35705_/Q _35641_/Q _21913_/X _21914_/X VGND VGND VPWR
+ VPWR _22200_/X sky130_fd_sc_hd__mux4_1
X_23180_ _32173_/Q _23111_/X _23182_/S VGND VGND VPWR VPWR _23181_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20392_ _20388_/X _20391_/X _20167_/X VGND VGND VPWR VPWR _20393_/D sky130_fd_sc_hd__o21ba_1
XFILLER_238_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32378_ _36027_/CLK _32378_/D VGND VGND VPWR VPWR _32378_/Q sky130_fd_sc_hd__dfxtp_1
X_35166_ _35166_/CLK _35166_/D VGND VGND VPWR VPWR _35166_/Q sky130_fd_sc_hd__dfxtp_1
X_22131_ _22127_/X _22130_/X _22089_/X _22090_/X VGND VGND VPWR VPWR _22146_/B sky130_fd_sc_hd__o211a_1
X_34117_ _34308_/CLK _34117_/D VGND VGND VPWR VPWR _34117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31329_ _35879_/Q input18/X _31337_/S VGND VGND VPWR VPWR _31330_/A sky130_fd_sc_hd__mux2_1
X_35097_ _35929_/CLK _35097_/D VGND VGND VPWR VPWR _35097_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput220 _32089_/Q VGND VGND VPWR VPWR D3[11] sky130_fd_sc_hd__buf_2
Xoutput231 _32099_/Q VGND VGND VPWR VPWR D3[21] sky130_fd_sc_hd__buf_2
XFILLER_161_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput242 _32109_/Q VGND VGND VPWR VPWR D3[31] sky130_fd_sc_hd__buf_2
XFILLER_82_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput253 _32119_/Q VGND VGND VPWR VPWR D3[41] sky130_fd_sc_hd__buf_2
X_22062_ _21952_/X _22060_/X _22061_/X _21955_/X VGND VGND VPWR VPWR _22062_/X sky130_fd_sc_hd__a22o_1
XTAP_6619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34048_ _34050_/CLK _34048_/D VGND VGND VPWR VPWR _34048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput264 _32129_/Q VGND VGND VPWR VPWR D3[51] sky130_fd_sc_hd__buf_2
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput275 _32139_/Q VGND VGND VPWR VPWR D3[61] sky130_fd_sc_hd__buf_2
Xclkbuf_6_3__f_CLK clkbuf_5_1_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_3__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_248_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21013_ _21013_/A VGND VGND VPWR VPWR _36183_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26870_ _26869_/X _33821_/Q _26882_/S VGND VGND VPWR VPWR _26871_/A sky130_fd_sc_hd__mux2_1
XTAP_5929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25821_ _25821_/A VGND VGND VPWR VPWR _33332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35999_ _36125_/CLK _35999_/D VGND VGND VPWR VPWR _35999_/Q sky130_fd_sc_hd__dfxtp_1
X_28540_ _28540_/A VGND VGND VPWR VPWR _34588_/D sky130_fd_sc_hd__clkbuf_1
X_25752_ _25752_/A VGND VGND VPWR VPWR _33299_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22964_ _22963_/X _32041_/Q _22970_/S VGND VGND VPWR VPWR _22965_/A sky130_fd_sc_hd__mux2_1
X_24703_ _23056_/X _32839_/Q _24707_/S VGND VGND VPWR VPWR _24704_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28471_ _26965_/X _34556_/Q _28477_/S VGND VGND VPWR VPWR _28472_/A sky130_fd_sc_hd__mux2_1
X_21915_ _35825_/Q _32202_/Q _35697_/Q _35633_/Q _21913_/X _21914_/X VGND VGND VPWR
+ VPWR _21915_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25683_ _33268_/Q _24363_/X _25685_/S VGND VGND VPWR VPWR _25684_/A sky130_fd_sc_hd__mux2_1
X_22895_ input56/X VGND VGND VPWR VPWR _22895_/X sky130_fd_sc_hd__buf_4
XFILLER_15_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27422_ _34060_/Q _24437_/X _27424_/S VGND VGND VPWR VPWR _27423_/A sky130_fd_sc_hd__mux2_1
X_24634_ _22954_/X _32806_/Q _24644_/S VGND VGND VPWR VPWR _24635_/A sky130_fd_sc_hd__mux2_1
X_21846_ _21842_/X _21845_/X _21736_/X _21737_/X VGND VGND VPWR VPWR _21863_/B sky130_fd_sc_hd__o211a_1
XFILLER_231_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27353_ _34027_/Q _24335_/X _27353_/S VGND VGND VPWR VPWR _27354_/A sky130_fd_sc_hd__mux2_1
X_24565_ _23056_/X _32775_/Q _24569_/S VGND VGND VPWR VPWR _24566_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21777_ _21663_/X _21775_/X _21776_/X _21667_/X VGND VGND VPWR VPWR _21777_/X sky130_fd_sc_hd__a22o_1
XFILLER_211_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26304_ _25026_/X _33561_/Q _26320_/S VGND VGND VPWR VPWR _26305_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_1248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23516_ _23010_/X _32312_/Q _23530_/S VGND VGND VPWR VPWR _23517_/A sky130_fd_sc_hd__mux2_1
X_27284_ _27284_/A VGND VGND VPWR VPWR _33994_/D sky130_fd_sc_hd__clkbuf_1
X_20728_ _35279_/Q _35215_/Q _35151_/Q _32271_/Q _20679_/X _20681_/X VGND VGND VPWR
+ VPWR _20728_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24496_ _22954_/X _32742_/Q _24506_/S VGND VGND VPWR VPWR _24497_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29023_ _29023_/A VGND VGND VPWR VPWR _34817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26235_ _26235_/A VGND VGND VPWR VPWR _33528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23447_ _23447_/A VGND VGND VPWR VPWR _32279_/D sky130_fd_sc_hd__clkbuf_1
X_20659_ _20659_/A VGND VGND VPWR VPWR _22447_/A sky130_fd_sc_hd__buf_12
XFILLER_221_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26166_ _26277_/S VGND VGND VPWR VPWR _26185_/S sky130_fd_sc_hd__buf_4
XFILLER_104_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23378_ _32248_/Q _23277_/X _23392_/S VGND VGND VPWR VPWR _23379_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25117_ _25115_/X _33014_/Q _25144_/S VGND VGND VPWR VPWR _25118_/A sky130_fd_sc_hd__mux2_1
X_22329_ _22155_/X _22325_/X _22328_/X _22158_/X VGND VGND VPWR VPWR _22329_/X sky130_fd_sc_hd__a22o_1
XFILLER_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26097_ _25119_/X _33463_/Q _26113_/S VGND VGND VPWR VPWR _26098_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_1147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29925_ _30057_/S VGND VGND VPWR VPWR _29944_/S sky130_fd_sc_hd__buf_6
X_25048_ _25047_/X _32992_/Q _25051_/S VGND VGND VPWR VPWR _25049_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17870_ _17870_/A VGND VGND VPWR VPWR _32000_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_215_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29856_ _35181_/Q _29148_/X _29872_/S VGND VGND VPWR VPWR _29857_/A sky130_fd_sc_hd__mux2_1
X_28807_ _26863_/X _34715_/Q _28819_/S VGND VGND VPWR VPWR _28808_/A sky130_fd_sc_hd__mux2_1
X_16821_ _16702_/X _16819_/X _16820_/X _16708_/X VGND VGND VPWR VPWR _16821_/X sky130_fd_sc_hd__a22o_1
X_29787_ _35149_/Q _29246_/X _29787_/S VGND VGND VPWR VPWR _29788_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26999_ input53/X VGND VGND VPWR VPWR _26999_/X sky130_fd_sc_hd__buf_4
XFILLER_59_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19540_ _32751_/Q _32687_/Q _32623_/Q _36079_/Q _19219_/X _19356_/X VGND VGND VPWR
+ VPWR _19540_/X sky130_fd_sc_hd__mux4_1
X_16752_ _35745_/Q _35105_/Q _34465_/Q _33825_/Q _16434_/X _16435_/X VGND VGND VPWR
+ VPWR _16752_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28738_ _28738_/A VGND VGND VPWR VPWR _34682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16683_ _33183_/Q _32543_/Q _35935_/Q _35871_/Q _16368_/X _16369_/X VGND VGND VPWR
+ VPWR _16683_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28669_ _28669_/A VGND VGND VPWR VPWR _34649_/D sky130_fd_sc_hd__clkbuf_1
X_19471_ _19467_/X _19470_/X _19428_/X VGND VGND VPWR VPWR _19493_/A sky130_fd_sc_hd__o21ba_1
XFILLER_62_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30700_ _35581_/Q _29197_/X _30704_/S VGND VGND VPWR VPWR _30701_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18422_ _18344_/X _18420_/X _18421_/X _18354_/X VGND VGND VPWR VPWR _18422_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31680_ _31680_/A _31680_/B VGND VGND VPWR VPWR _31813_/S sky130_fd_sc_hd__nor2_8
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _20067_/A VGND VGND VPWR VPWR _20158_/A sky130_fd_sc_hd__buf_12
X_30631_ _35548_/Q _29095_/X _30641_/S VGND VGND VPWR VPWR _30632_/A sky130_fd_sc_hd__mux2_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_230_CLK clkbuf_6_60__f_CLK/X VGND VGND VPWR VPWR _32901_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _17202_/X _17302_/X _17303_/X _17205_/X VGND VGND VPWR VPWR _17304_/X sky130_fd_sc_hd__a22o_1
X_33350_ _34053_/CLK _33350_/D VGND VGND VPWR VPWR _33350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18284_ _33742_/Q _33678_/Q _33614_/Q _33550_/Q _18280_/X _18283_/X VGND VGND VPWR
+ VPWR _18284_/X sky130_fd_sc_hd__mux4_1
X_30562_ _30562_/A VGND VGND VPWR VPWR _35515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32301_ _35500_/CLK _32301_/D VGND VGND VPWR VPWR _32301_/Q sky130_fd_sc_hd__dfxtp_1
X_17235_ _17195_/X _17233_/X _17234_/X _17200_/X VGND VGND VPWR VPWR _17235_/X sky130_fd_sc_hd__a22o_1
X_33281_ _36161_/CLK _33281_/D VGND VGND VPWR VPWR _33281_/Q sky130_fd_sc_hd__dfxtp_1
X_30493_ _30493_/A VGND VGND VPWR VPWR _35482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35020_ _35277_/CLK _35020_/D VGND VGND VPWR VPWR _35020_/Q sky130_fd_sc_hd__dfxtp_1
X_32232_ _35853_/CLK _32232_/D VGND VGND VPWR VPWR _32232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17166_ _34285_/Q _34221_/Q _34157_/Q _34093_/Q _17089_/X _17090_/X VGND VGND VPWR
+ VPWR _17166_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16117_ _32975_/Q _32911_/Q _32847_/Q _32783_/Q _16033_/X _16035_/X VGND VGND VPWR
+ VPWR _16117_/X sky130_fd_sc_hd__mux4_1
XFILLER_115_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32163_ _36130_/CLK _32163_/D VGND VGND VPWR VPWR _32163_/Q sky130_fd_sc_hd__dfxtp_1
X_17097_ _32747_/Q _32683_/Q _32619_/Q _36075_/Q _16919_/X _17056_/X VGND VGND VPWR
+ VPWR _17097_/X sky130_fd_sc_hd__mux4_1
X_31114_ _35777_/Q _29210_/X _31130_/S VGND VGND VPWR VPWR _31115_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16048_ _17978_/A VGND VGND VPWR VPWR _17994_/A sky130_fd_sc_hd__buf_12
XFILLER_100_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32094_ _35807_/CLK _32094_/D VGND VGND VPWR VPWR _32094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_297_CLK clkbuf_6_51__f_CLK/X VGND VGND VPWR VPWR _35709_/CLK sky130_fd_sc_hd__clkbuf_16
X_35922_ _35922_/CLK _35922_/D VGND VGND VPWR VPWR _35922_/Q sky130_fd_sc_hd__dfxtp_1
X_31045_ _31045_/A VGND VGND VPWR VPWR _35744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19807_ _20160_/A VGND VGND VPWR VPWR _19807_/X sky130_fd_sc_hd__clkbuf_4
X_35853_ _35853_/CLK _35853_/D VGND VGND VPWR VPWR _35853_/Q sky130_fd_sc_hd__dfxtp_1
X_17999_ _34564_/Q _32452_/Q _34436_/Q _34372_/Q _17931_/X _17932_/X VGND VGND VPWR
+ VPWR _17999_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34804_ _35250_/CLK _34804_/D VGND VGND VPWR VPWR _34804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19738_ _19734_/X _19737_/X _19461_/X VGND VGND VPWR VPWR _19739_/D sky130_fd_sc_hd__o21ba_1
X_35784_ _35784_/CLK _35784_/D VGND VGND VPWR VPWR _35784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32996_ _36069_/CLK _32996_/D VGND VGND VPWR VPWR _32996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34735_ _34932_/CLK _34735_/D VGND VGND VPWR VPWR _34735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31947_ _31947_/A VGND VGND VPWR VPWR _36172_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19669_ _33779_/Q _33715_/Q _33651_/Q _33587_/Q _19496_/X _19497_/X VGND VGND VPWR
+ VPWR _19669_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21700_ _32491_/Q _32363_/Q _32043_/Q _36011_/Q _21523_/X _21664_/X VGND VGND VPWR
+ VPWR _21700_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22680_ _35783_/Q _35143_/Q _34503_/Q _33863_/Q _22446_/X _22447_/X VGND VGND VPWR
+ VPWR _22680_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34666_ _34794_/CLK _34666_/D VGND VGND VPWR VPWR _34666_/Q sky130_fd_sc_hd__dfxtp_1
X_31878_ _31878_/A VGND VGND VPWR VPWR _36139_/D sky130_fd_sc_hd__clkbuf_1
X_33617_ _34259_/CLK _33617_/D VGND VGND VPWR VPWR _33617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21631_ _21627_/X _21630_/X _21383_/X _21384_/X VGND VGND VPWR VPWR _21646_/B sky130_fd_sc_hd__o211a_1
X_30829_ _23283_/X _35642_/Q _30839_/S VGND VGND VPWR VPWR _30830_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34597_ _36001_/CLK _34597_/D VGND VGND VPWR VPWR _34597_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_221_CLK clkbuf_6_55__f_CLK/X VGND VGND VPWR VPWR _34947_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_221_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24350_ _24350_/A VGND VGND VPWR VPWR _32687_/D sky130_fd_sc_hd__clkbuf_1
X_33548_ _33548_/CLK _33548_/D VGND VGND VPWR VPWR _33548_/Q sky130_fd_sc_hd__dfxtp_1
X_21562_ _35815_/Q _32191_/Q _35687_/Q _35623_/Q _21560_/X _21561_/X VGND VGND VPWR
+ VPWR _21562_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23301_ _32218_/Q _23300_/X _23301_/S VGND VGND VPWR VPWR _23302_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20513_ _20513_/A _20513_/B _20513_/C _20513_/D VGND VGND VPWR VPWR _20514_/A sky130_fd_sc_hd__or4_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24281_ _32665_/Q _24280_/X _24305_/S VGND VGND VPWR VPWR _24282_/A sky130_fd_sc_hd__mux2_1
X_21493_ _21489_/X _21492_/X _21383_/X _21384_/X VGND VGND VPWR VPWR _21510_/B sky130_fd_sc_hd__o211a_1
X_33479_ _33544_/CLK _33479_/D VGND VGND VPWR VPWR _33479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26020_ _26020_/A VGND VGND VPWR VPWR _33426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20444_ _18297_/X _20442_/X _20443_/X _18303_/X VGND VGND VPWR VPWR _20444_/X sky130_fd_sc_hd__a22o_1
X_35218_ _35282_/CLK _35218_/D VGND VGND VPWR VPWR _35218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23232_ _32195_/Q _23231_/X _23235_/S VGND VGND VPWR VPWR _23233_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36198_ _36200_/CLK _36198_/D VGND VGND VPWR VPWR _36198_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_88_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35149_ _35277_/CLK _35149_/D VGND VGND VPWR VPWR _35149_/Q sky130_fd_sc_hd__dfxtp_1
X_23163_ _32165_/Q _23090_/X _23182_/S VGND VGND VPWR VPWR _23164_/A sky130_fd_sc_hd__mux2_1
X_20375_ _32519_/Q _32391_/Q _32071_/Q _36039_/Q _20282_/X _20070_/X VGND VGND VPWR
+ VPWR _20375_/X sky130_fd_sc_hd__mux4_1
XTAP_7106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22114_ _22467_/A VGND VGND VPWR VPWR _22114_/X sky130_fd_sc_hd__clkbuf_2
XTAP_7139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23094_ _32144_/Q _23093_/X _23115_/S VGND VGND VPWR VPWR _23095_/A sky130_fd_sc_hd__mux2_1
X_27971_ _27971_/A VGND VGND VPWR VPWR _34318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_288_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _36092_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26922_ input26/X VGND VGND VPWR VPWR _26922_/X sky130_fd_sc_hd__buf_4
X_29710_ _35112_/Q _29132_/X _29716_/S VGND VGND VPWR VPWR _29711_/A sky130_fd_sc_hd__mux2_1
X_22045_ _21795_/X _22041_/X _22044_/X _21800_/X VGND VGND VPWR VPWR _22045_/X sky130_fd_sc_hd__a22o_1
XTAP_6449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29641_ _29641_/A VGND VGND VPWR VPWR _35079_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26853_ input2/X VGND VGND VPWR VPWR _26853_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25804_ _25084_/X _33324_/Q _25822_/S VGND VGND VPWR VPWR _25805_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29572_ _29572_/A VGND VGND VPWR VPWR _35046_/D sky130_fd_sc_hd__clkbuf_1
X_26784_ _33788_/Q _24388_/X _26790_/S VGND VGND VPWR VPWR _26785_/A sky130_fd_sc_hd__mux2_1
X_23996_ _22910_/X _32536_/Q _24014_/S VGND VGND VPWR VPWR _23997_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28523_ _28523_/A VGND VGND VPWR VPWR _34580_/D sky130_fd_sc_hd__clkbuf_1
X_25735_ _33293_/Q _24440_/X _25735_/S VGND VGND VPWR VPWR _25736_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22947_ _22947_/A VGND VGND VPWR VPWR _32035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_460_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _35942_/CLK sky130_fd_sc_hd__clkbuf_16
X_28454_ _26940_/X _34548_/Q _28456_/S VGND VGND VPWR VPWR _28455_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25666_ _25735_/S VGND VGND VPWR VPWR _25685_/S sky130_fd_sc_hd__buf_4
XFILLER_95_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22878_ _31545_/A input83/X _23561_/B VGND VGND VPWR VPWR _22879_/A sky130_fd_sc_hd__or3b_1
X_27405_ _27405_/A VGND VGND VPWR VPWR _34051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24617_ _22929_/X _32798_/Q _24623_/S VGND VGND VPWR VPWR _24618_/A sky130_fd_sc_hd__mux2_1
X_28385_ _26838_/X _34515_/Q _28393_/S VGND VGND VPWR VPWR _28386_/A sky130_fd_sc_hd__mux2_1
X_21829_ _21754_/X _21827_/X _21828_/X _21759_/X VGND VGND VPWR VPWR _21829_/X sky130_fd_sc_hd__a22o_1
X_25597_ _33229_/Q _24440_/X _25597_/S VGND VGND VPWR VPWR _25598_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_212_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _35847_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_197_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27336_ _27336_/A VGND VGND VPWR VPWR _34018_/D sky130_fd_sc_hd__clkbuf_1
X_24548_ _23031_/X _32767_/Q _24548_/S VGND VGND VPWR VPWR _24549_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27267_ _26984_/X _33986_/Q _27281_/S VGND VGND VPWR VPWR _27268_/A sky130_fd_sc_hd__mux2_1
X_24479_ _22929_/X _32734_/Q _24485_/S VGND VGND VPWR VPWR _24480_/A sky130_fd_sc_hd__mux2_1
X_29006_ _29006_/A VGND VGND VPWR VPWR _34809_/D sky130_fd_sc_hd__clkbuf_1
X_17020_ _17846_/A VGND VGND VPWR VPWR _17020_/X sky130_fd_sc_hd__buf_6
XFILLER_8_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26218_ _26218_/A VGND VGND VPWR VPWR _33520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1083 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27198_ _27198_/A VGND VGND VPWR VPWR _33953_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_15_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_15_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_109_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26149_ _26149_/A VGND VGND VPWR VPWR _33487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_784 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18971_ _18965_/X _18970_/X _18722_/X VGND VGND VPWR VPWR _18993_/A sky130_fd_sc_hd__o21ba_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_279_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _36154_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29908_ _35206_/Q _29225_/X _29914_/S VGND VGND VPWR VPWR _29909_/A sky130_fd_sc_hd__mux2_1
X_17922_ _35778_/Q _35138_/Q _34498_/Q _33858_/Q _17846_/X _17847_/X VGND VGND VPWR
+ VPWR _17922_/X sky130_fd_sc_hd__mux4_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17853_ _17853_/A VGND VGND VPWR VPWR _17853_/X sky130_fd_sc_hd__buf_2
XFILLER_113_1106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29839_ _35173_/Q _29123_/X _29851_/S VGND VGND VPWR VPWR _29840_/A sky130_fd_sc_hd__mux2_1
XTAP_6994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16804_ _17157_/A VGND VGND VPWR VPWR _16804_/X sky130_fd_sc_hd__buf_4
XFILLER_226_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32850_ _32978_/CLK _32850_/D VGND VGND VPWR VPWR _32850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17784_ _17778_/X _17783_/X _17500_/X VGND VGND VPWR VPWR _17792_/C sky130_fd_sc_hd__o21ba_1
X_31801_ _36103_/Q input53/X _31805_/S VGND VGND VPWR VPWR _31802_/A sky130_fd_sc_hd__mux2_1
X_19523_ _35310_/Q _35246_/Q _35182_/Q _32302_/Q _19306_/X _19307_/X VGND VGND VPWR
+ VPWR _19523_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16735_ _33761_/Q _33697_/Q _33633_/Q _33569_/Q _16490_/X _16491_/X VGND VGND VPWR
+ VPWR _16735_/X sky130_fd_sc_hd__mux4_1
XFILLER_207_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32781_ _36173_/CLK _32781_/D VGND VGND VPWR VPWR _32781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_451_CLK clkbuf_6_9__f_CLK/X VGND VGND VPWR VPWR _35300_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_207_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34520_ _35292_/CLK _34520_/D VGND VGND VPWR VPWR _34520_/Q sky130_fd_sc_hd__dfxtp_1
X_19454_ _19454_/A VGND VGND VPWR VPWR _19454_/X sky130_fd_sc_hd__clkbuf_4
X_31732_ _36070_/Q input17/X _31742_/S VGND VGND VPWR VPWR _31733_/A sky130_fd_sc_hd__mux2_1
X_16666_ _33503_/Q _33439_/Q _33375_/Q _33311_/Q _16417_/X _16418_/X VGND VGND VPWR
+ VPWR _16666_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18405_ _34255_/Q _34191_/Q _34127_/Q _34063_/Q _18305_/X _18307_/X VGND VGND VPWR
+ VPWR _18405_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34451_ _35730_/CLK _34451_/D VGND VGND VPWR VPWR _34451_/Q sky130_fd_sc_hd__dfxtp_1
X_31663_ _31663_/A VGND VGND VPWR VPWR _36037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19385_ _19381_/X _19384_/X _19108_/X VGND VGND VPWR VPWR _19386_/D sky130_fd_sc_hd__o21ba_1
X_16597_ _34013_/Q _33949_/Q _33885_/Q _32157_/Q _16314_/X _16315_/X VGND VGND VPWR
+ VPWR _16597_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_203_CLK clkbuf_6_52__f_CLK/X VGND VGND VPWR VPWR _35715_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_188_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33402_ _33787_/CLK _33402_/D VGND VGND VPWR VPWR _33402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18336_ _32974_/Q _32910_/Q _32846_/Q _32782_/Q _18333_/X _18335_/X VGND VGND VPWR
+ VPWR _18336_/X sky130_fd_sc_hd__mux4_1
X_30614_ _35540_/Q _29070_/X _30620_/S VGND VGND VPWR VPWR _30615_/A sky130_fd_sc_hd__mux2_1
X_34382_ _34638_/CLK _34382_/D VGND VGND VPWR VPWR _34382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31594_ _31594_/A VGND VGND VPWR VPWR _36004_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36121_ _36121_/CLK _36121_/D VGND VGND VPWR VPWR _36121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18267_ _35341_/Q _35277_/Q _35213_/Q _32333_/Q _16088_/X _16090_/X VGND VGND VPWR
+ VPWR _18267_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30545_ _30545_/A VGND VGND VPWR VPWR _35507_/D sky130_fd_sc_hd__clkbuf_1
X_33333_ _33780_/CLK _33333_/D VGND VGND VPWR VPWR _33333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36052_ _36052_/CLK _36052_/D VGND VGND VPWR VPWR _36052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17218_ _35566_/Q _35502_/Q _35438_/Q _35374_/Q _16897_/X _16898_/X VGND VGND VPWR
+ VPWR _17218_/X sky130_fd_sc_hd__mux4_1
X_18198_ _18194_/X _18197_/X _17842_/A _17843_/A VGND VGND VPWR VPWR _18213_/B sky130_fd_sc_hd__o211a_1
X_30476_ _30476_/A VGND VGND VPWR VPWR _35474_/D sky130_fd_sc_hd__clkbuf_1
X_33264_ _36081_/CLK _33264_/D VGND VGND VPWR VPWR _33264_/Q sky130_fd_sc_hd__dfxtp_1
X_35003_ _35515_/CLK _35003_/D VGND VGND VPWR VPWR _35003_/Q sky130_fd_sc_hd__dfxtp_1
X_17149_ _17149_/A VGND VGND VPWR VPWR _17149_/X sky130_fd_sc_hd__clkbuf_4
X_32215_ _33255_/CLK _32215_/D VGND VGND VPWR VPWR _32215_/Q sky130_fd_sc_hd__dfxtp_1
X_33195_ _35307_/CLK _33195_/D VGND VGND VPWR VPWR _33195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_16__f_CLK clkbuf_5_8_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_96_CLK/A sky130_fd_sc_hd__clkbuf_16
X_20160_ _20160_/A VGND VGND VPWR VPWR _20160_/X sky130_fd_sc_hd__buf_4
X_32146_ _34006_/CLK _32146_/D VGND VGND VPWR VPWR _32146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32077_ _36045_/CLK _32077_/D VGND VGND VPWR VPWR _32077_/Q sky130_fd_sc_hd__dfxtp_1
X_20091_ _20087_/X _20090_/X _19814_/X VGND VGND VPWR VPWR _20092_/D sky130_fd_sc_hd__o21ba_1
X_35905_ _35906_/CLK _35905_/D VGND VGND VPWR VPWR _35905_/Q sky130_fd_sc_hd__dfxtp_1
X_31028_ _35736_/Q _29082_/X _31046_/S VGND VGND VPWR VPWR _31029_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35836_ _35965_/CLK _35836_/D VGND VGND VPWR VPWR _35836_/Q sky130_fd_sc_hd__dfxtp_1
X_23850_ _23850_/A VGND VGND VPWR VPWR _32467_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22801_ _20577_/X _22799_/X _22800_/X _20587_/X VGND VGND VPWR VPWR _22801_/X sky130_fd_sc_hd__a22o_1
XFILLER_26_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35767_ _35833_/CLK _35767_/D VGND VGND VPWR VPWR _35767_/Q sky130_fd_sc_hd__dfxtp_1
X_23781_ _23781_/A VGND VGND VPWR VPWR _32435_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32979_ _36052_/CLK _32979_/D VGND VGND VPWR VPWR _32979_/Q sky130_fd_sc_hd__dfxtp_1
X_20993_ _20949_/X _20991_/X _20992_/X _20955_/X VGND VGND VPWR VPWR _20993_/X sky130_fd_sc_hd__a22o_1
XFILLER_25_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_609 _18435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25520_ _33192_/Q _24326_/X _25526_/S VGND VGND VPWR VPWR _25521_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_442_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _36007_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_225_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22732_ _32777_/Q _32713_/Q _32649_/Q _36105_/Q _22578_/X _21473_/A VGND VGND VPWR
+ VPWR _22732_/X sky130_fd_sc_hd__mux4_1
X_34718_ _34781_/CLK _34718_/D VGND VGND VPWR VPWR _34718_/Q sky130_fd_sc_hd__dfxtp_1
X_35698_ _35826_/CLK _35698_/D VGND VGND VPWR VPWR _35698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_958 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25451_ _25451_/A VGND VGND VPWR VPWR _33161_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22663_ _22663_/A _22663_/B _22663_/C _22663_/D VGND VGND VPWR VPWR _22664_/A sky130_fd_sc_hd__or4_4
X_34649_ _36201_/CLK _34649_/D VGND VGND VPWR VPWR _34649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24402_ _32704_/Q _24400_/X _24429_/S VGND VGND VPWR VPWR _24403_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28170_ _26919_/X _34413_/Q _28186_/S VGND VGND VPWR VPWR _28171_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21614_ _21614_/A _21614_/B _21614_/C _21614_/D VGND VGND VPWR VPWR _21615_/A sky130_fd_sc_hd__or4_4
XFILLER_240_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25382_ _25382_/A VGND VGND VPWR VPWR _33128_/D sky130_fd_sc_hd__clkbuf_1
X_22594_ _22594_/A VGND VGND VPWR VPWR _22594_/X sky130_fd_sc_hd__buf_6
XFILLER_146_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27121_ _26968_/X _33917_/Q _27125_/S VGND VGND VPWR VPWR _27122_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24333_ _32682_/Q _24332_/X _24336_/S VGND VGND VPWR VPWR _24334_/A sky130_fd_sc_hd__mux2_1
X_21545_ _21545_/A VGND VGND VPWR VPWR _36198_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27052_ _26866_/X _33884_/Q _27062_/S VGND VGND VPWR VPWR _27053_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24264_ input61/X VGND VGND VPWR VPWR _24264_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21476_ _21401_/X _21474_/X _21475_/X _21406_/X VGND VGND VPWR VPWR _21476_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26003_ _25180_/X _33419_/Q _26007_/S VGND VGND VPWR VPWR _26004_/A sky130_fd_sc_hd__mux2_1
X_23215_ _32189_/Q _23199_/X _23235_/S VGND VGND VPWR VPWR _23216_/A sky130_fd_sc_hd__mux2_1
X_20427_ _20201_/X _20425_/X _20426_/X _20206_/X VGND VGND VPWR VPWR _20427_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24195_ _23003_/X _32630_/Q _24213_/S VGND VGND VPWR VPWR _24196_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23146_ _32161_/Q _23145_/X _23146_/S VGND VGND VPWR VPWR _23147_/A sky130_fd_sc_hd__mux2_1
X_20358_ _20155_/X _20356_/X _20357_/X _20158_/X VGND VGND VPWR VPWR _20358_/X sky130_fd_sc_hd__a22o_1
XTAP_6202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1008 _17862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27954_ _34311_/Q _24422_/X _27958_/S VGND VGND VPWR VPWR _27955_/A sky130_fd_sc_hd__mux2_1
XANTENNA_1019 _17858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20289_ _20000_/X _20287_/X _20288_/X _20003_/X VGND VGND VPWR VPWR _20289_/X sky130_fd_sc_hd__a22o_1
X_23077_ input1/X VGND VGND VPWR VPWR _23077_/X sky130_fd_sc_hd__buf_4
XTAP_6246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26905_ _26905_/A VGND VGND VPWR VPWR _33832_/D sky130_fd_sc_hd__clkbuf_1
X_22028_ _22532_/A VGND VGND VPWR VPWR _22028_/X sky130_fd_sc_hd__buf_4
XTAP_6279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27885_ _34278_/Q _24320_/X _27895_/S VGND VGND VPWR VPWR _27886_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29624_ _29624_/A VGND VGND VPWR VPWR _35071_/D sky130_fd_sc_hd__clkbuf_1
X_26836_ _26835_/X _33810_/Q _26851_/S VGND VGND VPWR VPWR _26837_/A sky130_fd_sc_hd__mux2_1
XTAP_4844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29555_ _29555_/A VGND VGND VPWR VPWR _35038_/D sky130_fd_sc_hd__clkbuf_1
X_26767_ _33780_/Q _24363_/X _26769_/S VGND VGND VPWR VPWR _26768_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23979_ _22886_/X _32528_/Q _23993_/S VGND VGND VPWR VPWR _23980_/A sky130_fd_sc_hd__mux2_1
XTAP_4899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_433_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _34281_/CLK sky130_fd_sc_hd__clkbuf_16
X_16520_ _16873_/A VGND VGND VPWR VPWR _16520_/X sky130_fd_sc_hd__buf_4
XFILLER_244_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28506_ _27017_/X _34573_/Q _28506_/S VGND VGND VPWR VPWR _28507_/A sky130_fd_sc_hd__mux2_1
X_25718_ _25718_/A VGND VGND VPWR VPWR _33284_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_941 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26698_ _33747_/Q _24261_/X _26706_/S VGND VGND VPWR VPWR _26699_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29486_ _23297_/X _35006_/Q _29488_/S VGND VGND VPWR VPWR _29487_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16451_ _17157_/A VGND VGND VPWR VPWR _16451_/X sky130_fd_sc_hd__buf_4
XFILLER_232_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28437_ _28506_/S VGND VGND VPWR VPWR _28456_/S sky130_fd_sc_hd__clkbuf_8
X_25649_ _25649_/A VGND VGND VPWR VPWR _33251_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19170_ _35300_/Q _35236_/Q _35172_/Q _32292_/Q _18953_/X _18954_/X VGND VGND VPWR
+ VPWR _19170_/X sky130_fd_sc_hd__mux4_1
X_28368_ _28368_/A VGND VGND VPWR VPWR _34507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16382_ _33751_/Q _33687_/Q _33623_/Q _33559_/Q _16137_/X _16138_/X VGND VGND VPWR
+ VPWR _16382_/X sky130_fd_sc_hd__mux4_1
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18121_ _17860_/X _18119_/X _18120_/X _17865_/X VGND VGND VPWR VPWR _18121_/X sky130_fd_sc_hd__a22o_1
XFILLER_223_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27319_ _27319_/A VGND VGND VPWR VPWR _34010_/D sky130_fd_sc_hd__clkbuf_1
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28299_ _28299_/A VGND VGND VPWR VPWR _34474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30330_ _30735_/A _31410_/B VGND VGND VPWR VPWR _30463_/S sky130_fd_sc_hd__nand2_8
X_18052_ _35590_/Q _35526_/Q _35462_/Q _35398_/Q _17956_/X _17957_/X VGND VGND VPWR
+ VPWR _18052_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17003_ _16999_/X _17000_/X _17001_/X _17002_/X VGND VGND VPWR VPWR _17003_/X sky130_fd_sc_hd__a22o_1
X_30261_ _35373_/Q _29148_/X _30277_/S VGND VGND VPWR VPWR _30262_/A sky130_fd_sc_hd__mux2_1
XANTENNA_5 _32114_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32000_ _33946_/CLK _32000_/D VGND VGND VPWR VPWR _32000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30192_ _35341_/Q _29246_/X _30192_/S VGND VGND VPWR VPWR _30193_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18954_ _19307_/A VGND VGND VPWR VPWR _18954_/X sky130_fd_sc_hd__buf_4
XFILLER_98_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17905_ _34306_/Q _34242_/Q _34178_/Q _34114_/Q _17795_/X _17796_/X VGND VGND VPWR
+ VPWR _17905_/X sky130_fd_sc_hd__mux4_1
X_33951_ _34016_/CLK _33951_/D VGND VGND VPWR VPWR _33951_/Q sky130_fd_sc_hd__dfxtp_1
X_18885_ _35292_/Q _35228_/Q _35164_/Q _32284_/Q _18600_/X _18601_/X VGND VGND VPWR
+ VPWR _18885_/X sky130_fd_sc_hd__mux4_1
XTAP_6780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32902_ _36039_/CLK _32902_/D VGND VGND VPWR VPWR _32902_/Q sky130_fd_sc_hd__dfxtp_1
X_17836_ _32768_/Q _32704_/Q _32640_/Q _36096_/Q _17625_/X _17762_/X VGND VGND VPWR
+ VPWR _17836_/X sky130_fd_sc_hd__mux4_1
X_33882_ _33946_/CLK _33882_/D VGND VGND VPWR VPWR _33882_/Q sky130_fd_sc_hd__dfxtp_1
X_35621_ _35814_/CLK _35621_/D VGND VGND VPWR VPWR _35621_/Q sky130_fd_sc_hd__dfxtp_1
X_32833_ _36033_/CLK _32833_/D VGND VGND VPWR VPWR _32833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17767_ _17767_/A VGND VGND VPWR VPWR _17767_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_130_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_424_CLK clkbuf_6_36__f_CLK/X VGND VGND VPWR VPWR _34739_/CLK sky130_fd_sc_hd__clkbuf_16
X_19506_ _19502_/X _19503_/X _19504_/X _19505_/X VGND VGND VPWR VPWR _19506_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16718_ _35744_/Q _35104_/Q _34464_/Q _33824_/Q _16434_/X _16435_/X VGND VGND VPWR
+ VPWR _16718_/X sky130_fd_sc_hd__mux4_1
X_35552_ _35552_/CLK _35552_/D VGND VGND VPWR VPWR _35552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32764_ _36092_/CLK _32764_/D VGND VGND VPWR VPWR _32764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17698_ _17416_/X _17694_/X _17697_/X _17420_/X VGND VGND VPWR VPWR _17698_/X sky130_fd_sc_hd__a22o_1
XFILLER_63_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34503_ _35784_/CLK _34503_/D VGND VGND VPWR VPWR _34503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19437_ _20143_/A VGND VGND VPWR VPWR _19437_/X sky130_fd_sc_hd__clkbuf_4
X_31715_ _36062_/Q input8/X _31721_/S VGND VGND VPWR VPWR _31716_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16649_ _17865_/A VGND VGND VPWR VPWR _16649_/X sky130_fd_sc_hd__clkbuf_4
X_35483_ _35869_/CLK _35483_/D VGND VGND VPWR VPWR _35483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32695_ _36088_/CLK _32695_/D VGND VGND VPWR VPWR _32695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34434_ _34947_/CLK _34434_/D VGND VGND VPWR VPWR _34434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31646_ _31646_/A VGND VGND VPWR VPWR _36029_/D sky130_fd_sc_hd__clkbuf_1
X_19368_ _19363_/X _19365_/X _19366_/X _19367_/X VGND VGND VPWR VPWR _19368_/X sky130_fd_sc_hd__a22o_1
X_18319_ _32718_/Q _32654_/Q _32590_/Q _36046_/Q _20162_/A _20013_/A VGND VGND VPWR
+ VPWR _18319_/X sky130_fd_sc_hd__mux4_1
X_34365_ _35581_/CLK _34365_/D VGND VGND VPWR VPWR _34365_/Q sky130_fd_sc_hd__dfxtp_1
X_19299_ _20160_/A VGND VGND VPWR VPWR _19299_/X sky130_fd_sc_hd__clkbuf_4
X_31577_ _31577_/A VGND VGND VPWR VPWR _35996_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36104_ _36169_/CLK _36104_/D VGND VGND VPWR VPWR _36104_/Q sky130_fd_sc_hd__dfxtp_1
X_33316_ _33702_/CLK _33316_/D VGND VGND VPWR VPWR _33316_/Q sky130_fd_sc_hd__dfxtp_1
X_21330_ _35040_/Q _34976_/Q _34912_/Q _34848_/Q _21050_/X _21051_/X VGND VGND VPWR
+ VPWR _21330_/X sky130_fd_sc_hd__mux4_1
X_30528_ _30528_/A VGND VGND VPWR VPWR _35499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34296_ _34296_/CLK _34296_/D VGND VGND VPWR VPWR _34296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36035_ _36037_/CLK _36035_/D VGND VGND VPWR VPWR _36035_/Q sky130_fd_sc_hd__dfxtp_1
X_30459_ _23339_/X _35467_/Q _30463_/S VGND VGND VPWR VPWR _30460_/A sky130_fd_sc_hd__mux2_1
X_21261_ _21261_/A _21261_/B _21261_/C _21261_/D VGND VGND VPWR VPWR _21262_/A sky130_fd_sc_hd__or4_2
X_33247_ _34016_/CLK _33247_/D VGND VGND VPWR VPWR _33247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23000_ input33/X VGND VGND VPWR VPWR _23000_/X sky130_fd_sc_hd__buf_2
XFILLER_237_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20212_ _20208_/X _20209_/X _20210_/X _20211_/X VGND VGND VPWR VPWR _20212_/X sky130_fd_sc_hd__a22o_1
XFILLER_150_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21192_ _21192_/A VGND VGND VPWR VPWR _36188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33178_ _35864_/CLK _33178_/D VGND VGND VPWR VPWR _33178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20143_ _20143_/A VGND VGND VPWR VPWR _20143_/X sky130_fd_sc_hd__buf_4
XFILLER_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32129_ _35562_/CLK _32129_/D VGND VGND VPWR VPWR _32129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20074_ _20069_/X _20071_/X _20072_/X _20073_/X VGND VGND VPWR VPWR _20074_/X sky130_fd_sc_hd__a22o_1
X_24951_ _24951_/A VGND VGND VPWR VPWR _32955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23902_ _22972_/X _32492_/Q _23920_/S VGND VGND VPWR VPWR _23903_/A sky130_fd_sc_hd__mux2_1
X_27670_ _34176_/Q _24400_/X _27688_/S VGND VGND VPWR VPWR _27671_/A sky130_fd_sc_hd__mux2_1
XTAP_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24882_ _24882_/A VGND VGND VPWR VPWR _32922_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26621_ _25094_/X _33711_/Q _26633_/S VGND VGND VPWR VPWR _26622_/A sky130_fd_sc_hd__mux2_1
X_23833_ _23833_/A VGND VGND VPWR VPWR _32460_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35819_ _35819_/CLK _35819_/D VGND VGND VPWR VPWR _35819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_406 _36211_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_415_CLK clkbuf_6_35__f_CLK/X VGND VGND VPWR VPWR _35308_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_417 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26552_ _24989_/X _33678_/Q _26570_/S VGND VGND VPWR VPWR _26553_/A sky130_fd_sc_hd__mux2_1
X_29340_ _29340_/A VGND VGND VPWR VPWR _34936_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23764_ _23764_/A VGND VGND VPWR VPWR _32427_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_428 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20976_ _34518_/Q _32406_/Q _34390_/Q _34326_/Q _20766_/X _20767_/X VGND VGND VPWR
+ VPWR _20976_/X sky130_fd_sc_hd__mux4_1
XANTENNA_439 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25503_ _33184_/Q _24301_/X _25505_/S VGND VGND VPWR VPWR _25504_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22715_ _22711_/X _22714_/X _22453_/X VGND VGND VPWR VPWR _22723_/C sky130_fd_sc_hd__o21ba_1
XFILLER_214_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29271_ _29382_/S VGND VGND VPWR VPWR _29290_/S sky130_fd_sc_hd__buf_4
XFILLER_92_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26483_ _25091_/X _33646_/Q _26497_/S VGND VGND VPWR VPWR _26484_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23695_ _23695_/A VGND VGND VPWR VPWR _32396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28222_ _26996_/X _34438_/Q _28228_/S VGND VGND VPWR VPWR _28223_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25434_ _25150_/X _33153_/Q _25450_/S VGND VGND VPWR VPWR _25435_/A sky130_fd_sc_hd__mux2_1
X_22646_ _33030_/Q _32966_/Q _32902_/Q _32838_/Q _20580_/X _20583_/X VGND VGND VPWR
+ VPWR _22646_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28153_ _26894_/X _34405_/Q _28165_/S VGND VGND VPWR VPWR _28154_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25365_ _25365_/A VGND VGND VPWR VPWR _33120_/D sky130_fd_sc_hd__clkbuf_1
X_22577_ _22573_/X _22576_/X _22434_/X VGND VGND VPWR VPWR _22603_/A sky130_fd_sc_hd__o21ba_1
XFILLER_139_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27104_ _26943_/X _33909_/Q _27104_/S VGND VGND VPWR VPWR _27105_/A sky130_fd_sc_hd__mux2_1
X_24316_ _24316_/A VGND VGND VPWR VPWR _32676_/D sky130_fd_sc_hd__clkbuf_1
X_28084_ _28084_/A VGND VGND VPWR VPWR _34372_/D sky130_fd_sc_hd__clkbuf_1
X_21528_ _35814_/Q _32190_/Q _35686_/Q _35622_/Q _21207_/X _21208_/X VGND VGND VPWR
+ VPWR _21528_/X sky130_fd_sc_hd__mux4_1
X_25296_ _25146_/X _33088_/Q _25314_/S VGND VGND VPWR VPWR _25297_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27035_ _26841_/X _33876_/Q _27041_/S VGND VGND VPWR VPWR _27036_/A sky130_fd_sc_hd__mux2_1
X_24247_ _32654_/Q _24244_/X _24274_/S VGND VGND VPWR VPWR _24248_/A sky130_fd_sc_hd__mux2_1
X_21459_ _32996_/Q _32932_/Q _32868_/Q _32804_/Q _21236_/X _21237_/X VGND VGND VPWR
+ VPWR _21459_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24178_ _22979_/X _32622_/Q _24192_/S VGND VGND VPWR VPWR _24179_/A sky130_fd_sc_hd__mux2_1
XTAP_6010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23129_ _23129_/A VGND VGND VPWR VPWR _32155_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_968 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28986_ _34800_/Q _24351_/X _28996_/S VGND VGND VPWR VPWR _28987_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_6_62__f_CLK clkbuf_5_31_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_62__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XTAP_6043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput97 _31966_/Q VGND VGND VPWR VPWR D1[16] sky130_fd_sc_hd__buf_2
XFILLER_49_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27937_ _34303_/Q _24397_/X _27937_/S VGND VGND VPWR VPWR _27938_/A sky130_fd_sc_hd__mux2_1
XTAP_6076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18670_ _33174_/Q _32534_/Q _35926_/Q _35862_/Q _18668_/X _18669_/X VGND VGND VPWR
+ VPWR _18670_/X sky130_fd_sc_hd__mux4_1
XTAP_5375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27868_ _34270_/Q _24295_/X _27874_/S VGND VGND VPWR VPWR _27869_/A sky130_fd_sc_hd__mux2_1
XTAP_5386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ _33530_/Q _33466_/Q _33402_/Q _33338_/Q _17476_/X _17477_/X VGND VGND VPWR
+ VPWR _17621_/X sky130_fd_sc_hd__mux4_1
X_29607_ _35063_/Q _29179_/X _29623_/S VGND VGND VPWR VPWR _29608_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26819_ _33805_/Q _24440_/X _26819_/S VGND VGND VPWR VPWR _26820_/A sky130_fd_sc_hd__mux2_1
XTAP_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27799_ _27799_/A VGND VGND VPWR VPWR _34237_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_930 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_406_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _35947_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29538_ _29538_/A VGND VGND VPWR VPWR _35030_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ _34296_/Q _34232_/Q _34168_/Q _34104_/Q _17442_/X _17443_/X VGND VGND VPWR
+ VPWR _17552_/X sky130_fd_sc_hd__mux4_1
XTAP_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_940 _29382_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_951 _29652_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16503_ _33242_/Q _36122_/Q _33114_/Q _33050_/Q _16352_/X _16353_/X VGND VGND VPWR
+ VPWR _16503_/X sky130_fd_sc_hd__mux4_1
XANTENNA_962 _30057_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17483_ _32758_/Q _32694_/Q _32630_/Q _36086_/Q _17272_/X _17409_/X VGND VGND VPWR
+ VPWR _17483_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29469_ _29517_/S VGND VGND VPWR VPWR _29488_/S sky130_fd_sc_hd__buf_4
XFILLER_60_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_944 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_973 _31813_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_984 _17795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31500_ _23277_/X _35960_/Q _31514_/S VGND VGND VPWR VPWR _31501_/A sky130_fd_sc_hd__mux2_1
XANTENNA_995 _17956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19222_ _19002_/X _19220_/X _19221_/X _19008_/X VGND VGND VPWR VPWR _19222_/X sky130_fd_sc_hd__a22o_1
X_16434_ _17994_/A VGND VGND VPWR VPWR _16434_/X sky130_fd_sc_hd__buf_6
XFILLER_34_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32480_ _36001_/CLK _32480_/D VGND VGND VPWR VPWR _32480_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16365_ _35734_/Q _35094_/Q _34454_/Q _33814_/Q _16049_/X _16051_/X VGND VGND VPWR
+ VPWR _16365_/X sky130_fd_sc_hd__mux4_1
X_31431_ _31431_/A VGND VGND VPWR VPWR _35927_/D sky130_fd_sc_hd__clkbuf_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19153_ _19149_/X _19150_/X _19151_/X _19152_/X VGND VGND VPWR VPWR _19153_/X sky130_fd_sc_hd__a22o_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18104_ _17149_/A _18102_/X _18103_/X _17152_/A VGND VGND VPWR VPWR _18104_/X sky130_fd_sc_hd__a22o_1
XFILLER_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31362_ _31362_/A VGND VGND VPWR VPWR _35894_/D sky130_fd_sc_hd__clkbuf_1
X_34150_ _34277_/CLK _34150_/D VGND VGND VPWR VPWR _34150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16296_ _17865_/A VGND VGND VPWR VPWR _16296_/X sky130_fd_sc_hd__buf_4
XFILLER_117_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19084_ _20143_/A VGND VGND VPWR VPWR _19084_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_195_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30313_ _35398_/Q _29225_/X _30319_/S VGND VGND VPWR VPWR _30314_/A sky130_fd_sc_hd__mux2_1
X_33101_ _34316_/CLK _33101_/D VGND VGND VPWR VPWR _33101_/Q sky130_fd_sc_hd__dfxtp_1
X_18035_ _33798_/Q _33734_/Q _33670_/Q _33606_/Q _17902_/X _17903_/X VGND VGND VPWR
+ VPWR _18035_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31293_ _35862_/Q input63/X _31295_/S VGND VGND VPWR VPWR _31294_/A sky130_fd_sc_hd__mux2_1
X_34081_ _36124_/CLK _34081_/D VGND VGND VPWR VPWR _34081_/Q sky130_fd_sc_hd__dfxtp_1
X_33032_ _35909_/CLK _33032_/D VGND VGND VPWR VPWR _33032_/Q sky130_fd_sc_hd__dfxtp_1
X_30244_ _35365_/Q _29123_/X _30256_/S VGND VGND VPWR VPWR _30245_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30175_ _30175_/A VGND VGND VPWR VPWR _35332_/D sky130_fd_sc_hd__clkbuf_1
X_19986_ _19848_/X _19984_/X _19985_/X _19853_/X VGND VGND VPWR VPWR _19986_/X sky130_fd_sc_hd__a22o_1
XFILLER_140_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18937_ _20130_/A VGND VGND VPWR VPWR _18937_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_101_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34983_ _35943_/CLK _34983_/D VGND VGND VPWR VPWR _34983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1350 _21757_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1361 _23133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1372 _25314_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33934_ _34262_/CLK _33934_/D VGND VGND VPWR VPWR _33934_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1383 _30598_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18868_ _33244_/Q _36124_/Q _33116_/Q _33052_/Q _18652_/X _18653_/X VGND VGND VPWR
+ VPWR _18868_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1394 input87/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17819_ _17502_/X _17817_/X _17818_/X _17505_/X VGND VGND VPWR VPWR _17819_/X sky130_fd_sc_hd__a22o_1
XFILLER_132_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33865_ _35845_/CLK _33865_/D VGND VGND VPWR VPWR _33865_/Q sky130_fd_sc_hd__dfxtp_1
X_18799_ _20165_/A VGND VGND VPWR VPWR _18799_/X sky130_fd_sc_hd__buf_4
XFILLER_208_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35604_ _35669_/CLK _35604_/D VGND VGND VPWR VPWR _35604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20830_ _22595_/A VGND VGND VPWR VPWR _20830_/X sky130_fd_sc_hd__buf_4
X_32816_ _33009_/CLK _32816_/D VGND VGND VPWR VPWR _32816_/Q sky130_fd_sc_hd__dfxtp_1
X_33796_ _34309_/CLK _33796_/D VGND VGND VPWR VPWR _33796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35535_ _35597_/CLK _35535_/D VGND VGND VPWR VPWR _35535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20761_ _20656_/X _20759_/X _20760_/X _20668_/X VGND VGND VPWR VPWR _20761_/X sky130_fd_sc_hd__a22o_1
X_32747_ _35187_/CLK _32747_/D VGND VGND VPWR VPWR _32747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22500_ _22500_/A VGND VGND VPWR VPWR _36225_/D sky130_fd_sc_hd__clkbuf_1
X_35466_ _35978_/CLK _35466_/D VGND VGND VPWR VPWR _35466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23480_ _22957_/X _32295_/Q _23488_/S VGND VGND VPWR VPWR _23481_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20692_ _22462_/A VGND VGND VPWR VPWR _20692_/X sky130_fd_sc_hd__buf_4
XFILLER_126_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32678_ _36135_/CLK _32678_/D VGND VGND VPWR VPWR _32678_/Q sky130_fd_sc_hd__dfxtp_1
X_22431_ _33536_/Q _33472_/Q _33408_/Q _33344_/Q _22429_/X _22430_/X VGND VGND VPWR
+ VPWR _22431_/X sky130_fd_sc_hd__mux4_1
X_34417_ _35052_/CLK _34417_/D VGND VGND VPWR VPWR _34417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31629_ _31629_/A VGND VGND VPWR VPWR _36021_/D sky130_fd_sc_hd__clkbuf_1
X_35397_ _36168_/CLK _35397_/D VGND VGND VPWR VPWR _35397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25150_ input47/X VGND VGND VPWR VPWR _25150_/X sky130_fd_sc_hd__buf_2
XFILLER_176_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22362_ _22362_/A VGND VGND VPWR VPWR _22362_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_136_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34348_ _35307_/CLK _34348_/D VGND VGND VPWR VPWR _34348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24101_ _24101_/A VGND VGND VPWR VPWR _32586_/D sky130_fd_sc_hd__clkbuf_1
X_21313_ _32992_/Q _32928_/Q _32864_/Q _32800_/Q _21236_/X _21237_/X VGND VGND VPWR
+ VPWR _21313_/X sky130_fd_sc_hd__mux4_1
X_25081_ input22/X VGND VGND VPWR VPWR _25081_/X sky130_fd_sc_hd__buf_2
X_22293_ _22008_/X _22291_/X _22292_/X _22014_/X VGND VGND VPWR VPWR _22293_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34279_ _34279_/CLK _34279_/D VGND VGND VPWR VPWR _34279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24032_ _24032_/A VGND VGND VPWR VPWR _32553_/D sky130_fd_sc_hd__clkbuf_1
X_36018_ _36018_/CLK _36018_/D VGND VGND VPWR VPWR _36018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21244_ _22458_/A VGND VGND VPWR VPWR _21244_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_85_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28840_ _26912_/X _34731_/Q _28840_/S VGND VGND VPWR VPWR _28841_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21175_ _35804_/Q _32179_/Q _35676_/Q _35612_/Q _20854_/X _20855_/X VGND VGND VPWR
+ VPWR _21175_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20126_ _33792_/Q _33728_/Q _33664_/Q _33600_/Q _19849_/X _19850_/X VGND VGND VPWR
+ VPWR _20126_/X sky130_fd_sc_hd__mux4_1
X_28771_ _28771_/A VGND VGND VPWR VPWR _34698_/D sky130_fd_sc_hd__clkbuf_1
X_25983_ _25150_/X _33409_/Q _25999_/S VGND VGND VPWR VPWR _25984_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20057_ _33534_/Q _33470_/Q _33406_/Q _33342_/Q _19776_/X _19777_/X VGND VGND VPWR
+ VPWR _20057_/X sky130_fd_sc_hd__mux4_1
X_27722_ _27722_/A VGND VGND VPWR VPWR _34200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24934_ _24934_/A VGND VGND VPWR VPWR _32947_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24865_ _24865_/A VGND VGND VPWR VPWR _32914_/D sky130_fd_sc_hd__clkbuf_1
X_27653_ _34168_/Q _24376_/X _27667_/S VGND VGND VPWR VPWR _27654_/A sky130_fd_sc_hd__mux2_1
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23816_ _23047_/X _32452_/Q _23826_/S VGND VGND VPWR VPWR _23817_/A sky130_fd_sc_hd__mux2_1
XFILLER_233_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_203 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26604_ _25069_/X _33703_/Q _26612_/S VGND VGND VPWR VPWR _26605_/A sky130_fd_sc_hd__mux2_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27584_ _27584_/A VGND VGND VPWR VPWR _34135_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_214 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_225 _32136_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24796_ _22991_/X _32882_/Q _24802_/S VGND VGND VPWR VPWR _24797_/A sky130_fd_sc_hd__mux2_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_236 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26535_ _25168_/X _33671_/Q _26539_/S VGND VGND VPWR VPWR _26536_/A sky130_fd_sc_hd__mux2_1
XANTENNA_247 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29323_ _29323_/A VGND VGND VPWR VPWR _34928_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23747_ _22945_/X _32419_/Q _23763_/S VGND VGND VPWR VPWR _23748_/A sky130_fd_sc_hd__mux2_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20959_ _32470_/Q _32342_/Q _32022_/Q _35990_/Q _20817_/X _20958_/X VGND VGND VPWR
+ VPWR _20959_/X sky130_fd_sc_hd__mux4_1
XANTENNA_269 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29254_ _29254_/A VGND VGND VPWR VPWR _34895_/D sky130_fd_sc_hd__clkbuf_1
X_26466_ _25066_/X _33638_/Q _26476_/S VGND VGND VPWR VPWR _26467_/A sky130_fd_sc_hd__mux2_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23678_ _32388_/Q _23316_/X _23688_/S VGND VGND VPWR VPWR _23679_/A sky130_fd_sc_hd__mux2_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28205_ _26971_/X _34430_/Q _28207_/S VGND VGND VPWR VPWR _28206_/A sky130_fd_sc_hd__mux2_1
X_25417_ _25125_/X _33145_/Q _25429_/S VGND VGND VPWR VPWR _25418_/A sky130_fd_sc_hd__mux2_1
X_22629_ _34565_/Q _32453_/Q _34437_/Q _34373_/Q _22531_/X _22532_/X VGND VGND VPWR
+ VPWR _22629_/X sky130_fd_sc_hd__mux4_1
X_29185_ input38/X VGND VGND VPWR VPWR _29185_/X sky130_fd_sc_hd__clkbuf_4
X_26397_ _26397_/A VGND VGND VPWR VPWR _33605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16150_ _33232_/Q _36112_/Q _33104_/Q _33040_/Q _16020_/X _16021_/X VGND VGND VPWR
+ VPWR _16150_/X sky130_fd_sc_hd__mux4_1
X_28136_ _26869_/X _34397_/Q _28144_/S VGND VGND VPWR VPWR _28137_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25348_ _25022_/X _33112_/Q _25366_/S VGND VGND VPWR VPWR _25349_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16081_ _17007_/A VGND VGND VPWR VPWR _16081_/X sky130_fd_sc_hd__buf_4
X_28067_ _28067_/A VGND VGND VPWR VPWR _34364_/D sky130_fd_sc_hd__clkbuf_1
X_25279_ _25122_/X _33080_/Q _25293_/S VGND VGND VPWR VPWR _25280_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27018_ _27017_/X _33869_/Q _27018_/S VGND VGND VPWR VPWR _27019_/A sky130_fd_sc_hd__mux2_1
X_19840_ _35319_/Q _35255_/Q _35191_/Q _32311_/Q _19659_/X _19660_/X VGND VGND VPWR
+ VPWR _19840_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19771_ _19771_/A _19771_/B _19771_/C _19771_/D VGND VGND VPWR VPWR _19772_/A sky130_fd_sc_hd__or4_2
X_28969_ _34792_/Q _24326_/X _28975_/S VGND VGND VPWR VPWR _28970_/A sky130_fd_sc_hd__mux2_1
X_16983_ _16849_/X _16981_/X _16982_/X _16852_/X VGND VGND VPWR VPWR _16983_/X sky130_fd_sc_hd__a22o_1
XFILLER_27_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18722_ _20134_/A VGND VGND VPWR VPWR _18722_/X sky130_fd_sc_hd__buf_2
XFILLER_114_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31980_ _34970_/CLK _31980_/D VGND VGND VPWR VPWR _31980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18653_ _20203_/A VGND VGND VPWR VPWR _18653_/X sky130_fd_sc_hd__clkbuf_4
X_30931_ _30931_/A VGND VGND VPWR VPWR _35690_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17604_ _17957_/A VGND VGND VPWR VPWR _17604_/X sky130_fd_sc_hd__buf_4
XTAP_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33650_ _34227_/CLK _33650_/D VGND VGND VPWR VPWR _33650_/Q sky130_fd_sc_hd__dfxtp_1
X_30862_ _23336_/X _35658_/Q _30868_/S VGND VGND VPWR VPWR _30863_/A sky130_fd_sc_hd__mux2_1
X_18584_ _20130_/A VGND VGND VPWR VPWR _18584_/X sky130_fd_sc_hd__buf_4
XTAP_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32601_ _36059_/CLK _32601_/D VGND VGND VPWR VPWR _32601_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17535_ _35575_/Q _35511_/Q _35447_/Q _35383_/Q _17250_/X _17251_/X VGND VGND VPWR
+ VPWR _17535_/X sky130_fd_sc_hd__mux4_1
X_33581_ _34283_/CLK _33581_/D VGND VGND VPWR VPWR _33581_/Q sky130_fd_sc_hd__dfxtp_1
X_30793_ _23228_/X _35625_/Q _30797_/S VGND VGND VPWR VPWR _30794_/A sky130_fd_sc_hd__mux2_1
XANTENNA_770 _22538_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_781 _22604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35320_ _35320_/CLK _35320_/D VGND VGND VPWR VPWR _35320_/Q sky130_fd_sc_hd__dfxtp_1
X_32532_ _36115_/CLK _32532_/D VGND VGND VPWR VPWR _32532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_792 _22694_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17466_ _17149_/X _17464_/X _17465_/X _17152_/X VGND VGND VPWR VPWR _17466_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_774 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19205_ _19096_/X _19203_/X _19204_/X _19099_/X VGND VGND VPWR VPWR _19205_/X sky130_fd_sc_hd__a22o_1
X_16417_ _17795_/A VGND VGND VPWR VPWR _16417_/X sky130_fd_sc_hd__buf_4
X_35251_ _36074_/CLK _35251_/D VGND VGND VPWR VPWR _35251_/Q sky130_fd_sc_hd__dfxtp_1
X_32463_ _36041_/CLK _32463_/D VGND VGND VPWR VPWR _32463_/Q sky130_fd_sc_hd__dfxtp_1
X_17397_ _17154_/X _17395_/X _17396_/X _17159_/X VGND VGND VPWR VPWR _17397_/X sky130_fd_sc_hd__a22o_1
XFILLER_207_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34202_ _34202_/CLK _34202_/D VGND VGND VPWR VPWR _34202_/Q sky130_fd_sc_hd__dfxtp_1
X_31414_ _23090_/X _35919_/Q _31430_/S VGND VGND VPWR VPWR _31415_/A sky130_fd_sc_hd__mux2_1
X_19136_ _34531_/Q _32419_/Q _34403_/Q _34339_/Q _18819_/X _18820_/X VGND VGND VPWR
+ VPWR _19136_/X sky130_fd_sc_hd__mux4_1
X_16348_ _16344_/X _16347_/X _16011_/X VGND VGND VPWR VPWR _16380_/A sky130_fd_sc_hd__o21ba_2
XFILLER_173_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35182_ _35500_/CLK _35182_/D VGND VGND VPWR VPWR _35182_/Q sky130_fd_sc_hd__dfxtp_1
X_32394_ _36109_/CLK _32394_/D VGND VGND VPWR VPWR _32394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34133_ _34197_/CLK _34133_/D VGND VGND VPWR VPWR _34133_/Q sky130_fd_sc_hd__dfxtp_1
X_16279_ _32724_/Q _32660_/Q _32596_/Q _36052_/Q _16213_/X _17713_/A VGND VGND VPWR
+ VPWR _16279_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19067_ _33762_/Q _33698_/Q _33634_/Q _33570_/Q _18790_/X _18791_/X VGND VGND VPWR
+ VPWR _19067_/X sky130_fd_sc_hd__mux4_1
X_31345_ _31345_/A VGND VGND VPWR VPWR _35886_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18018_ _18014_/X _18017_/X _17842_/X _17843_/X VGND VGND VPWR VPWR _18033_/B sky130_fd_sc_hd__o211a_1
XFILLER_160_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34064_ _35021_/CLK _34064_/D VGND VGND VPWR VPWR _34064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31276_ _31408_/S VGND VGND VPWR VPWR _31295_/S sky130_fd_sc_hd__buf_4
XFILLER_218_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33015_ _36087_/CLK _33015_/D VGND VGND VPWR VPWR _33015_/Q sky130_fd_sc_hd__dfxtp_1
X_30227_ _35357_/Q _29098_/X _30235_/S VGND VGND VPWR VPWR _30228_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30158_ _30158_/A VGND VGND VPWR VPWR _35324_/D sky130_fd_sc_hd__clkbuf_1
X_19969_ _35771_/Q _35131_/Q _34491_/Q _33851_/Q _19793_/X _19794_/X VGND VGND VPWR
+ VPWR _19969_/X sky130_fd_sc_hd__mux4_1
XFILLER_87_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1063 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34966_ _35028_/CLK _34966_/D VGND VGND VPWR VPWR _34966_/Q sky130_fd_sc_hd__dfxtp_1
X_22980_ _22979_/X _32046_/Q _23001_/S VGND VGND VPWR VPWR _22981_/A sky130_fd_sc_hd__mux2_1
X_30089_ _30089_/A VGND VGND VPWR VPWR _35291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1180 _21333_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1191 _22883_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33917_ _34046_/CLK _33917_/D VGND VGND VPWR VPWR _33917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21931_ _33778_/Q _33714_/Q _33650_/Q _33586_/Q _21796_/X _21797_/X VGND VGND VPWR
+ VPWR _21931_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34897_ _36204_/CLK _34897_/D VGND VGND VPWR VPWR _34897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_880 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24650_ _24650_/A VGND VGND VPWR VPWR _32813_/D sky130_fd_sc_hd__clkbuf_1
X_33848_ _35768_/CLK _33848_/D VGND VGND VPWR VPWR _33848_/Q sky130_fd_sc_hd__dfxtp_1
X_21862_ _21858_/X _21861_/X _21761_/X VGND VGND VPWR VPWR _21863_/D sky130_fd_sc_hd__o21ba_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23601_ _23601_/A VGND VGND VPWR VPWR _32351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20813_ _22578_/A VGND VGND VPWR VPWR _20813_/X sky130_fd_sc_hd__buf_6
X_24581_ _24581_/A VGND VGND VPWR VPWR _31815_/B sky130_fd_sc_hd__buf_12
XFILLER_82_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21793_ _21793_/A _21793_/B _21793_/C _21793_/D VGND VGND VPWR VPWR _21794_/A sky130_fd_sc_hd__or4_1
XFILLER_35_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33779_ _33779_/CLK _33779_/D VGND VGND VPWR VPWR _33779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26320_ _25050_/X _33569_/Q _26320_/S VGND VGND VPWR VPWR _26321_/A sky130_fd_sc_hd__mux2_1
XFILLER_247_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23532_ _23559_/S VGND VGND VPWR VPWR _23551_/S sky130_fd_sc_hd__buf_6
X_35518_ _35970_/CLK _35518_/D VGND VGND VPWR VPWR _35518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20744_ _33488_/Q _33424_/Q _33360_/Q _33296_/Q _20598_/X _20599_/X VGND VGND VPWR
+ VPWR _20744_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26251_ _25146_/X _33536_/Q _26269_/S VGND VGND VPWR VPWR _26252_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35449_ _35578_/CLK _35449_/D VGND VGND VPWR VPWR _35449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23463_ _22932_/X _32287_/Q _23467_/S VGND VGND VPWR VPWR _23464_/A sky130_fd_sc_hd__mux2_1
X_20675_ _22531_/A VGND VGND VPWR VPWR _20675_/X sky130_fd_sc_hd__buf_6
XFILLER_137_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25202_ _25202_/A VGND VGND VPWR VPWR _33043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22414_ _33215_/Q _32575_/Q _35967_/Q _35903_/Q _22380_/X _22381_/X VGND VGND VPWR
+ VPWR _22414_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26182_ _26182_/A VGND VGND VPWR VPWR _33503_/D sky130_fd_sc_hd__clkbuf_1
X_23394_ _23421_/S VGND VGND VPWR VPWR _23413_/S sky130_fd_sc_hd__buf_4
XFILLER_13_1127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25133_ _25133_/A VGND VGND VPWR VPWR _33019_/D sky130_fd_sc_hd__clkbuf_1
X_22345_ _34813_/Q _34749_/Q _34685_/Q _34621_/Q _22241_/X _22242_/X VGND VGND VPWR
+ VPWR _22345_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29941_ _29941_/A VGND VGND VPWR VPWR _35221_/D sky130_fd_sc_hd__clkbuf_1
X_25064_ _25063_/X _32997_/Q _25082_/S VGND VGND VPWR VPWR _25065_/A sky130_fd_sc_hd__mux2_1
X_22276_ _35323_/Q _35259_/Q _35195_/Q _32315_/Q _21959_/X _21960_/X VGND VGND VPWR
+ VPWR _22276_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24015_ _24015_/A VGND VGND VPWR VPWR _32545_/D sky130_fd_sc_hd__clkbuf_1
X_21227_ _21089_/X _21225_/X _21226_/X _21094_/X VGND VGND VPWR VPWR _21227_/X sky130_fd_sc_hd__a22o_1
X_29872_ _35189_/Q _29172_/X _29872_/S VGND VGND VPWR VPWR _29873_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28823_ _28823_/A VGND VGND VPWR VPWR _34722_/D sky130_fd_sc_hd__clkbuf_1
X_21158_ _21158_/A VGND VGND VPWR VPWR _36187_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20109_ _20105_/X _20108_/X _19789_/X _19790_/X VGND VGND VPWR VPWR _20124_/B sky130_fd_sc_hd__o211a_1
X_28754_ _26984_/X _34690_/Q _28768_/S VGND VGND VPWR VPWR _28755_/A sky130_fd_sc_hd__mux2_1
X_25966_ _25125_/X _33401_/Q _25978_/S VGND VGND VPWR VPWR _25967_/A sky130_fd_sc_hd__mux2_1
X_21089_ _22501_/A VGND VGND VPWR VPWR _21089_/X sky130_fd_sc_hd__buf_4
XFILLER_247_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27705_ _27705_/A VGND VGND VPWR VPWR _34192_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24917_ _24917_/A VGND VGND VPWR VPWR _32939_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25897_ _25022_/X _33368_/Q _25915_/S VGND VGND VPWR VPWR _25898_/A sky130_fd_sc_hd__mux2_1
X_28685_ _28685_/A VGND VGND VPWR VPWR _34657_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27636_ _34160_/Q _24351_/X _27646_/S VGND VGND VPWR VPWR _27637_/A sky130_fd_sc_hd__mux2_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24848_ _23068_/X _32907_/Q _24852_/S VGND VGND VPWR VPWR _24849_/A sky130_fd_sc_hd__mux2_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27567_ _34127_/Q _24249_/X _27583_/S VGND VGND VPWR VPWR _27568_/A sky130_fd_sc_hd__mux2_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24779_ _22966_/X _32874_/Q _24781_/S VGND VGND VPWR VPWR _24780_/A sky130_fd_sc_hd__mux2_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _16999_/X _17318_/X _17319_/X _17002_/X VGND VGND VPWR VPWR _17320_/X sky130_fd_sc_hd__a22o_1
X_29306_ _29306_/A VGND VGND VPWR VPWR _34920_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26518_ _25143_/X _33663_/Q _26518_/S VGND VGND VPWR VPWR _26519_/A sky130_fd_sc_hd__mux2_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27498_ _27498_/A VGND VGND VPWR VPWR _34095_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29237_ input57/X VGND VGND VPWR VPWR _29237_/X sky130_fd_sc_hd__buf_2
XFILLER_35_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17251_ _17957_/A VGND VGND VPWR VPWR _17251_/X sky130_fd_sc_hd__buf_4
XFILLER_230_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26449_ _25041_/X _33630_/Q _26455_/S VGND VGND VPWR VPWR _26450_/A sky130_fd_sc_hd__mux2_1
X_16202_ _16087_/X _16200_/X _16201_/X _16097_/X VGND VGND VPWR VPWR _16202_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17182_ _35565_/Q _35501_/Q _35437_/Q _35373_/Q _16897_/X _16898_/X VGND VGND VPWR
+ VPWR _17182_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29168_ _29168_/A VGND VGND VPWR VPWR _34867_/D sky130_fd_sc_hd__clkbuf_1
X_16133_ _16129_/X _16132_/X _16100_/X VGND VGND VPWR VPWR _16134_/D sky130_fd_sc_hd__o21ba_1
X_28119_ _26844_/X _34389_/Q _28123_/S VGND VGND VPWR VPWR _28120_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29099_ _34845_/Q _29098_/X _29111_/S VGND VGND VPWR VPWR _29100_/A sky130_fd_sc_hd__mux2_1
X_31130_ _35785_/Q _29234_/X _31130_/S VGND VGND VPWR VPWR _31131_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16064_ _17762_/A VGND VGND VPWR VPWR _17932_/A sky130_fd_sc_hd__buf_12
XFILLER_142_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31061_ _35752_/Q _29132_/X _31067_/S VGND VGND VPWR VPWR _31062_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30012_ _35255_/Q _29179_/X _30028_/S VGND VGND VPWR VPWR _30013_/A sky130_fd_sc_hd__mux2_1
X_19823_ _19502_/X _19821_/X _19822_/X _19505_/X VGND VGND VPWR VPWR _19823_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34820_ _35779_/CLK _34820_/D VGND VGND VPWR VPWR _34820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19754_ _33013_/Q _32949_/Q _32885_/Q _32821_/Q _19642_/X _19643_/X VGND VGND VPWR
+ VPWR _19754_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16966_ _33191_/Q _32551_/Q _35943_/Q _35879_/Q _16721_/X _16722_/X VGND VGND VPWR
+ VPWR _16966_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18705_ _34775_/Q _34711_/Q _34647_/Q _34583_/Q _18529_/X _18530_/X VGND VGND VPWR
+ VPWR _18705_/X sky130_fd_sc_hd__mux4_1
XFILLER_231_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34751_ _35837_/CLK _34751_/D VGND VGND VPWR VPWR _34751_/Q sky130_fd_sc_hd__dfxtp_1
X_31963_ _35166_/CLK _31963_/D VGND VGND VPWR VPWR _31963_/Q sky130_fd_sc_hd__dfxtp_1
X_19685_ _35827_/Q _32205_/Q _35699_/Q _35635_/Q _19613_/X _19614_/X VGND VGND VPWR
+ VPWR _19685_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16897_ _17956_/A VGND VGND VPWR VPWR _16897_/X sky130_fd_sc_hd__buf_4
XFILLER_209_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33702_ _33702_/CLK _33702_/D VGND VGND VPWR VPWR _33702_/Q sky130_fd_sc_hd__dfxtp_1
X_18636_ _34517_/Q _32405_/Q _34389_/Q _34325_/Q _18466_/X _18467_/X VGND VGND VPWR
+ VPWR _18636_/X sky130_fd_sc_hd__mux4_1
X_30914_ _35682_/Q _29113_/X _30932_/S VGND VGND VPWR VPWR _30915_/A sky130_fd_sc_hd__mux2_1
XTAP_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34682_ _35771_/CLK _34682_/D VGND VGND VPWR VPWR _34682_/Q sky130_fd_sc_hd__dfxtp_1
X_31894_ _23261_/X _36147_/Q _31898_/S VGND VGND VPWR VPWR _31895_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33633_ _34145_/CLK _33633_/D VGND VGND VPWR VPWR _33633_/Q sky130_fd_sc_hd__dfxtp_1
X_30845_ _30845_/A VGND VGND VPWR VPWR _35649_/D sky130_fd_sc_hd__clkbuf_1
X_18567_ _35027_/Q _34963_/Q _34899_/Q _34835_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _18567_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17518_ _33783_/Q _33719_/Q _33655_/Q _33591_/Q _17196_/X _17197_/X VGND VGND VPWR
+ VPWR _17518_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33564_ _34010_/CLK _33564_/D VGND VGND VPWR VPWR _33564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18498_ _35281_/Q _35217_/Q _35153_/Q _32273_/Q _18379_/X _18381_/X VGND VGND VPWR
+ VPWR _18498_/X sky130_fd_sc_hd__mux4_1
X_30776_ _23145_/X _35617_/Q _30776_/S VGND VGND VPWR VPWR _30777_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35303_ _35303_/CLK _35303_/D VGND VGND VPWR VPWR _35303_/Q sky130_fd_sc_hd__dfxtp_1
X_32515_ _36037_/CLK _32515_/D VGND VGND VPWR VPWR _32515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17449_ _17445_/X _17448_/X _17128_/X VGND VGND VPWR VPWR _17471_/A sky130_fd_sc_hd__o21ba_1
X_33495_ _34001_/CLK _33495_/D VGND VGND VPWR VPWR _33495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35234_ _35298_/CLK _35234_/D VGND VGND VPWR VPWR _35234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20460_ _20208_/X _20458_/X _20459_/X _20211_/X VGND VGND VPWR VPWR _20460_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32446_ _35581_/CLK _32446_/D VGND VGND VPWR VPWR _32446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19119_ _32739_/Q _32675_/Q _32611_/Q _36067_/Q _18866_/X _19003_/X VGND VGND VPWR
+ VPWR _19119_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35165_ _35293_/CLK _35165_/D VGND VGND VPWR VPWR _35165_/Q sky130_fd_sc_hd__dfxtp_1
X_20391_ _20160_/X _20389_/X _20390_/X _20165_/X VGND VGND VPWR VPWR _20391_/X sky130_fd_sc_hd__a22o_1
XFILLER_203_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32377_ _36025_/CLK _32377_/D VGND VGND VPWR VPWR _32377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34116_ _34308_/CLK _34116_/D VGND VGND VPWR VPWR _34116_/Q sky130_fd_sc_hd__dfxtp_1
X_22130_ _22016_/X _22128_/X _22129_/X _22020_/X VGND VGND VPWR VPWR _22130_/X sky130_fd_sc_hd__a22o_1
X_31328_ _31328_/A VGND VGND VPWR VPWR _35878_/D sky130_fd_sc_hd__clkbuf_1
Xoutput210 _36234_/Q VGND VGND VPWR VPWR D2[60] sky130_fd_sc_hd__buf_2
X_35096_ _35738_/CLK _35096_/D VGND VGND VPWR VPWR _35096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput221 _32090_/Q VGND VGND VPWR VPWR D3[12] sky130_fd_sc_hd__buf_2
XFILLER_245_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput232 _32100_/Q VGND VGND VPWR VPWR D3[22] sky130_fd_sc_hd__buf_2
XFILLER_86_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34047_ _34303_/CLK _34047_/D VGND VGND VPWR VPWR _34047_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput243 _32110_/Q VGND VGND VPWR VPWR D3[32] sky130_fd_sc_hd__buf_2
X_22061_ _33205_/Q _32565_/Q _35957_/Q _35893_/Q _22027_/X _22028_/X VGND VGND VPWR
+ VPWR _22061_/X sky130_fd_sc_hd__mux4_1
XTAP_6609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31259_ _35846_/Q input52/X _31265_/S VGND VGND VPWR VPWR _31260_/A sky130_fd_sc_hd__mux2_1
Xoutput254 _32120_/Q VGND VGND VPWR VPWR D3[42] sky130_fd_sc_hd__buf_2
XFILLER_99_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput265 _32130_/Q VGND VGND VPWR VPWR D3[52] sky130_fd_sc_hd__buf_2
Xoutput276 _32140_/Q VGND VGND VPWR VPWR D3[62] sky130_fd_sc_hd__buf_2
X_21012_ _21012_/A _21012_/B _21012_/C _21012_/D VGND VGND VPWR VPWR _21013_/A sky130_fd_sc_hd__or4_1
XFILLER_138_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25820_ _25109_/X _33332_/Q _25822_/S VGND VGND VPWR VPWR _25821_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35998_ _36062_/CLK _35998_/D VGND VGND VPWR VPWR _35998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25751_ _25007_/X _33299_/Q _25759_/S VGND VGND VPWR VPWR _25752_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34949_ _35781_/CLK _34949_/D VGND VGND VPWR VPWR _34949_/Q sky130_fd_sc_hd__dfxtp_1
X_22963_ input20/X VGND VGND VPWR VPWR _22963_/X sky130_fd_sc_hd__clkbuf_4
X_24702_ _24702_/A VGND VGND VPWR VPWR _32838_/D sky130_fd_sc_hd__clkbuf_1
X_21914_ _22396_/A VGND VGND VPWR VPWR _21914_/X sky130_fd_sc_hd__buf_4
X_28470_ _28470_/A VGND VGND VPWR VPWR _34555_/D sky130_fd_sc_hd__clkbuf_1
X_25682_ _25682_/A VGND VGND VPWR VPWR _33267_/D sky130_fd_sc_hd__clkbuf_1
X_22894_ _22894_/A VGND VGND VPWR VPWR _32018_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27421_ _27421_/A VGND VGND VPWR VPWR _34059_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24633_ _24633_/A VGND VGND VPWR VPWR _32805_/D sky130_fd_sc_hd__clkbuf_1
X_21845_ _21663_/X _21843_/X _21844_/X _21667_/X VGND VGND VPWR VPWR _21845_/X sky130_fd_sc_hd__a22o_1
XFILLER_203_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24564_ _24564_/A VGND VGND VPWR VPWR _32774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27352_ _27352_/A VGND VGND VPWR VPWR _34026_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21776_ _33005_/Q _32941_/Q _32877_/Q _32813_/Q _21589_/X _21590_/X VGND VGND VPWR
+ VPWR _21776_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26303_ _26303_/A VGND VGND VPWR VPWR _33560_/D sky130_fd_sc_hd__clkbuf_1
X_23515_ _23515_/A VGND VGND VPWR VPWR _32311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27283_ _27008_/X _33994_/Q _27289_/S VGND VGND VPWR VPWR _27284_/A sky130_fd_sc_hd__mux2_1
X_20727_ _34767_/Q _34703_/Q _34639_/Q _34575_/Q _20675_/X _20676_/X VGND VGND VPWR
+ VPWR _20727_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24495_ _24495_/A VGND VGND VPWR VPWR _32741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29022_ _34817_/Q _24404_/X _29038_/S VGND VGND VPWR VPWR _29023_/A sky130_fd_sc_hd__mux2_1
X_26234_ _25122_/X _33528_/Q _26248_/S VGND VGND VPWR VPWR _26235_/A sky130_fd_sc_hd__mux2_1
X_23446_ _22907_/X _32279_/Q _23446_/S VGND VGND VPWR VPWR _23447_/A sky130_fd_sc_hd__mux2_1
X_20658_ _22446_/A VGND VGND VPWR VPWR _20658_/X sky130_fd_sc_hd__buf_8
XFILLER_149_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26165_ _26165_/A VGND VGND VPWR VPWR _33495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23377_ _23377_/A VGND VGND VPWR VPWR _32247_/D sky130_fd_sc_hd__clkbuf_1
X_20589_ _22395_/A VGND VGND VPWR VPWR _20589_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25116_ _25187_/S VGND VGND VPWR VPWR _25144_/S sky130_fd_sc_hd__buf_4
X_22328_ _34045_/Q _33981_/Q _33917_/Q _32253_/Q _22326_/X _22327_/X VGND VGND VPWR
+ VPWR _22328_/X sky130_fd_sc_hd__mux4_1
X_26096_ _26096_/A VGND VGND VPWR VPWR _33462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_944 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29924_ _29924_/A _30059_/A VGND VGND VPWR VPWR _30057_/S sky130_fd_sc_hd__nor2_8
XFILLER_139_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25047_ input10/X VGND VGND VPWR VPWR _25047_/X sky130_fd_sc_hd__clkbuf_4
X_22259_ _32763_/Q _32699_/Q _32635_/Q _36091_/Q _22225_/X _22009_/X VGND VGND VPWR
+ VPWR _22259_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29855_ _29855_/A VGND VGND VPWR VPWR _35180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28806_ _28806_/A VGND VGND VPWR VPWR _34714_/D sky130_fd_sc_hd__clkbuf_1
X_16820_ _33251_/Q _36131_/Q _33123_/Q _33059_/Q _16705_/X _16706_/X VGND VGND VPWR
+ VPWR _16820_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29786_ _29786_/A VGND VGND VPWR VPWR _35148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26998_ _26998_/A VGND VGND VPWR VPWR _33862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28737_ _26959_/X _34682_/Q _28747_/S VGND VGND VPWR VPWR _28738_/A sky130_fd_sc_hd__mux2_1
X_16751_ _35809_/Q _32185_/Q _35681_/Q _35617_/Q _16607_/X _16608_/X VGND VGND VPWR
+ VPWR _16751_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_1136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25949_ _25100_/X _33393_/Q _25957_/S VGND VGND VPWR VPWR _25950_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19470_ _19149_/X _19468_/X _19469_/X _19152_/X VGND VGND VPWR VPWR _19470_/X sky130_fd_sc_hd__a22o_1
XFILLER_234_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16682_ _35551_/Q _35487_/Q _35423_/Q _35359_/Q _16544_/X _16545_/X VGND VGND VPWR
+ VPWR _16682_/X sky130_fd_sc_hd__mux4_1
X_28668_ _26857_/X _34649_/Q _28684_/S VGND VGND VPWR VPWR _28669_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18421_ _35727_/Q _35087_/Q _34447_/Q _33807_/Q _18349_/X _18351_/X VGND VGND VPWR
+ VPWR _18421_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27619_ _34152_/Q _24326_/X _27625_/S VGND VGND VPWR VPWR _27620_/A sky130_fd_sc_hd__mux2_1
XFILLER_234_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28599_ _28599_/A VGND VGND VPWR VPWR _34616_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18352_ _35726_/Q _35086_/Q _34446_/Q _33806_/Q _18349_/X _18351_/X VGND VGND VPWR
+ VPWR _18352_/X sky130_fd_sc_hd__mux4_1
X_30630_ _30630_/A VGND VGND VPWR VPWR _35547_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _34033_/Q _33969_/Q _33905_/Q _32241_/Q _17020_/X _17021_/X VGND VGND VPWR
+ VPWR _17303_/X sky130_fd_sc_hd__mux4_1
X_18283_ _20203_/A VGND VGND VPWR VPWR _18283_/X sky130_fd_sc_hd__buf_6
X_30561_ _23286_/X _35515_/Q _30569_/S VGND VGND VPWR VPWR _30562_/A sky130_fd_sc_hd__mux2_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32300_ _35564_/CLK _32300_/D VGND VGND VPWR VPWR _32300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17234_ _34287_/Q _34223_/Q _34159_/Q _34095_/Q _17089_/X _17090_/X VGND VGND VPWR
+ VPWR _17234_/X sky130_fd_sc_hd__mux4_1
X_33280_ _36160_/CLK _33280_/D VGND VGND VPWR VPWR _33280_/Q sky130_fd_sc_hd__dfxtp_1
X_30492_ _23124_/X _35482_/Q _30506_/S VGND VGND VPWR VPWR _30493_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32231_ _35787_/CLK _32231_/D VGND VGND VPWR VPWR _32231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17165_ _33773_/Q _33709_/Q _33645_/Q _33581_/Q _16843_/X _16844_/X VGND VGND VPWR
+ VPWR _17165_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16116_ _32463_/Q _32335_/Q _32015_/Q _35983_/Q _16028_/X _17863_/A VGND VGND VPWR
+ VPWR _16116_/X sky130_fd_sc_hd__mux4_1
X_32162_ _36130_/CLK _32162_/D VGND VGND VPWR VPWR _32162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17096_ _17092_/X _17095_/X _16775_/X VGND VGND VPWR VPWR _17118_/A sky130_fd_sc_hd__o21ba_1
XFILLER_127_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31113_ _31113_/A VGND VGND VPWR VPWR _35776_/D sky130_fd_sc_hd__clkbuf_1
X_16047_ _35790_/Q _32164_/Q _35662_/Q _35598_/Q _16045_/X _16046_/X VGND VGND VPWR
+ VPWR _16047_/X sky130_fd_sc_hd__mux4_1
XFILLER_115_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32093_ _35807_/CLK _32093_/D VGND VGND VPWR VPWR _32093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35921_ _35921_/CLK _35921_/D VGND VGND VPWR VPWR _35921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31044_ _35744_/Q _29107_/X _31046_/S VGND VGND VPWR VPWR _31045_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19806_ _19802_/X _19803_/X _19804_/X _19805_/X VGND VGND VPWR VPWR _19806_/X sky130_fd_sc_hd__a22o_1
X_35852_ _35852_/CLK _35852_/D VGND VGND VPWR VPWR _35852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17998_ _17855_/X _17996_/X _17997_/X _17858_/X VGND VGND VPWR VPWR _17998_/X sky130_fd_sc_hd__a22o_1
X_34803_ _35250_/CLK _34803_/D VGND VGND VPWR VPWR _34803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19737_ _19454_/X _19735_/X _19736_/X _19459_/X VGND VGND VPWR VPWR _19737_/X sky130_fd_sc_hd__a22o_1
X_35783_ _35845_/CLK _35783_/D VGND VGND VPWR VPWR _35783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16949_ _33511_/Q _33447_/Q _33383_/Q _33319_/Q _16770_/X _16771_/X VGND VGND VPWR
+ VPWR _16949_/X sky130_fd_sc_hd__mux4_1
X_32995_ _36067_/CLK _32995_/D VGND VGND VPWR VPWR _32995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34734_ _35308_/CLK _34734_/D VGND VGND VPWR VPWR _34734_/Q sky130_fd_sc_hd__dfxtp_1
X_31946_ _23342_/X _36172_/Q _31948_/S VGND VGND VPWR VPWR _31947_/A sky130_fd_sc_hd__mux2_1
X_19668_ _19668_/A VGND VGND VPWR VPWR _32114_/D sky130_fd_sc_hd__buf_2
XFILLER_237_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18619_ _32725_/Q _32661_/Q _32597_/Q _36053_/Q _18513_/X _20013_/A VGND VGND VPWR
+ VPWR _18619_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34665_ _34792_/CLK _34665_/D VGND VGND VPWR VPWR _34665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19599_ _33777_/Q _33713_/Q _33649_/Q _33585_/Q _19496_/X _19497_/X VGND VGND VPWR
+ VPWR _19599_/X sky130_fd_sc_hd__mux4_1
X_31877_ _23234_/X _36139_/Q _31877_/S VGND VGND VPWR VPWR _31878_/A sky130_fd_sc_hd__mux2_1
X_33616_ _34194_/CLK _33616_/D VGND VGND VPWR VPWR _33616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_1221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_39__f_CLK clkbuf_5_19_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_39__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_21630_ _21310_/X _21628_/X _21629_/X _21314_/X VGND VGND VPWR VPWR _21630_/X sky130_fd_sc_hd__a22o_1
X_30828_ _30828_/A VGND VGND VPWR VPWR _35641_/D sky130_fd_sc_hd__clkbuf_1
X_34596_ _35928_/CLK _34596_/D VGND VGND VPWR VPWR _34596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33547_ _36041_/CLK _33547_/D VGND VGND VPWR VPWR _33547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21561_ _22396_/A VGND VGND VPWR VPWR _21561_/X sky130_fd_sc_hd__buf_4
XFILLER_244_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30759_ _30759_/A VGND VGND VPWR VPWR _35608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23300_ input44/X VGND VGND VPWR VPWR _23300_/X sky130_fd_sc_hd__buf_4
XFILLER_60_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20512_ _20508_/X _20511_/X _20167_/A VGND VGND VPWR VPWR _20513_/D sky130_fd_sc_hd__o21ba_1
XFILLER_193_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24280_ input3/X VGND VGND VPWR VPWR _24280_/X sky130_fd_sc_hd__buf_4
X_33478_ _34053_/CLK _33478_/D VGND VGND VPWR VPWR _33478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21492_ _21310_/X _21490_/X _21491_/X _21314_/X VGND VGND VPWR VPWR _21492_/X sky130_fd_sc_hd__a22o_1
XFILLER_197_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35217_ _36216_/CLK _35217_/D VGND VGND VPWR VPWR _35217_/Q sky130_fd_sc_hd__dfxtp_1
X_23231_ input21/X VGND VGND VPWR VPWR _23231_/X sky130_fd_sc_hd__buf_4
X_20443_ _33225_/Q _32585_/Q _35977_/Q _35913_/Q _18375_/X _18376_/X VGND VGND VPWR
+ VPWR _20443_/X sky130_fd_sc_hd__mux4_1
X_32429_ _35500_/CLK _32429_/D VGND VGND VPWR VPWR _32429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36197_ _36200_/CLK _36197_/D VGND VGND VPWR VPWR _36197_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_101_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35148_ _35853_/CLK _35148_/D VGND VGND VPWR VPWR _35148_/Q sky130_fd_sc_hd__dfxtp_1
X_23162_ _23162_/A VGND VGND VPWR VPWR _32164_/D sky130_fd_sc_hd__clkbuf_1
X_20374_ _20061_/X _20372_/X _20373_/X _20067_/X VGND VGND VPWR VPWR _20374_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22113_ _22107_/X _22108_/X _22111_/X _22112_/X VGND VGND VPWR VPWR _22113_/X sky130_fd_sc_hd__a22o_1
XTAP_7129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35079_ _35079_/CLK _35079_/D VGND VGND VPWR VPWR _35079_/Q sky130_fd_sc_hd__dfxtp_1
X_27970_ _26821_/X _34318_/Q _27988_/S VGND VGND VPWR VPWR _27971_/A sky130_fd_sc_hd__mux2_1
X_23093_ input23/X VGND VGND VPWR VPWR _23093_/X sky130_fd_sc_hd__buf_4
XTAP_6406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26921_ _26921_/A VGND VGND VPWR VPWR _33837_/D sky130_fd_sc_hd__clkbuf_1
X_22044_ _34293_/Q _34229_/Q _34165_/Q _34101_/Q _22042_/X _22043_/X VGND VGND VPWR
+ VPWR _22044_/X sky130_fd_sc_hd__mux4_1
XTAP_6439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29640_ _35079_/Q _29228_/X _29644_/S VGND VGND VPWR VPWR _29641_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_1389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26852_ _26852_/A VGND VGND VPWR VPWR _33815_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25803_ _25872_/S VGND VGND VPWR VPWR _25822_/S sky130_fd_sc_hd__buf_4
XFILLER_214_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29571_ _35046_/Q _29126_/X _29581_/S VGND VGND VPWR VPWR _29572_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26783_ _26783_/A VGND VGND VPWR VPWR _33787_/D sky130_fd_sc_hd__clkbuf_1
X_23995_ _24106_/S VGND VGND VPWR VPWR _24014_/S sky130_fd_sc_hd__buf_4
XFILLER_169_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28522_ _26841_/X _34580_/Q _28528_/S VGND VGND VPWR VPWR _28523_/A sky130_fd_sc_hd__mux2_1
X_25734_ _25734_/A VGND VGND VPWR VPWR _33292_/D sky130_fd_sc_hd__clkbuf_1
X_22946_ _22945_/X _32035_/Q _22970_/S VGND VGND VPWR VPWR _22947_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28453_ _28453_/A VGND VGND VPWR VPWR _34547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22877_ input88/X input87/X input86/X input89/X VGND VGND VPWR VPWR _23561_/B sky130_fd_sc_hd__and4_2
XFILLER_141_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25665_ _25665_/A VGND VGND VPWR VPWR _33259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27404_ _34051_/Q _24410_/X _27416_/S VGND VGND VPWR VPWR _27405_/A sky130_fd_sc_hd__mux2_1
X_21828_ _35054_/Q _34990_/Q _34926_/Q _34862_/Q _21756_/X _21757_/X VGND VGND VPWR
+ VPWR _21828_/X sky130_fd_sc_hd__mux4_1
X_24616_ _24616_/A VGND VGND VPWR VPWR _32797_/D sky130_fd_sc_hd__clkbuf_1
X_25596_ _25596_/A VGND VGND VPWR VPWR _33228_/D sky130_fd_sc_hd__clkbuf_1
X_28384_ _28384_/A VGND VGND VPWR VPWR _34514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24547_ _24547_/A VGND VGND VPWR VPWR _32766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27335_ _34018_/Q _24307_/X _27353_/S VGND VGND VPWR VPWR _27336_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21759_ _21759_/A VGND VGND VPWR VPWR _21759_/X sky130_fd_sc_hd__buf_4
XFILLER_19_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27266_ _27266_/A VGND VGND VPWR VPWR _33985_/D sky130_fd_sc_hd__clkbuf_1
X_24478_ _24478_/A VGND VGND VPWR VPWR _32733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29005_ _34809_/Q _24379_/X _29017_/S VGND VGND VPWR VPWR _29006_/A sky130_fd_sc_hd__mux2_1
X_23429_ _23429_/A VGND VGND VPWR VPWR _32270_/D sky130_fd_sc_hd__clkbuf_1
X_26217_ _25097_/X _33520_/Q _26227_/S VGND VGND VPWR VPWR _26218_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27197_ _26881_/X _33953_/Q _27197_/S VGND VGND VPWR VPWR _27198_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26148_ _24995_/X _33487_/Q _26164_/S VGND VGND VPWR VPWR _26149_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26079_ _26079_/A VGND VGND VPWR VPWR _33454_/D sky130_fd_sc_hd__clkbuf_1
X_18970_ _18796_/X _18966_/X _18969_/X _18799_/X VGND VGND VPWR VPWR _18970_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29907_ _29907_/A VGND VGND VPWR VPWR _35205_/D sky130_fd_sc_hd__clkbuf_1
X_17921_ _35842_/Q _32221_/Q _35714_/Q _35650_/Q _17666_/X _17667_/X VGND VGND VPWR
+ VPWR _17921_/X sky130_fd_sc_hd__mux4_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17852_ _17705_/X _17850_/X _17851_/X _17708_/X VGND VGND VPWR VPWR _17852_/X sky130_fd_sc_hd__a22o_1
X_29838_ _29838_/A VGND VGND VPWR VPWR _35172_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16803_ _17862_/A VGND VGND VPWR VPWR _16803_/X sky130_fd_sc_hd__clkbuf_8
X_29769_ _35140_/Q _29219_/X _29779_/S VGND VGND VPWR VPWR _29770_/A sky130_fd_sc_hd__mux2_1
X_17783_ _17705_/X _17779_/X _17782_/X _17708_/X VGND VGND VPWR VPWR _17783_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31800_ _31800_/A VGND VGND VPWR VPWR _36102_/D sky130_fd_sc_hd__clkbuf_1
X_19522_ _34798_/Q _34734_/Q _34670_/Q _34606_/Q _19235_/X _19236_/X VGND VGND VPWR
+ VPWR _19522_/X sky130_fd_sc_hd__mux4_1
X_16734_ _16734_/A VGND VGND VPWR VPWR _31968_/D sky130_fd_sc_hd__clkbuf_1
X_32780_ _36109_/CLK _32780_/D VGND VGND VPWR VPWR _32780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19453_ _19449_/X _19450_/X _19451_/X _19452_/X VGND VGND VPWR VPWR _19453_/X sky130_fd_sc_hd__a22o_1
X_31731_ _31731_/A VGND VGND VPWR VPWR _36069_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16665_ _16489_/X _16663_/X _16664_/X _16494_/X VGND VGND VPWR VPWR _16665_/X sky130_fd_sc_hd__a22o_1
XFILLER_228_1238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18404_ _33743_/Q _33679_/Q _33615_/Q _33551_/Q _18280_/X _18283_/X VGND VGND VPWR
+ VPWR _18404_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34450_ _35729_/CLK _34450_/D VGND VGND VPWR VPWR _34450_/Q sky130_fd_sc_hd__dfxtp_1
X_31662_ _36037_/Q input51/X _31670_/S VGND VGND VPWR VPWR _31663_/A sky130_fd_sc_hd__mux2_1
X_19384_ _19101_/X _19382_/X _19383_/X _19106_/X VGND VGND VPWR VPWR _19384_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16596_ _33501_/Q _33437_/Q _33373_/Q _33309_/Q _16417_/X _16418_/X VGND VGND VPWR
+ VPWR _16596_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33401_ _34298_/CLK _33401_/D VGND VGND VPWR VPWR _33401_/Q sky130_fd_sc_hd__dfxtp_1
X_30613_ _30613_/A VGND VGND VPWR VPWR _35539_/D sky130_fd_sc_hd__clkbuf_1
X_18335_ _20130_/A VGND VGND VPWR VPWR _18335_/X sky130_fd_sc_hd__clkbuf_4
X_34381_ _35597_/CLK _34381_/D VGND VGND VPWR VPWR _34381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31593_ _36004_/Q input15/X _31607_/S VGND VGND VPWR VPWR _31594_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36120_ _36123_/CLK _36120_/D VGND VGND VPWR VPWR _36120_/Q sky130_fd_sc_hd__dfxtp_1
X_33332_ _33780_/CLK _33332_/D VGND VGND VPWR VPWR _33332_/Q sky130_fd_sc_hd__dfxtp_1
X_18266_ _34829_/Q _34765_/Q _34701_/Q _34637_/Q _17994_/X _17995_/X VGND VGND VPWR
+ VPWR _18266_/X sky130_fd_sc_hd__mux4_1
X_30544_ _23261_/X _35507_/Q _30548_/S VGND VGND VPWR VPWR _30545_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36051_ _36052_/CLK _36051_/D VGND VGND VPWR VPWR _36051_/Q sky130_fd_sc_hd__dfxtp_1
X_17217_ _16994_/X _17215_/X _17216_/X _16997_/X VGND VGND VPWR VPWR _17217_/X sky130_fd_sc_hd__a22o_1
X_33263_ _36081_/CLK _33263_/D VGND VGND VPWR VPWR _33263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18197_ _17154_/A _18195_/X _18196_/X _17159_/A VGND VGND VPWR VPWR _18197_/X sky130_fd_sc_hd__a22o_1
X_30475_ _23099_/X _35474_/Q _30485_/S VGND VGND VPWR VPWR _30476_/A sky130_fd_sc_hd__mux2_1
X_35002_ _35002_/CLK _35002_/D VGND VGND VPWR VPWR _35002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32214_ _35965_/CLK _32214_/D VGND VGND VPWR VPWR _32214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17148_ _17143_/X _17146_/X _17147_/X VGND VGND VPWR VPWR _17163_/C sky130_fd_sc_hd__o21ba_1
X_33194_ _35946_/CLK _33194_/D VGND VGND VPWR VPWR _33194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32145_ _36228_/CLK _32145_/D VGND VGND VPWR VPWR _32145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17079_ _34794_/Q _34730_/Q _34666_/Q _34602_/Q _16935_/X _16936_/X VGND VGND VPWR
+ VPWR _17079_/X sky130_fd_sc_hd__mux4_1
XFILLER_171_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32076_ _35532_/CLK _32076_/D VGND VGND VPWR VPWR _32076_/Q sky130_fd_sc_hd__dfxtp_1
X_20090_ _19807_/X _20088_/X _20089_/X _19812_/X VGND VGND VPWR VPWR _20090_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_830 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35904_ _35971_/CLK _35904_/D VGND VGND VPWR VPWR _35904_/Q sky130_fd_sc_hd__dfxtp_1
X_31027_ _31138_/S VGND VGND VPWR VPWR _31046_/S sky130_fd_sc_hd__buf_4
XFILLER_242_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35835_ _35965_/CLK _35835_/D VGND VGND VPWR VPWR _35835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22800_ _35787_/Q _35147_/Q _34507_/Q _33867_/Q _20708_/X _20709_/X VGND VGND VPWR
+ VPWR _22800_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23780_ _22994_/X _32435_/Q _23784_/S VGND VGND VPWR VPWR _23781_/A sky130_fd_sc_hd__mux2_1
X_32978_ _32978_/CLK _32978_/D VGND VGND VPWR VPWR _32978_/Q sky130_fd_sc_hd__dfxtp_1
X_20992_ _33239_/Q _36119_/Q _33111_/Q _33047_/Q _20952_/X _20953_/X VGND VGND VPWR
+ VPWR _20992_/X sky130_fd_sc_hd__mux4_1
X_35766_ _35766_/CLK _35766_/D VGND VGND VPWR VPWR _35766_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22731_ _22727_/X _22730_/X _22434_/X VGND VGND VPWR VPWR _22753_/A sky130_fd_sc_hd__o21ba_2
X_31929_ _31929_/A VGND VGND VPWR VPWR _36163_/D sky130_fd_sc_hd__clkbuf_1
X_34717_ _35034_/CLK _34717_/D VGND VGND VPWR VPWR _34717_/Q sky130_fd_sc_hd__dfxtp_1
X_35697_ _35954_/CLK _35697_/D VGND VGND VPWR VPWR _35697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25450_ _25174_/X _33161_/Q _25450_/S VGND VGND VPWR VPWR _25451_/A sky130_fd_sc_hd__mux2_1
X_22662_ _22658_/X _22661_/X _22467_/X VGND VGND VPWR VPWR _22663_/D sky130_fd_sc_hd__o21ba_1
X_34648_ _34777_/CLK _34648_/D VGND VGND VPWR VPWR _34648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24401_ _24401_/A VGND VGND VPWR VPWR _24429_/S sky130_fd_sc_hd__buf_6
XFILLER_80_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21613_ _21609_/X _21612_/X _21408_/X VGND VGND VPWR VPWR _21614_/D sky130_fd_sc_hd__o21ba_1
XFILLER_197_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25381_ _25072_/X _33128_/Q _25387_/S VGND VGND VPWR VPWR _25382_/A sky130_fd_sc_hd__mux2_1
X_22593_ _22589_/X _22592_/X _22453_/X VGND VGND VPWR VPWR _22603_/C sky130_fd_sc_hd__o21ba_1
X_34579_ _36189_/CLK _34579_/D VGND VGND VPWR VPWR _34579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27120_ _27120_/A VGND VGND VPWR VPWR _33916_/D sky130_fd_sc_hd__clkbuf_1
X_24332_ input21/X VGND VGND VPWR VPWR _24332_/X sky130_fd_sc_hd__buf_4
XFILLER_181_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21544_ _21544_/A _21544_/B _21544_/C _21544_/D VGND VGND VPWR VPWR _21545_/A sky130_fd_sc_hd__or4_4
X_27051_ _27051_/A VGND VGND VPWR VPWR _33883_/D sky130_fd_sc_hd__clkbuf_1
X_24263_ _24263_/A VGND VGND VPWR VPWR _32659_/D sky130_fd_sc_hd__clkbuf_1
X_21475_ _35044_/Q _34980_/Q _34916_/Q _34852_/Q _21403_/X _21404_/X VGND VGND VPWR
+ VPWR _21475_/X sky130_fd_sc_hd__mux4_1
XFILLER_217_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26002_ _26002_/A VGND VGND VPWR VPWR _33418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23214_ _23214_/A VGND VGND VPWR VPWR _32188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20426_ _34313_/Q _34249_/Q _34185_/Q _34121_/Q _18345_/X _18346_/X VGND VGND VPWR
+ VPWR _20426_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24194_ _24242_/S VGND VGND VPWR VPWR _24213_/S sky130_fd_sc_hd__buf_4
XFILLER_140_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23145_ input11/X VGND VGND VPWR VPWR _23145_/X sky130_fd_sc_hd__buf_4
X_20357_ _35334_/Q _35270_/Q _35206_/Q _32326_/Q _18388_/X _18390_/X VGND VGND VPWR
+ VPWR _20357_/X sky130_fd_sc_hd__mux4_1
XFILLER_218_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27953_ _27953_/A VGND VGND VPWR VPWR _34310_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23076_ _23076_/A VGND VGND VPWR VPWR _32077_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_1009 _17908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20288_ _35780_/Q _35140_/Q _34500_/Q _33860_/Q _20146_/X _20147_/X VGND VGND VPWR
+ VPWR _20288_/X sky130_fd_sc_hd__mux4_1
XTAP_6236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26904_ _26903_/X _33832_/Q _26913_/S VGND VGND VPWR VPWR _26905_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22027_ _22531_/A VGND VGND VPWR VPWR _22027_/X sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_130_CLK clkbuf_6_23__f_CLK/X VGND VGND VPWR VPWR _34194_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27884_ _27884_/A VGND VGND VPWR VPWR _34277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29623_ _35071_/Q _29203_/X _29623_/S VGND VGND VPWR VPWR _29624_/A sky130_fd_sc_hd__mux2_1
XTAP_5568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26835_ input45/X VGND VGND VPWR VPWR _26835_/X sky130_fd_sc_hd__buf_4
XFILLER_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29554_ _35038_/Q _29101_/X _29560_/S VGND VGND VPWR VPWR _29555_/A sky130_fd_sc_hd__mux2_1
XTAP_4878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26766_ _26766_/A VGND VGND VPWR VPWR _33779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23978_ _23978_/A VGND VGND VPWR VPWR _32527_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28505_ _28505_/A VGND VGND VPWR VPWR _34572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25717_ _33284_/Q _24413_/X _25727_/S VGND VGND VPWR VPWR _25718_/A sky130_fd_sc_hd__mux2_1
X_29485_ _29485_/A VGND VGND VPWR VPWR _35005_/D sky130_fd_sc_hd__clkbuf_1
X_22929_ input8/X VGND VGND VPWR VPWR _22929_/X sky130_fd_sc_hd__buf_4
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26697_ _26697_/A VGND VGND VPWR VPWR _33746_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28436_ _28436_/A VGND VGND VPWR VPWR _34539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16450_ _17862_/A VGND VGND VPWR VPWR _16450_/X sky130_fd_sc_hd__buf_4
XFILLER_16_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25648_ _33251_/Q _24311_/X _25664_/S VGND VGND VPWR VPWR _25649_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28367_ _34507_/Q _24434_/X _28371_/S VGND VGND VPWR VPWR _28368_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_6_22__f_CLK clkbuf_5_11_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_22__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_197_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _35966_/CLK sky130_fd_sc_hd__clkbuf_16
X_16381_ _16381_/A VGND VGND VPWR VPWR _31958_/D sky130_fd_sc_hd__clkbuf_1
X_25579_ _33220_/Q _24413_/X _25589_/S VGND VGND VPWR VPWR _25580_/A sky130_fd_sc_hd__mux2_1
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18120_ _35080_/Q _35016_/Q _34952_/Q _34888_/Q _17862_/X _17863_/X VGND VGND VPWR
+ VPWR _18120_/X sky130_fd_sc_hd__mux4_1
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27318_ _34010_/Q _24283_/X _27332_/S VGND VGND VPWR VPWR _27319_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28298_ _34474_/Q _24332_/X _28300_/S VGND VGND VPWR VPWR _28299_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18051_ _15977_/X _18049_/X _18050_/X _15987_/X VGND VGND VPWR VPWR _18051_/X sky130_fd_sc_hd__a22o_1
XFILLER_200_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27249_ _27249_/A VGND VGND VPWR VPWR _33977_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17002_ _17865_/A VGND VGND VPWR VPWR _17002_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_6_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30260_ _30260_/A VGND VGND VPWR VPWR _35372_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_6 _32114_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30191_ _30191_/A VGND VGND VPWR VPWR _35340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18953_ _20012_/A VGND VGND VPWR VPWR _18953_/X sky130_fd_sc_hd__buf_6
XFILLER_193_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_969 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17904_ _33794_/Q _33730_/Q _33666_/Q _33602_/Q _17902_/X _17903_/X VGND VGND VPWR
+ VPWR _17904_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33950_ _34205_/CLK _33950_/D VGND VGND VPWR VPWR _33950_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_121_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _36232_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18884_ _34780_/Q _34716_/Q _34652_/Q _34588_/Q _18882_/X _18883_/X VGND VGND VPWR
+ VPWR _18884_/X sky130_fd_sc_hd__mux4_1
XTAP_6770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32901_ _32901_/CLK _32901_/D VGND VGND VPWR VPWR _32901_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17835_ _17828_/X _17833_/X _17834_/X VGND VGND VPWR VPWR _17869_/A sky130_fd_sc_hd__o21ba_1
XFILLER_86_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33881_ _35284_/CLK _33881_/D VGND VGND VPWR VPWR _33881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32832_ _32962_/CLK _32832_/D VGND VGND VPWR VPWR _32832_/Q sky130_fd_sc_hd__dfxtp_1
X_35620_ _35811_/CLK _35620_/D VGND VGND VPWR VPWR _35620_/Q sky130_fd_sc_hd__dfxtp_1
X_17766_ _33278_/Q _36158_/Q _33150_/Q _33086_/Q _17764_/X _17765_/X VGND VGND VPWR
+ VPWR _17766_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_920 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19505_ _20211_/A VGND VGND VPWR VPWR _19505_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_235_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35551_ _35744_/CLK _35551_/D VGND VGND VPWR VPWR _35551_/Q sky130_fd_sc_hd__dfxtp_1
X_16717_ _35808_/Q _32184_/Q _35680_/Q _35616_/Q _16607_/X _16608_/X VGND VGND VPWR
+ VPWR _16717_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32763_ _33083_/CLK _32763_/D VGND VGND VPWR VPWR _32763_/Q sky130_fd_sc_hd__dfxtp_1
X_17697_ _33020_/Q _32956_/Q _32892_/Q _32828_/Q _17695_/X _17696_/X VGND VGND VPWR
+ VPWR _17697_/X sky130_fd_sc_hd__mux4_1
X_34502_ _35784_/CLK _34502_/D VGND VGND VPWR VPWR _34502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19436_ _20142_/A VGND VGND VPWR VPWR _19436_/X sky130_fd_sc_hd__clkbuf_4
X_31714_ _31714_/A VGND VGND VPWR VPWR _36061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16648_ _33182_/Q _32542_/Q _35934_/Q _35870_/Q _16368_/X _16369_/X VGND VGND VPWR
+ VPWR _16648_/X sky130_fd_sc_hd__mux4_1
X_35482_ _35801_/CLK _35482_/D VGND VGND VPWR VPWR _35482_/Q sky130_fd_sc_hd__dfxtp_1
X_32694_ _36087_/CLK _32694_/D VGND VGND VPWR VPWR _32694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34433_ _36038_/CLK _34433_/D VGND VGND VPWR VPWR _34433_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_188_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _35517_/CLK sky130_fd_sc_hd__clkbuf_16
X_31645_ _36029_/Q input42/X _31649_/S VGND VGND VPWR VPWR _31646_/A sky130_fd_sc_hd__mux2_1
X_19367_ _20211_/A VGND VGND VPWR VPWR _19367_/X sky130_fd_sc_hd__clkbuf_8
X_16579_ _33180_/Q _32540_/Q _35932_/Q _35868_/Q _16368_/X _16369_/X VGND VGND VPWR
+ VPWR _16579_/X sky130_fd_sc_hd__mux4_1
X_18318_ _20062_/A VGND VGND VPWR VPWR _20013_/A sky130_fd_sc_hd__buf_4
X_34364_ _35580_/CLK _34364_/D VGND VGND VPWR VPWR _34364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19298_ _19294_/X _19295_/X _19296_/X _19297_/X VGND VGND VPWR VPWR _19298_/X sky130_fd_sc_hd__a22o_1
X_31576_ _35996_/Q input6/X _31586_/S VGND VGND VPWR VPWR _31577_/A sky130_fd_sc_hd__mux2_1
X_36103_ _36103_/CLK _36103_/D VGND VGND VPWR VPWR _36103_/Q sky130_fd_sc_hd__dfxtp_1
X_33315_ _36055_/CLK _33315_/D VGND VGND VPWR VPWR _33315_/Q sky130_fd_sc_hd__dfxtp_1
X_18249_ _34061_/Q _33997_/Q _33933_/Q _32269_/Q _16058_/X _16060_/X VGND VGND VPWR
+ VPWR _18249_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30527_ _23234_/X _35499_/Q _30527_/S VGND VGND VPWR VPWR _30528_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34295_ _34295_/CLK _34295_/D VGND VGND VPWR VPWR _34295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36034_ _36034_/CLK _36034_/D VGND VGND VPWR VPWR _36034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21260_ _21256_/X _21259_/X _21055_/X VGND VGND VPWR VPWR _21261_/D sky130_fd_sc_hd__o21ba_1
X_33246_ _36127_/CLK _33246_/D VGND VGND VPWR VPWR _33246_/Q sky130_fd_sc_hd__dfxtp_1
X_30458_ _30458_/A VGND VGND VPWR VPWR _35466_/D sky130_fd_sc_hd__clkbuf_1
X_20211_ _20211_/A VGND VGND VPWR VPWR _20211_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_102_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_360_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _34032_/CLK sky130_fd_sc_hd__clkbuf_16
X_33177_ _35929_/CLK _33177_/D VGND VGND VPWR VPWR _33177_/Q sky130_fd_sc_hd__dfxtp_1
X_21191_ _21191_/A _21191_/B _21191_/C _21191_/D VGND VGND VPWR VPWR _21192_/A sky130_fd_sc_hd__or4_2
XFILLER_104_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30389_ _30389_/A VGND VGND VPWR VPWR _35433_/D sky130_fd_sc_hd__clkbuf_1
X_20142_ _20142_/A VGND VGND VPWR VPWR _20142_/X sky130_fd_sc_hd__buf_4
X_32128_ _35814_/CLK _32128_/D VGND VGND VPWR VPWR _32128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20073_ _20073_/A VGND VGND VPWR VPWR _20073_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_112_CLK clkbuf_6_20__f_CLK/X VGND VGND VPWR VPWR _35282_/CLK sky130_fd_sc_hd__clkbuf_16
X_32059_ _36028_/CLK _32059_/D VGND VGND VPWR VPWR _32059_/Q sky130_fd_sc_hd__dfxtp_1
X_24950_ _23019_/X _32955_/Q _24958_/S VGND VGND VPWR VPWR _24951_/A sky130_fd_sc_hd__mux2_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23901_ _23970_/S VGND VGND VPWR VPWR _23920_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_245_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24881_ _22917_/X _32922_/Q _24895_/S VGND VGND VPWR VPWR _24882_/A sky130_fd_sc_hd__mux2_1
XTAP_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26620_ _26620_/A VGND VGND VPWR VPWR _33710_/D sky130_fd_sc_hd__clkbuf_1
X_23832_ _23071_/X _32460_/Q _23834_/S VGND VGND VPWR VPWR _23833_/A sky130_fd_sc_hd__mux2_1
XTAP_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35818_ _35818_/CLK _35818_/D VGND VGND VPWR VPWR _35818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_407 _36211_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_14_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_14_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_26551_ _26683_/S VGND VGND VPWR VPWR _26570_/S sky130_fd_sc_hd__clkbuf_8
X_23763_ _22969_/X _32427_/Q _23763_/S VGND VGND VPWR VPWR _23764_/A sky130_fd_sc_hd__mux2_1
XANTENNA_418 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20975_ _20674_/X _20973_/X _20974_/X _20684_/X VGND VGND VPWR VPWR _20975_/X sky130_fd_sc_hd__a22o_1
X_35749_ _35749_/CLK _35749_/D VGND VGND VPWR VPWR _35749_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_429 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25502_ _25502_/A VGND VGND VPWR VPWR _33183_/D sky130_fd_sc_hd__clkbuf_1
X_22714_ _20597_/X _22712_/X _22713_/X _20603_/X VGND VGND VPWR VPWR _22714_/X sky130_fd_sc_hd__a22o_1
X_29270_ _29270_/A VGND VGND VPWR VPWR _34903_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23694_ _32396_/Q _23342_/X _23696_/S VGND VGND VPWR VPWR _23695_/A sky130_fd_sc_hd__mux2_1
X_26482_ _26482_/A VGND VGND VPWR VPWR _33645_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28221_ _28221_/A VGND VGND VPWR VPWR _34437_/D sky130_fd_sc_hd__clkbuf_1
X_22645_ _32518_/Q _32390_/Q _32070_/Q _36038_/Q _22582_/X _22370_/X VGND VGND VPWR
+ VPWR _22645_/X sky130_fd_sc_hd__mux4_1
X_25433_ _25433_/A VGND VGND VPWR VPWR _33152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_179_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _36041_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_29_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_29_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_28152_ _28152_/A VGND VGND VPWR VPWR _34404_/D sky130_fd_sc_hd__clkbuf_1
X_25364_ _25047_/X _33120_/Q _25366_/S VGND VGND VPWR VPWR _25365_/A sky130_fd_sc_hd__mux2_1
X_22576_ _22508_/X _22574_/X _22575_/X _22511_/X VGND VGND VPWR VPWR _22576_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27103_ _27103_/A VGND VGND VPWR VPWR _33908_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21527_ _21522_/X _21526_/X _21383_/X _21384_/X VGND VGND VPWR VPWR _21544_/B sky130_fd_sc_hd__o211a_1
X_24315_ _32676_/Q _24314_/X _24336_/S VGND VGND VPWR VPWR _24316_/A sky130_fd_sc_hd__mux2_1
X_28083_ _26990_/X _34372_/Q _28093_/S VGND VGND VPWR VPWR _28084_/A sky130_fd_sc_hd__mux2_1
X_25295_ _25322_/S VGND VGND VPWR VPWR _25314_/S sky130_fd_sc_hd__buf_6
XFILLER_166_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27034_ _27034_/A VGND VGND VPWR VPWR _33875_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24246_ _24441_/S VGND VGND VPWR VPWR _24274_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_182_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21458_ _32484_/Q _32356_/Q _32036_/Q _36004_/Q _21170_/X _21311_/X VGND VGND VPWR
+ VPWR _21458_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20409_ _35848_/Q _32228_/Q _35720_/Q _35656_/Q _18289_/X _18291_/X VGND VGND VPWR
+ VPWR _20409_/X sky130_fd_sc_hd__mux4_1
XFILLER_134_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24177_ _24177_/A VGND VGND VPWR VPWR _32621_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21389_ _35746_/Q _35106_/Q _34466_/Q _33826_/Q _21387_/X _21388_/X VGND VGND VPWR
+ VPWR _21389_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_351_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _34228_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_150_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23128_ _32155_/Q _23127_/X _23146_/S VGND VGND VPWR VPWR _23129_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28985_ _28985_/A VGND VGND VPWR VPWR _34799_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23059_ input54/X VGND VGND VPWR VPWR _23059_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_103_CLK clkbuf_leaf_80_CLK/A VGND VGND VPWR VPWR _35730_/CLK sky130_fd_sc_hd__clkbuf_16
X_27936_ _27936_/A VGND VGND VPWR VPWR _34302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput98 _31967_/Q VGND VGND VPWR VPWR D1[17] sky130_fd_sc_hd__buf_2
XTAP_6066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27867_ _27867_/A VGND VGND VPWR VPWR _34269_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ _17548_/X _17618_/X _17619_/X _17553_/X VGND VGND VPWR VPWR _17620_/X sky130_fd_sc_hd__a22o_1
X_29606_ _29606_/A VGND VGND VPWR VPWR _35062_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26818_ _26818_/A VGND VGND VPWR VPWR _33804_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27798_ _34237_/Q _24391_/X _27802_/S VGND VGND VPWR VPWR _27799_/A sky130_fd_sc_hd__mux2_1
XTAP_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29537_ _35030_/Q _29076_/X _29539_/S VGND VGND VPWR VPWR _29538_/A sky130_fd_sc_hd__mux2_1
XTAP_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _33784_/Q _33720_/Q _33656_/Q _33592_/Q _17549_/X _17550_/X VGND VGND VPWR
+ VPWR _17551_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26749_ _26749_/A VGND VGND VPWR VPWR _33771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_930 _29247_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _32730_/Q _32666_/Q _32602_/Q _36058_/Q _16213_/X _16350_/X VGND VGND VPWR
+ VPWR _16502_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_941 _29382_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_952 _29652_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29468_ _29468_/A VGND VGND VPWR VPWR _34997_/D sky130_fd_sc_hd__clkbuf_1
X_17482_ _17475_/X _17480_/X _17481_/X VGND VGND VPWR VPWR _17516_/A sky130_fd_sc_hd__o21ba_1
XANTENNA_963 _30057_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_974 _31948_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1006 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19221_ _33254_/Q _36134_/Q _33126_/Q _33062_/Q _19005_/X _19006_/X VGND VGND VPWR
+ VPWR _19221_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_985 _17795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28419_ _26888_/X _34531_/Q _28435_/S VGND VGND VPWR VPWR _28420_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_956 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16433_ _35800_/Q _32175_/Q _35672_/Q _35608_/Q _16254_/X _16255_/X VGND VGND VPWR
+ VPWR _16433_/X sky130_fd_sc_hd__mux4_1
XANTENNA_996 _17956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29399_ _29399_/A VGND VGND VPWR VPWR _34964_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31430_ _23114_/X _35927_/Q _31430_/S VGND VGND VPWR VPWR _31431_/A sky130_fd_sc_hd__mux2_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19152_ _20211_/A VGND VGND VPWR VPWR _19152_/X sky130_fd_sc_hd__buf_4
X_16364_ _35798_/Q _32173_/Q _35670_/Q _35606_/Q _16254_/X _16255_/X VGND VGND VPWR
+ VPWR _16364_/X sky130_fd_sc_hd__mux4_1
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18103_ _33288_/Q _36168_/Q _33160_/Q _33096_/Q _16028_/X _17157_/A VGND VGND VPWR
+ VPWR _18103_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19083_ _20142_/A VGND VGND VPWR VPWR _19083_/X sky130_fd_sc_hd__clkbuf_4
X_31361_ _35894_/Q input35/X _31379_/S VGND VGND VPWR VPWR _31362_/A sky130_fd_sc_hd__mux2_1
X_16295_ _33172_/Q _32532_/Q _35924_/Q _35860_/Q _16063_/X _16065_/X VGND VGND VPWR
+ VPWR _16295_/X sky130_fd_sc_hd__mux4_1
X_33100_ _36170_/CLK _33100_/D VGND VGND VPWR VPWR _33100_/Q sky130_fd_sc_hd__dfxtp_1
X_18034_ _18034_/A VGND VGND VPWR VPWR _32005_/D sky130_fd_sc_hd__clkbuf_2
X_30312_ _30312_/A VGND VGND VPWR VPWR _35397_/D sky130_fd_sc_hd__clkbuf_1
X_34080_ _34080_/CLK _34080_/D VGND VGND VPWR VPWR _34080_/Q sky130_fd_sc_hd__dfxtp_1
X_31292_ _31292_/A VGND VGND VPWR VPWR _35861_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33031_ _34752_/CLK _33031_/D VGND VGND VPWR VPWR _33031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30243_ _30243_/A VGND VGND VPWR VPWR _35364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_342_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _34293_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_113_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30174_ _35332_/Q _29219_/X _30184_/S VGND VGND VPWR VPWR _30175_/A sky130_fd_sc_hd__mux2_1
X_19985_ _34300_/Q _34236_/Q _34172_/Q _34108_/Q _19742_/X _19743_/X VGND VGND VPWR
+ VPWR _19985_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18936_ _20129_/A VGND VGND VPWR VPWR _18936_/X sky130_fd_sc_hd__buf_4
XANTENNA_1340 _20203_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34982_ _35239_/CLK _34982_/D VGND VGND VPWR VPWR _34982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1351 _21757_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1362 _24244_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33933_ _34060_/CLK _33933_/D VGND VGND VPWR VPWR _33933_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1373 _25872_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18867_ _32732_/Q _32668_/Q _32604_/Q _36060_/Q _18866_/X _18650_/X VGND VGND VPWR
+ VPWR _18867_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1384 _31003_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1395 input87/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17818_ _35327_/Q _35263_/Q _35199_/Q _32319_/Q _17712_/X _17713_/X VGND VGND VPWR
+ VPWR _17818_/X sky130_fd_sc_hd__mux4_1
X_33864_ _35847_/CLK _33864_/D VGND VGND VPWR VPWR _33864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18798_ _34010_/Q _33946_/Q _33882_/Q _32154_/Q _18614_/X _18615_/X VGND VGND VPWR
+ VPWR _18798_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35603_ _35797_/CLK _35603_/D VGND VGND VPWR VPWR _35603_/Q sky130_fd_sc_hd__dfxtp_1
X_32815_ _33007_/CLK _32815_/D VGND VGND VPWR VPWR _32815_/Q sky130_fd_sc_hd__dfxtp_1
X_17749_ _35069_/Q _35005_/Q _34941_/Q _34877_/Q _17509_/X _17510_/X VGND VGND VPWR
+ VPWR _17749_/X sky130_fd_sc_hd__mux4_1
X_33795_ _33795_/CLK _33795_/D VGND VGND VPWR VPWR _33795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35534_ _35793_/CLK _35534_/D VGND VGND VPWR VPWR _35534_/Q sky130_fd_sc_hd__dfxtp_1
X_20760_ _33168_/Q _32528_/Q _35920_/Q _35856_/Q _20663_/X _20665_/X VGND VGND VPWR
+ VPWR _20760_/X sky130_fd_sc_hd__mux4_1
X_32746_ _36139_/CLK _32746_/D VGND VGND VPWR VPWR _32746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19419_ _19419_/A VGND VGND VPWR VPWR _32107_/D sky130_fd_sc_hd__clkbuf_1
X_35465_ _35975_/CLK _35465_/D VGND VGND VPWR VPWR _35465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20691_ _34510_/Q _32398_/Q _34382_/Q _34318_/Q _20688_/X _20690_/X VGND VGND VPWR
+ VPWR _20691_/X sky130_fd_sc_hd__mux4_1
X_32677_ _36070_/CLK _32677_/D VGND VGND VPWR VPWR _32677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22430_ _22430_/A VGND VGND VPWR VPWR _22430_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_182_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34416_ _35052_/CLK _34416_/D VGND VGND VPWR VPWR _34416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31628_ _36021_/Q input33/X _31628_/S VGND VGND VPWR VPWR _31629_/A sky130_fd_sc_hd__mux2_1
X_35396_ _35715_/CLK _35396_/D VGND VGND VPWR VPWR _35396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22361_ _22361_/A VGND VGND VPWR VPWR _22361_/X sky130_fd_sc_hd__clkbuf_4
X_34347_ _35944_/CLK _34347_/D VGND VGND VPWR VPWR _34347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31559_ _35988_/Q input61/X _31565_/S VGND VGND VPWR VPWR _31560_/A sky130_fd_sc_hd__mux2_1
X_24100_ _23065_/X _32586_/Q _24106_/S VGND VGND VPWR VPWR _24101_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21312_ _32480_/Q _32352_/Q _32032_/Q _36000_/Q _21170_/X _21311_/X VGND VGND VPWR
+ VPWR _21312_/X sky130_fd_sc_hd__mux4_1
X_25080_ _25080_/A VGND VGND VPWR VPWR _33002_/D sky130_fd_sc_hd__clkbuf_1
X_22292_ _33276_/Q _36156_/Q _33148_/Q _33084_/Q _22011_/X _22012_/X VGND VGND VPWR
+ VPWR _22292_/X sky130_fd_sc_hd__mux4_1
X_34278_ _34278_/CLK _34278_/D VGND VGND VPWR VPWR _34278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1044 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36017_ _36076_/CLK _36017_/D VGND VGND VPWR VPWR _36017_/Q sky130_fd_sc_hd__dfxtp_1
X_24031_ _22963_/X _32553_/Q _24035_/S VGND VGND VPWR VPWR _24032_/A sky130_fd_sc_hd__mux2_1
X_33229_ _35917_/CLK _33229_/D VGND VGND VPWR VPWR _33229_/Q sky130_fd_sc_hd__dfxtp_1
X_21243_ _35742_/Q _35102_/Q _34462_/Q _33822_/Q _21034_/X _21035_/X VGND VGND VPWR
+ VPWR _21243_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_333_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _36025_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21174_ _21169_/X _21173_/X _21030_/X _21031_/X VGND VGND VPWR VPWR _21191_/B sky130_fd_sc_hd__o211a_1
XFILLER_172_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20125_ _20125_/A VGND VGND VPWR VPWR _32127_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_63_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28770_ _27008_/X _34698_/Q _28776_/S VGND VGND VPWR VPWR _28771_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25982_ _25982_/A VGND VGND VPWR VPWR _33408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27721_ _34200_/Q _24276_/X _27739_/S VGND VGND VPWR VPWR _27722_/A sky130_fd_sc_hd__mux2_1
X_20056_ _19848_/X _20054_/X _20055_/X _19853_/X VGND VGND VPWR VPWR _20056_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24933_ _22994_/X _32947_/Q _24937_/S VGND VGND VPWR VPWR _24934_/A sky130_fd_sc_hd__mux2_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27652_ _27652_/A VGND VGND VPWR VPWR _34167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24864_ _22892_/X _32914_/Q _24874_/S VGND VGND VPWR VPWR _24865_/A sky130_fd_sc_hd__mux2_1
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26603_ _26603_/A VGND VGND VPWR VPWR _33702_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23815_ _23815_/A VGND VGND VPWR VPWR _32451_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_204 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27583_ _34135_/Q _24273_/X _27583_/S VGND VGND VPWR VPWR _27584_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24795_ _24795_/A VGND VGND VPWR VPWR _32881_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_215 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_226 _32136_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29322_ _23250_/X _34928_/Q _29332_/S VGND VGND VPWR VPWR _29323_/A sky130_fd_sc_hd__mux2_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26534_ _26534_/A VGND VGND VPWR VPWR _33670_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_248 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_259 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20958_ _22370_/A VGND VGND VPWR VPWR _20958_/X sky130_fd_sc_hd__buf_4
X_23746_ _23746_/A VGND VGND VPWR VPWR _32418_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29253_ _23090_/X _34895_/Q _29269_/S VGND VGND VPWR VPWR _29254_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26465_ _26465_/A VGND VGND VPWR VPWR _33637_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23677_ _23677_/A VGND VGND VPWR VPWR _32387_/D sky130_fd_sc_hd__clkbuf_1
X_20889_ _35796_/Q _32170_/Q _35668_/Q _35604_/Q _20854_/X _20855_/X VGND VGND VPWR
+ VPWR _20889_/X sky130_fd_sc_hd__mux4_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28204_ _28204_/A VGND VGND VPWR VPWR _34429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25416_ _25416_/A VGND VGND VPWR VPWR _33144_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22628_ _22455_/X _22626_/X _22627_/X _22458_/X VGND VGND VPWR VPWR _22628_/X sky130_fd_sc_hd__a22o_1
XFILLER_224_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29184_ _29184_/A VGND VGND VPWR VPWR _34872_/D sky130_fd_sc_hd__clkbuf_1
X_26396_ _25162_/X _33605_/Q _26404_/S VGND VGND VPWR VPWR _26397_/A sky130_fd_sc_hd__mux2_1
X_28135_ _28135_/A VGND VGND VPWR VPWR _34396_/D sky130_fd_sc_hd__clkbuf_1
X_22559_ _33219_/Q _32579_/Q _35971_/Q _35907_/Q _22380_/X _22381_/X VGND VGND VPWR
+ VPWR _22559_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25347_ _25458_/S VGND VGND VPWR VPWR _25366_/S sky130_fd_sc_hd__buf_4
XFILLER_220_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16080_ _17762_/A VGND VGND VPWR VPWR _17007_/A sky130_fd_sc_hd__buf_12
XFILLER_154_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28066_ _26965_/X _34364_/Q _28072_/S VGND VGND VPWR VPWR _28067_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25278_ _25278_/A VGND VGND VPWR VPWR _33079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27017_ input60/X VGND VGND VPWR VPWR _27017_/X sky130_fd_sc_hd__clkbuf_4
X_24229_ _24229_/A VGND VGND VPWR VPWR _32646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_324_CLK clkbuf_6_38__f_CLK/X VGND VGND VPWR VPWR _35700_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_194_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19770_ _19766_/X _19769_/X _19461_/X VGND VGND VPWR VPWR _19771_/D sky130_fd_sc_hd__o21ba_1
XFILLER_231_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28968_ _28968_/A VGND VGND VPWR VPWR _34791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16982_ _34024_/Q _33960_/Q _33896_/Q _32215_/Q _16667_/X _16668_/X VGND VGND VPWR
+ VPWR _16982_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18721_ _18443_/X _18719_/X _18720_/X _18446_/X VGND VGND VPWR VPWR _18721_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27919_ _34294_/Q _24369_/X _27937_/S VGND VGND VPWR VPWR _27920_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28899_ _26999_/X _34759_/Q _28903_/S VGND VGND VPWR VPWR _28900_/A sky130_fd_sc_hd__mux2_1
XTAP_5151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18652_ _20202_/A VGND VGND VPWR VPWR _18652_/X sky130_fd_sc_hd__buf_4
XFILLER_7_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30930_ _35690_/Q _29138_/X _30932_/S VGND VGND VPWR VPWR _30931_/A sky130_fd_sc_hd__mux2_1
XTAP_5195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17603_ _17956_/A VGND VGND VPWR VPWR _17603_/X sky130_fd_sc_hd__buf_4
XTAP_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30861_ _30861_/A VGND VGND VPWR VPWR _35657_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18583_ _20129_/A VGND VGND VPWR VPWR _18583_/X sky130_fd_sc_hd__buf_4
XFILLER_131_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32600_ _32666_/CLK _32600_/D VGND VGND VPWR VPWR _32600_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17534_ _17347_/X _17532_/X _17533_/X _17350_/X VGND VGND VPWR VPWR _17534_/X sky130_fd_sc_hd__a22o_1
XTAP_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33580_ _34283_/CLK _33580_/D VGND VGND VPWR VPWR _33580_/Q sky130_fd_sc_hd__dfxtp_1
X_30792_ _30792_/A VGND VGND VPWR VPWR _35624_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_760 _22500_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_771 _22538_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32531_ _36114_/CLK _32531_/D VGND VGND VPWR VPWR _32531_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_782 _22604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17465_ _35317_/Q _35253_/Q _35189_/Q _32309_/Q _17359_/X _17360_/X VGND VGND VPWR
+ VPWR _17465_/X sky130_fd_sc_hd__mux4_1
XANTENNA_793 _22694_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19204_ _35301_/Q _35237_/Q _35173_/Q _32293_/Q _18953_/X _18954_/X VGND VGND VPWR
+ VPWR _19204_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16416_ _16136_/X _16414_/X _16415_/X _16141_/X VGND VGND VPWR VPWR _16416_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_786 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35250_ _35250_/CLK _35250_/D VGND VGND VPWR VPWR _35250_/Q sky130_fd_sc_hd__dfxtp_1
X_32462_ _35982_/CLK _32462_/D VGND VGND VPWR VPWR _32462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17396_ _35059_/Q _34995_/Q _34931_/Q _34867_/Q _17156_/X _17157_/X VGND VGND VPWR
+ VPWR _17396_/X sky130_fd_sc_hd__mux4_1
X_34201_ _35671_/CLK _34201_/D VGND VGND VPWR VPWR _34201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31413_ _31413_/A VGND VGND VPWR VPWR _35918_/D sky130_fd_sc_hd__clkbuf_1
X_19135_ _19096_/X _19133_/X _19134_/X _19099_/X VGND VGND VPWR VPWR _19135_/X sky130_fd_sc_hd__a22o_1
X_16347_ _16143_/X _16345_/X _16346_/X _16146_/X VGND VGND VPWR VPWR _16347_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35181_ _35307_/CLK _35181_/D VGND VGND VPWR VPWR _35181_/Q sky130_fd_sc_hd__dfxtp_1
X_32393_ _36107_/CLK _32393_/D VGND VGND VPWR VPWR _32393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34132_ _34260_/CLK _34132_/D VGND VGND VPWR VPWR _34132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31344_ _35886_/Q input26/X _31358_/S VGND VGND VPWR VPWR _31345_/A sky130_fd_sc_hd__mux2_1
X_19066_ _19066_/A VGND VGND VPWR VPWR _32097_/D sky130_fd_sc_hd__clkbuf_1
X_16278_ _16274_/X _16277_/X _16011_/X VGND VGND VPWR VPWR _16308_/A sky130_fd_sc_hd__o21ba_2
XFILLER_146_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18017_ _17769_/X _18015_/X _18016_/X _17773_/X VGND VGND VPWR VPWR _18017_/X sky130_fd_sc_hd__a22o_1
X_34063_ _35021_/CLK _34063_/D VGND VGND VPWR VPWR _34063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31275_ _31275_/A _31275_/B VGND VGND VPWR VPWR _31408_/S sky130_fd_sc_hd__nor2_8
Xclkbuf_leaf_315_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _35768_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_126_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33014_ _36087_/CLK _33014_/D VGND VGND VPWR VPWR _33014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30226_ _30226_/A VGND VGND VPWR VPWR _35356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30157_ _35324_/Q _29194_/X _30163_/S VGND VGND VPWR VPWR _30158_/A sky130_fd_sc_hd__mux2_1
X_19968_ _35835_/Q _32213_/Q _35707_/Q _35643_/Q _19966_/X _19967_/X VGND VGND VPWR
+ VPWR _19968_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18919_ _34525_/Q _32413_/Q _34397_/Q _34333_/Q _18819_/X _18820_/X VGND VGND VPWR
+ VPWR _18919_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34965_ _34967_/CLK _34965_/D VGND VGND VPWR VPWR _34965_/Q sky130_fd_sc_hd__dfxtp_1
X_30088_ _35291_/Q _29092_/X _30100_/S VGND VGND VPWR VPWR _30089_/A sky130_fd_sc_hd__mux2_1
XANTENNA_1170 _22447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19899_ _19895_/X _19898_/X _19789_/X _19790_/X VGND VGND VPWR VPWR _19916_/B sky130_fd_sc_hd__o211a_1
XFILLER_80_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1181 _21589_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1192 _22889_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33916_ _34171_/CLK _33916_/D VGND VGND VPWR VPWR _33916_/Q sky130_fd_sc_hd__dfxtp_1
X_21930_ _21930_/A VGND VGND VPWR VPWR _36209_/D sky130_fd_sc_hd__buf_6
X_34896_ _35026_/CLK _34896_/D VGND VGND VPWR VPWR _34896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21861_ _21754_/X _21859_/X _21860_/X _21759_/X VGND VGND VPWR VPWR _21861_/X sky130_fd_sc_hd__a22o_1
XFILLER_209_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33847_ _34809_/CLK _33847_/D VGND VGND VPWR VPWR _33847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20812_ _20808_/X _20811_/X _20611_/X VGND VGND VPWR VPWR _20838_/A sky130_fd_sc_hd__o21ba_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23600_ _32351_/Q _23139_/X _23604_/S VGND VGND VPWR VPWR _23601_/A sky130_fd_sc_hd__mux2_1
X_24580_ input86/X _30329_/B input88/X VGND VGND VPWR VPWR _24581_/A sky130_fd_sc_hd__and3b_1
X_21792_ _21788_/X _21791_/X _21761_/X VGND VGND VPWR VPWR _21793_/D sky130_fd_sc_hd__o21ba_1
X_33778_ _34288_/CLK _33778_/D VGND VGND VPWR VPWR _33778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23531_ _23531_/A VGND VGND VPWR VPWR _32319_/D sky130_fd_sc_hd__clkbuf_1
X_35517_ _35517_/CLK _35517_/D VGND VGND VPWR VPWR _35517_/Q sky130_fd_sc_hd__dfxtp_1
X_20743_ _22460_/A VGND VGND VPWR VPWR _20743_/X sky130_fd_sc_hd__buf_4
X_32729_ _36119_/CLK _32729_/D VGND VGND VPWR VPWR _32729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26250_ _26277_/S VGND VGND VPWR VPWR _26269_/S sky130_fd_sc_hd__buf_4
XFILLER_168_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23462_ _23462_/A VGND VGND VPWR VPWR _32286_/D sky130_fd_sc_hd__clkbuf_1
X_20674_ _21749_/A VGND VGND VPWR VPWR _20674_/X sky130_fd_sc_hd__buf_4
X_35448_ _35638_/CLK _35448_/D VGND VGND VPWR VPWR _35448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22413_ _35583_/Q _35519_/Q _35455_/Q _35391_/Q _22203_/X _22204_/X VGND VGND VPWR
+ VPWR _22413_/X sky130_fd_sc_hd__mux4_1
X_25201_ _25007_/X _33043_/Q _25209_/S VGND VGND VPWR VPWR _25202_/A sky130_fd_sc_hd__mux2_1
X_23393_ _23393_/A VGND VGND VPWR VPWR _32255_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26181_ _25044_/X _33503_/Q _26185_/S VGND VGND VPWR VPWR _26182_/A sky130_fd_sc_hd__mux2_1
X_35379_ _35827_/CLK _35379_/D VGND VGND VPWR VPWR _35379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22344_ _22340_/X _22343_/X _22100_/X VGND VGND VPWR VPWR _22352_/C sky130_fd_sc_hd__o21ba_1
XFILLER_148_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25132_ _25131_/X _33019_/Q _25144_/S VGND VGND VPWR VPWR _25133_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29940_ _35221_/Q _29073_/X _29944_/S VGND VGND VPWR VPWR _29941_/A sky130_fd_sc_hd__mux2_1
X_25063_ input16/X VGND VGND VPWR VPWR _25063_/X sky130_fd_sc_hd__buf_2
X_22275_ _34811_/Q _34747_/Q _34683_/Q _34619_/Q _22241_/X _22242_/X VGND VGND VPWR
+ VPWR _22275_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_306_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _35579_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24014_ _22938_/X _32545_/Q _24014_/S VGND VGND VPWR VPWR _24015_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21226_ _34270_/Q _34206_/Q _34142_/Q _34078_/Q _20983_/X _20984_/X VGND VGND VPWR
+ VPWR _21226_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29871_ _29871_/A VGND VGND VPWR VPWR _35188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28822_ _26884_/X _34722_/Q _28840_/S VGND VGND VPWR VPWR _28823_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21157_ _21157_/A _21157_/B _21157_/C _21157_/D VGND VGND VPWR VPWR _21158_/A sky130_fd_sc_hd__or4_2
X_20108_ _20069_/X _20106_/X _20107_/X _20073_/X VGND VGND VPWR VPWR _20108_/X sky130_fd_sc_hd__a22o_1
X_28753_ _28753_/A VGND VGND VPWR VPWR _34689_/D sky130_fd_sc_hd__clkbuf_1
X_21088_ _21088_/A VGND VGND VPWR VPWR _36185_/D sky130_fd_sc_hd__clkbuf_1
X_25965_ _25965_/A VGND VGND VPWR VPWR _33400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27704_ _34192_/Q _24252_/X _27718_/S VGND VGND VPWR VPWR _27705_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20039_ _35773_/Q _35133_/Q _34493_/Q _33853_/Q _19793_/X _19794_/X VGND VGND VPWR
+ VPWR _20039_/X sky130_fd_sc_hd__mux4_1
X_24916_ _22969_/X _32939_/Q _24916_/S VGND VGND VPWR VPWR _24917_/A sky130_fd_sc_hd__mux2_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28684_ _26881_/X _34657_/Q _28684_/S VGND VGND VPWR VPWR _28685_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25896_ _26007_/S VGND VGND VPWR VPWR _25915_/S sky130_fd_sc_hd__buf_4
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27635_ _27635_/A VGND VGND VPWR VPWR _34159_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24847_ _24847_/A VGND VGND VPWR VPWR _32906_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27566_ _27566_/A VGND VGND VPWR VPWR _34126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24778_ _24778_/A VGND VGND VPWR VPWR _32873_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29305_ _23223_/X _34920_/Q _29311_/S VGND VGND VPWR VPWR _29306_/A sky130_fd_sc_hd__mux2_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26517_ _26517_/A VGND VGND VPWR VPWR _33662_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23729_ _23729_/A VGND VGND VPWR VPWR _32410_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27497_ _26925_/X _34095_/Q _27509_/S VGND VGND VPWR VPWR _27498_/A sky130_fd_sc_hd__mux2_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29236_ _29236_/A VGND VGND VPWR VPWR _34889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _17956_/A VGND VGND VPWR VPWR _17250_/X sky130_fd_sc_hd__buf_6
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26448_ _26448_/A VGND VGND VPWR VPWR _33629_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16201_ _35025_/Q _34961_/Q _34897_/Q _34833_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _16201_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17181_ _16994_/X _17179_/X _17180_/X _16997_/X VGND VGND VPWR VPWR _17181_/X sky130_fd_sc_hd__a22o_1
X_29167_ _34867_/Q _29166_/X _29173_/S VGND VGND VPWR VPWR _29168_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26379_ _25137_/X _33597_/Q _26383_/S VGND VGND VPWR VPWR _26380_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16132_ _16087_/X _16130_/X _16131_/X _16097_/X VGND VGND VPWR VPWR _16132_/X sky130_fd_sc_hd__a22o_1
X_28118_ _28118_/A VGND VGND VPWR VPWR _34388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29098_ input7/X VGND VGND VPWR VPWR _29098_/X sky130_fd_sc_hd__buf_4
XFILLER_196_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16063_ _17931_/A VGND VGND VPWR VPWR _16063_/X sky130_fd_sc_hd__buf_6
X_28049_ _26940_/X _34356_/Q _28051_/S VGND VGND VPWR VPWR _28050_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31060_ _31060_/A VGND VGND VPWR VPWR _35751_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_1192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30011_ _30011_/A VGND VGND VPWR VPWR _35254_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19822_ _34039_/Q _33975_/Q _33911_/Q _32247_/Q _19673_/X _19674_/X VGND VGND VPWR
+ VPWR _19822_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16965_ _35559_/Q _35495_/Q _35431_/Q _35367_/Q _16897_/X _16898_/X VGND VGND VPWR
+ VPWR _16965_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19753_ _32501_/Q _32373_/Q _32053_/Q _36021_/Q _19576_/X _19717_/X VGND VGND VPWR
+ VPWR _19753_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18704_ _18700_/X _18703_/X _18371_/X VGND VGND VPWR VPWR _18712_/C sky130_fd_sc_hd__o21ba_1
X_34750_ _36031_/CLK _34750_/D VGND VGND VPWR VPWR _34750_/Q sky130_fd_sc_hd__dfxtp_1
X_31962_ _35166_/CLK _31962_/D VGND VGND VPWR VPWR _31962_/Q sky130_fd_sc_hd__dfxtp_1
X_19684_ _19680_/X _19683_/X _19436_/X _19437_/X VGND VGND VPWR VPWR _19699_/B sky130_fd_sc_hd__o211a_1
X_16896_ _16641_/X _16894_/X _16895_/X _16644_/X VGND VGND VPWR VPWR _16896_/X sky130_fd_sc_hd__a22o_1
XFILLER_231_1097 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18635_ _18374_/X _18633_/X _18634_/X _18384_/X VGND VGND VPWR VPWR _18635_/X sky130_fd_sc_hd__a22o_1
X_33701_ _33702_/CLK _33701_/D VGND VGND VPWR VPWR _33701_/Q sky130_fd_sc_hd__dfxtp_1
X_30913_ _31003_/S VGND VGND VPWR VPWR _30932_/S sky130_fd_sc_hd__buf_4
XTAP_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34681_ _34745_/CLK _34681_/D VGND VGND VPWR VPWR _34681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31893_ _31893_/A VGND VGND VPWR VPWR _36146_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33632_ _34080_/CLK _33632_/D VGND VGND VPWR VPWR _33632_/Q sky130_fd_sc_hd__dfxtp_1
X_30844_ _23307_/X _35649_/Q _30860_/S VGND VGND VPWR VPWR _30845_/A sky130_fd_sc_hd__mux2_1
X_18566_ _34515_/Q _32403_/Q _34387_/Q _34323_/Q _18466_/X _18467_/X VGND VGND VPWR
+ VPWR _18566_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17517_ _17517_/A VGND VGND VPWR VPWR _31990_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_220_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33563_ _34267_/CLK _33563_/D VGND VGND VPWR VPWR _33563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18497_ _34769_/Q _34705_/Q _34641_/Q _34577_/Q _18375_/X _18376_/X VGND VGND VPWR
+ VPWR _18497_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30775_ _30775_/A VGND VGND VPWR VPWR _35616_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_590 _19457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32514_ _32962_/CLK _32514_/D VGND VGND VPWR VPWR _32514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35302_ _35302_/CLK _35302_/D VGND VGND VPWR VPWR _35302_/Q sky130_fd_sc_hd__dfxtp_1
X_17448_ _17202_/X _17446_/X _17447_/X _17205_/X VGND VGND VPWR VPWR _17448_/X sky130_fd_sc_hd__a22o_1
XFILLER_221_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33494_ _34001_/CLK _33494_/D VGND VGND VPWR VPWR _33494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32445_ _35581_/CLK _32445_/D VGND VGND VPWR VPWR _32445_/Q sky130_fd_sc_hd__dfxtp_1
X_35233_ _35296_/CLK _35233_/D VGND VGND VPWR VPWR _35233_/Q sky130_fd_sc_hd__dfxtp_1
X_17379_ _33267_/Q _36147_/Q _33139_/Q _33075_/Q _17058_/X _17059_/X VGND VGND VPWR
+ VPWR _17379_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_92_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _36185_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19118_ _19114_/X _19117_/X _19075_/X VGND VGND VPWR VPWR _19140_/A sky130_fd_sc_hd__o21ba_1
X_35164_ _35164_/CLK _35164_/D VGND VGND VPWR VPWR _35164_/Q sky130_fd_sc_hd__dfxtp_1
X_20390_ _35079_/Q _35015_/Q _34951_/Q _34887_/Q _20162_/X _20163_/X VGND VGND VPWR
+ VPWR _20390_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32376_ _36025_/CLK _32376_/D VGND VGND VPWR VPWR _32376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34115_ _34243_/CLK _34115_/D VGND VGND VPWR VPWR _34115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31327_ _35878_/Q input17/X _31337_/S VGND VGND VPWR VPWR _31328_/A sky130_fd_sc_hd__mux2_1
X_19049_ _19010_/X _19047_/X _19048_/X _19014_/X VGND VGND VPWR VPWR _19049_/X sky130_fd_sc_hd__a22o_1
X_35095_ _35733_/CLK _35095_/D VGND VGND VPWR VPWR _35095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput200 _36225_/Q VGND VGND VPWR VPWR D2[51] sky130_fd_sc_hd__buf_2
XFILLER_160_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput211 _36235_/Q VGND VGND VPWR VPWR D2[61] sky130_fd_sc_hd__buf_2
Xoutput222 _32091_/Q VGND VGND VPWR VPWR D3[13] sky130_fd_sc_hd__buf_2
X_34046_ _34046_/CLK _34046_/D VGND VGND VPWR VPWR _34046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput233 _32101_/Q VGND VGND VPWR VPWR D3[23] sky130_fd_sc_hd__buf_2
X_22060_ _35573_/Q _35509_/Q _35445_/Q _35381_/Q _21850_/X _21851_/X VGND VGND VPWR
+ VPWR _22060_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31258_ _31258_/A VGND VGND VPWR VPWR _35845_/D sky130_fd_sc_hd__clkbuf_1
Xoutput244 _32111_/Q VGND VGND VPWR VPWR D3[33] sky130_fd_sc_hd__buf_2
XFILLER_138_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput255 _32121_/Q VGND VGND VPWR VPWR D3[43] sky130_fd_sc_hd__buf_2
XFILLER_160_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21011_ _21007_/X _21010_/X _20700_/X VGND VGND VPWR VPWR _21012_/D sky130_fd_sc_hd__o21ba_1
XFILLER_138_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput266 _32131_/Q VGND VGND VPWR VPWR D3[53] sky130_fd_sc_hd__buf_2
XFILLER_99_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30209_ _30209_/A VGND VGND VPWR VPWR _35348_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput277 _32141_/Q VGND VGND VPWR VPWR D3[63] sky130_fd_sc_hd__buf_2
XTAP_5909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31189_ _31189_/A VGND VGND VPWR VPWR _35812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35997_ _36129_/CLK _35997_/D VGND VGND VPWR VPWR _35997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25750_ _25750_/A VGND VGND VPWR VPWR _33298_/D sky130_fd_sc_hd__clkbuf_1
X_34948_ _35779_/CLK _34948_/D VGND VGND VPWR VPWR _34948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22962_ _22962_/A VGND VGND VPWR VPWR _32040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24701_ _23053_/X _32838_/Q _24707_/S VGND VGND VPWR VPWR _24702_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21913_ _22395_/A VGND VGND VPWR VPWR _21913_/X sky130_fd_sc_hd__buf_6
XFILLER_28_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25681_ _33267_/Q _24360_/X _25685_/S VGND VGND VPWR VPWR _25682_/A sky130_fd_sc_hd__mux2_1
X_34879_ _35982_/CLK _34879_/D VGND VGND VPWR VPWR _34879_/Q sky130_fd_sc_hd__dfxtp_1
X_22893_ _22892_/X _32018_/Q _22908_/S VGND VGND VPWR VPWR _22894_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27420_ _34059_/Q _24434_/X _27424_/S VGND VGND VPWR VPWR _27421_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24632_ _22951_/X _32805_/Q _24644_/S VGND VGND VPWR VPWR _24633_/A sky130_fd_sc_hd__mux2_1
X_21844_ _33007_/Q _32943_/Q _32879_/Q _32815_/Q _21589_/X _21590_/X VGND VGND VPWR
+ VPWR _21844_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27351_ _34026_/Q _24332_/X _27353_/S VGND VGND VPWR VPWR _27352_/A sky130_fd_sc_hd__mux2_1
X_24563_ _23053_/X _32774_/Q _24569_/S VGND VGND VPWR VPWR _24564_/A sky130_fd_sc_hd__mux2_1
X_21775_ _32493_/Q _32365_/Q _32045_/Q _36013_/Q _21523_/X _21664_/X VGND VGND VPWR
+ VPWR _21775_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26302_ _25022_/X _33560_/Q _26320_/S VGND VGND VPWR VPWR _26303_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_786 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20726_ _20722_/X _20725_/X _20671_/X VGND VGND VPWR VPWR _20734_/C sky130_fd_sc_hd__o21ba_1
X_23514_ _23007_/X _32311_/Q _23530_/S VGND VGND VPWR VPWR _23515_/A sky130_fd_sc_hd__mux2_1
X_27282_ _27282_/A VGND VGND VPWR VPWR _33993_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24494_ _22951_/X _32741_/Q _24506_/S VGND VGND VPWR VPWR _24495_/A sky130_fd_sc_hd__mux2_1
X_29021_ _29021_/A VGND VGND VPWR VPWR _34816_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26233_ _26233_/A VGND VGND VPWR VPWR _33527_/D sky130_fd_sc_hd__clkbuf_1
X_20657_ _20657_/A VGND VGND VPWR VPWR _22446_/A sky130_fd_sc_hd__buf_12
X_23445_ _23445_/A VGND VGND VPWR VPWR _32278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_83_CLK clkbuf_leaf_87_CLK/A VGND VGND VPWR VPWR _35927_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_183_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26164_ _25019_/X _33495_/Q _26164_/S VGND VGND VPWR VPWR _26165_/A sky130_fd_sc_hd__mux2_1
X_23376_ _32247_/Q _23274_/X _23392_/S VGND VGND VPWR VPWR _23377_/A sky130_fd_sc_hd__mux2_1
X_20588_ _20657_/A VGND VGND VPWR VPWR _22395_/A sky130_fd_sc_hd__buf_12
XFILLER_164_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25115_ input35/X VGND VGND VPWR VPWR _25115_/X sky130_fd_sc_hd__buf_2
X_22327_ _22447_/A VGND VGND VPWR VPWR _22327_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_124_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26095_ _25115_/X _33462_/Q _26113_/S VGND VGND VPWR VPWR _26096_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29923_ _29923_/A VGND VGND VPWR VPWR _35213_/D sky130_fd_sc_hd__clkbuf_1
X_22258_ _22254_/X _22257_/X _22081_/X VGND VGND VPWR VPWR _22282_/A sky130_fd_sc_hd__o21ba_1
X_25046_ _25046_/A VGND VGND VPWR VPWR _32991_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21209_ _35805_/Q _32180_/Q _35677_/Q _35613_/Q _21207_/X _21208_/X VGND VGND VPWR
+ VPWR _21209_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29854_ _35180_/Q _29144_/X _29872_/S VGND VGND VPWR VPWR _29855_/A sky130_fd_sc_hd__mux2_1
X_22189_ _33529_/Q _33465_/Q _33401_/Q _33337_/Q _22076_/X _22077_/X VGND VGND VPWR
+ VPWR _22189_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28805_ _26860_/X _34714_/Q _28819_/S VGND VGND VPWR VPWR _28806_/A sky130_fd_sc_hd__mux2_1
X_29785_ _35148_/Q _29243_/X _29787_/S VGND VGND VPWR VPWR _29786_/A sky130_fd_sc_hd__mux2_1
X_26997_ _26996_/X _33862_/Q _27006_/S VGND VGND VPWR VPWR _26998_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16750_ _16746_/X _16749_/X _16430_/X _16431_/X VGND VGND VPWR VPWR _16765_/B sky130_fd_sc_hd__o211a_2
X_28736_ _28736_/A VGND VGND VPWR VPWR _34681_/D sky130_fd_sc_hd__clkbuf_1
X_25948_ _25948_/A VGND VGND VPWR VPWR _33392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16681_ _16641_/X _16679_/X _16680_/X _16644_/X VGND VGND VPWR VPWR _16681_/X sky130_fd_sc_hd__a22o_1
X_28667_ _28667_/A VGND VGND VPWR VPWR _34648_/D sky130_fd_sc_hd__clkbuf_1
X_25879_ _25879_/A VGND VGND VPWR VPWR _33359_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18420_ _35791_/Q _32165_/Q _35663_/Q _35599_/Q _18345_/X _18346_/X VGND VGND VPWR
+ VPWR _18420_/X sky130_fd_sc_hd__mux4_1
X_27618_ _27618_/A VGND VGND VPWR VPWR _34151_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28598_ _26953_/X _34616_/Q _28612_/S VGND VGND VPWR VPWR _28599_/A sky130_fd_sc_hd__mux2_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _20295_/A VGND VGND VPWR VPWR _18351_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_163_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27549_ _27002_/X _34120_/Q _27551_/S VGND VGND VPWR VPWR _27550_/A sky130_fd_sc_hd__mux2_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17302_ _33521_/Q _33457_/Q _33393_/Q _33329_/Q _17123_/X _17124_/X VGND VGND VPWR
+ VPWR _17302_/X sky130_fd_sc_hd__mux4_1
XFILLER_199_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18282_ _18359_/A VGND VGND VPWR VPWR _20203_/A sky130_fd_sc_hd__buf_12
X_30560_ _30560_/A VGND VGND VPWR VPWR _35514_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29219_ input50/X VGND VGND VPWR VPWR _29219_/X sky130_fd_sc_hd__buf_2
XFILLER_187_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17233_ _33775_/Q _33711_/Q _33647_/Q _33583_/Q _17196_/X _17197_/X VGND VGND VPWR
+ VPWR _17233_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30491_ _30491_/A VGND VGND VPWR VPWR _35481_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_74_CLK clkbuf_leaf_76_CLK/A VGND VGND VPWR VPWR _33234_/CLK sky130_fd_sc_hd__clkbuf_16
X_32230_ _35852_/CLK _32230_/D VGND VGND VPWR VPWR _32230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17164_ _17164_/A VGND VGND VPWR VPWR _31980_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16115_ _16014_/X _16113_/X _16114_/X _16023_/X VGND VGND VPWR VPWR _16115_/X sky130_fd_sc_hd__a22o_1
XFILLER_183_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32161_ _34271_/CLK _32161_/D VGND VGND VPWR VPWR _32161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17095_ _16849_/X _17093_/X _17094_/X _16852_/X VGND VGND VPWR VPWR _17095_/X sky130_fd_sc_hd__a22o_1
X_31112_ _35776_/Q _29206_/X _31130_/S VGND VGND VPWR VPWR _31113_/A sky130_fd_sc_hd__mux2_1
X_16046_ _17796_/A VGND VGND VPWR VPWR _16046_/X sky130_fd_sc_hd__buf_6
XFILLER_115_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32092_ _35040_/CLK _32092_/D VGND VGND VPWR VPWR _32092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35920_ _35921_/CLK _35920_/D VGND VGND VPWR VPWR _35920_/Q sky130_fd_sc_hd__dfxtp_1
X_31043_ _31043_/A VGND VGND VPWR VPWR _35743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19805_ _20158_/A VGND VGND VPWR VPWR _19805_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35851_ _35851_/CLK _35851_/D VGND VGND VPWR VPWR _35851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17997_ _35332_/Q _35268_/Q _35204_/Q _32324_/Q _17712_/X _17713_/X VGND VGND VPWR
+ VPWR _17997_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34802_ _35061_/CLK _34802_/D VGND VGND VPWR VPWR _34802_/Q sky130_fd_sc_hd__dfxtp_1
X_19736_ _35060_/Q _34996_/Q _34932_/Q _34868_/Q _19456_/X _19457_/X VGND VGND VPWR
+ VPWR _19736_/X sky130_fd_sc_hd__mux4_1
X_16948_ _16842_/X _16946_/X _16947_/X _16847_/X VGND VGND VPWR VPWR _16948_/X sky130_fd_sc_hd__a22o_1
X_35782_ _35845_/CLK _35782_/D VGND VGND VPWR VPWR _35782_/Q sky130_fd_sc_hd__dfxtp_1
X_32994_ _32994_/CLK _32994_/D VGND VGND VPWR VPWR _32994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34733_ _35304_/CLK _34733_/D VGND VGND VPWR VPWR _34733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31945_ _31945_/A VGND VGND VPWR VPWR _36171_/D sky130_fd_sc_hd__clkbuf_1
X_16879_ _16879_/A VGND VGND VPWR VPWR _31972_/D sky130_fd_sc_hd__clkbuf_1
X_19667_ _19667_/A _19667_/B _19667_/C _19667_/D VGND VGND VPWR VPWR _19668_/A sky130_fd_sc_hd__or4_2
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18618_ _18612_/X _18617_/X _18311_/X VGND VGND VPWR VPWR _18640_/A sky130_fd_sc_hd__o21ba_1
XFILLER_53_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19598_ _19598_/A VGND VGND VPWR VPWR _32112_/D sky130_fd_sc_hd__buf_2
X_34664_ _34922_/CLK _34664_/D VGND VGND VPWR VPWR _34664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31876_ _31876_/A VGND VGND VPWR VPWR _36138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33615_ _34256_/CLK _33615_/D VGND VGND VPWR VPWR _33615_/Q sky130_fd_sc_hd__dfxtp_1
X_30827_ _23280_/X _35641_/Q _30839_/S VGND VGND VPWR VPWR _30828_/A sky130_fd_sc_hd__mux2_1
X_18549_ _18314_/X _18547_/X _18548_/X _18323_/X VGND VGND VPWR VPWR _18549_/X sky130_fd_sc_hd__a22o_1
XFILLER_244_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34595_ _35928_/CLK _34595_/D VGND VGND VPWR VPWR _34595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21560_ _22395_/A VGND VGND VPWR VPWR _21560_/X sky130_fd_sc_hd__buf_4
X_33546_ _36107_/CLK _33546_/D VGND VGND VPWR VPWR _33546_/Q sky130_fd_sc_hd__dfxtp_1
X_30758_ _23117_/X _35608_/Q _30776_/S VGND VGND VPWR VPWR _30759_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20511_ _18356_/X _20509_/X _20510_/X _18368_/X VGND VGND VPWR VPWR _20511_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33477_ _34050_/CLK _33477_/D VGND VGND VPWR VPWR _33477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21491_ _32997_/Q _32933_/Q _32869_/Q _32805_/Q _21236_/X _21237_/X VGND VGND VPWR
+ VPWR _21491_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_65_CLK clkbuf_leaf_66_CLK/A VGND VGND VPWR VPWR _32983_/CLK sky130_fd_sc_hd__clkbuf_16
X_30689_ _30689_/A VGND VGND VPWR VPWR _35575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23230_ _23230_/A VGND VGND VPWR VPWR _32194_/D sky130_fd_sc_hd__clkbuf_1
X_20442_ _35593_/Q _35529_/Q _35465_/Q _35401_/Q _20256_/X _20257_/X VGND VGND VPWR
+ VPWR _20442_/X sky130_fd_sc_hd__mux4_1
X_35216_ _35281_/CLK _35216_/D VGND VGND VPWR VPWR _35216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32428_ _35500_/CLK _32428_/D VGND VGND VPWR VPWR _32428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36196_ _36196_/CLK _36196_/D VGND VGND VPWR VPWR _36196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23161_ _32164_/Q _23077_/X _23182_/S VGND VGND VPWR VPWR _23162_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35147_ _35147_/CLK _35147_/D VGND VGND VPWR VPWR _35147_/Q sky130_fd_sc_hd__dfxtp_1
X_20373_ _33287_/Q _36167_/Q _33159_/Q _33095_/Q _20064_/X _20065_/X VGND VGND VPWR
+ VPWR _20373_/X sky130_fd_sc_hd__mux4_1
X_32359_ _34792_/CLK _32359_/D VGND VGND VPWR VPWR _32359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22112_ _22465_/A VGND VGND VPWR VPWR _22112_/X sky130_fd_sc_hd__buf_2
XFILLER_88_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35078_ _35078_/CLK _35078_/D VGND VGND VPWR VPWR _35078_/Q sky130_fd_sc_hd__dfxtp_1
X_23092_ _23092_/A VGND VGND VPWR VPWR _32143_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22043_ _22557_/A VGND VGND VPWR VPWR _22043_/X sky130_fd_sc_hd__buf_4
X_26920_ _26919_/X _33837_/Q _26944_/S VGND VGND VPWR VPWR _26921_/A sky130_fd_sc_hd__mux2_1
X_34029_ _36085_/CLK _34029_/D VGND VGND VPWR VPWR _34029_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26851_ _26850_/X _33815_/Q _26851_/S VGND VGND VPWR VPWR _26852_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25802_ _25802_/A VGND VGND VPWR VPWR _33323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29570_ _29570_/A VGND VGND VPWR VPWR _35045_/D sky130_fd_sc_hd__clkbuf_1
X_26782_ _33787_/Q _24385_/X _26790_/S VGND VGND VPWR VPWR _26783_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23994_ _23994_/A VGND VGND VPWR VPWR _32535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28521_ _28521_/A VGND VGND VPWR VPWR _34579_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25733_ _33292_/Q _24437_/X _25735_/S VGND VGND VPWR VPWR _25734_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22945_ input14/X VGND VGND VPWR VPWR _22945_/X sky130_fd_sc_hd__buf_2
XFILLER_90_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28452_ _26937_/X _34547_/Q _28456_/S VGND VGND VPWR VPWR _28453_/A sky130_fd_sc_hd__mux2_1
X_25664_ _33259_/Q _24335_/X _25664_/S VGND VGND VPWR VPWR _25665_/A sky130_fd_sc_hd__mux2_1
X_22876_ input85/X input84/X VGND VGND VPWR VPWR _31545_/A sky130_fd_sc_hd__nand2_8
XFILLER_55_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27403_ _27403_/A VGND VGND VPWR VPWR _34050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24615_ _22926_/X _32797_/Q _24623_/S VGND VGND VPWR VPWR _24616_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28383_ _26835_/X _34514_/Q _28393_/S VGND VGND VPWR VPWR _28384_/A sky130_fd_sc_hd__mux2_1
X_21827_ _34542_/Q _32430_/Q _34414_/Q _34350_/Q _21825_/X _21826_/X VGND VGND VPWR
+ VPWR _21827_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25595_ _33228_/Q _24437_/X _25597_/S VGND VGND VPWR VPWR _25596_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27334_ _27424_/S VGND VGND VPWR VPWR _27353_/S sky130_fd_sc_hd__buf_4
X_24546_ _23028_/X _32766_/Q _24548_/S VGND VGND VPWR VPWR _24547_/A sky130_fd_sc_hd__mux2_1
X_21758_ _35052_/Q _34988_/Q _34924_/Q _34860_/Q _21756_/X _21757_/X VGND VGND VPWR
+ VPWR _21758_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20709_ _22447_/A VGND VGND VPWR VPWR _20709_/X sky130_fd_sc_hd__buf_4
X_27265_ _26981_/X _33985_/Q _27281_/S VGND VGND VPWR VPWR _27266_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24477_ _22926_/X _32733_/Q _24485_/S VGND VGND VPWR VPWR _24478_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1030 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_931 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_CLK clkbuf_leaf_57_CLK/A VGND VGND VPWR VPWR _34276_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21689_ _22556_/A VGND VGND VPWR VPWR _21689_/X sky130_fd_sc_hd__buf_6
X_29004_ _29004_/A VGND VGND VPWR VPWR _34808_/D sky130_fd_sc_hd__clkbuf_1
X_26216_ _26216_/A VGND VGND VPWR VPWR _33519_/D sky130_fd_sc_hd__clkbuf_1
X_23428_ _22875_/X _32270_/Q _23446_/S VGND VGND VPWR VPWR _23429_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27196_ _27196_/A VGND VGND VPWR VPWR _33952_/D sky130_fd_sc_hd__clkbuf_1
X_26147_ _26147_/A VGND VGND VPWR VPWR _33486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23359_ _32239_/Q _23247_/X _23371_/S VGND VGND VPWR VPWR _23360_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26078_ _25091_/X _33454_/Q _26092_/S VGND VGND VPWR VPWR _26079_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29906_ _35205_/Q _29222_/X _29914_/S VGND VGND VPWR VPWR _29907_/A sky130_fd_sc_hd__mux2_1
X_17920_ _17916_/X _17919_/X _17842_/X _17843_/X VGND VGND VPWR VPWR _17937_/B sky130_fd_sc_hd__o211a_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25029_ input4/X VGND VGND VPWR VPWR _25029_/X sky130_fd_sc_hd__buf_2
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17851_ _33216_/Q _32576_/Q _35968_/Q _35904_/Q _17780_/X _17781_/X VGND VGND VPWR
+ VPWR _17851_/X sky130_fd_sc_hd__mux4_1
XTAP_6963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29837_ _35172_/Q _29120_/X _29851_/S VGND VGND VPWR VPWR _29838_/A sky130_fd_sc_hd__mux2_1
XTAP_6974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_45__f_CLK clkbuf_5_22_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_45__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XTAP_6985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16802_ _34530_/Q _32418_/Q _34402_/Q _34338_/Q _16519_/X _16520_/X VGND VGND VPWR
+ VPWR _16802_/X sky130_fd_sc_hd__mux4_1
XTAP_6996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17782_ _33214_/Q _32574_/Q _35966_/Q _35902_/Q _17780_/X _17781_/X VGND VGND VPWR
+ VPWR _17782_/X sky130_fd_sc_hd__mux4_1
X_29768_ _29768_/A VGND VGND VPWR VPWR _35139_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19521_ _19517_/X _19520_/X _19447_/X VGND VGND VPWR VPWR _19531_/C sky130_fd_sc_hd__o21ba_1
X_16733_ _16733_/A _16733_/B _16733_/C _16733_/D VGND VGND VPWR VPWR _16734_/A sky130_fd_sc_hd__or4_1
X_28719_ _28719_/A VGND VGND VPWR VPWR _34673_/D sky130_fd_sc_hd__clkbuf_1
X_29699_ _29699_/A VGND VGND VPWR VPWR _35106_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19452_ _19452_/A VGND VGND VPWR VPWR _19452_/X sky130_fd_sc_hd__clkbuf_4
X_31730_ _36069_/Q input16/X _31742_/S VGND VGND VPWR VPWR _31731_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16664_ _34271_/Q _34207_/Q _34143_/Q _34079_/Q _16383_/X _16384_/X VGND VGND VPWR
+ VPWR _16664_/X sky130_fd_sc_hd__mux4_1
XFILLER_234_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18403_ _18403_/A VGND VGND VPWR VPWR _32078_/D sky130_fd_sc_hd__clkbuf_1
X_31661_ _31661_/A VGND VGND VPWR VPWR _36036_/D sky130_fd_sc_hd__clkbuf_1
X_19383_ _35050_/Q _34986_/Q _34922_/Q _34858_/Q _19103_/X _19104_/X VGND VGND VPWR
+ VPWR _19383_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16595_ _16489_/X _16593_/X _16594_/X _16494_/X VGND VGND VPWR VPWR _16595_/X sky130_fd_sc_hd__a22o_1
XFILLER_76_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18334_ _18359_/A VGND VGND VPWR VPWR _20130_/A sky130_fd_sc_hd__buf_12
X_30612_ _35539_/Q _29067_/X _30620_/S VGND VGND VPWR VPWR _30613_/A sky130_fd_sc_hd__mux2_1
X_33400_ _34297_/CLK _33400_/D VGND VGND VPWR VPWR _33400_/Q sky130_fd_sc_hd__dfxtp_1
X_34380_ _35981_/CLK _34380_/D VGND VGND VPWR VPWR _34380_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31592_ _31592_/A VGND VGND VPWR VPWR _36003_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33331_ _33779_/CLK _33331_/D VGND VGND VPWR VPWR _33331_/Q sky130_fd_sc_hd__dfxtp_1
X_18265_ _18261_/X _18264_/X _17853_/A VGND VGND VPWR VPWR _18273_/C sky130_fd_sc_hd__o21ba_1
X_30543_ _30543_/A VGND VGND VPWR VPWR _35506_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_47_CLK clkbuf_leaf_50_CLK/A VGND VGND VPWR VPWR _36065_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_204_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17216_ _35758_/Q _35118_/Q _34478_/Q _33838_/Q _17140_/X _17141_/X VGND VGND VPWR
+ VPWR _17216_/X sky130_fd_sc_hd__mux4_1
XFILLER_198_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36050_ _36050_/CLK _36050_/D VGND VGND VPWR VPWR _36050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33262_ _33262_/CLK _33262_/D VGND VGND VPWR VPWR _33262_/Q sky130_fd_sc_hd__dfxtp_1
X_18196_ _33035_/Q _32971_/Q _32907_/Q _32843_/Q _15980_/X _15983_/X VGND VGND VPWR
+ VPWR _18196_/X sky130_fd_sc_hd__mux4_1
X_30474_ _30474_/A VGND VGND VPWR VPWR _35473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32213_ _35965_/CLK _32213_/D VGND VGND VPWR VPWR _32213_/Q sky130_fd_sc_hd__dfxtp_1
X_35001_ _35386_/CLK _35001_/D VGND VGND VPWR VPWR _35001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17147_ _17853_/A VGND VGND VPWR VPWR _17147_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33193_ _35947_/CLK _33193_/D VGND VGND VPWR VPWR _33193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32144_ _34001_/CLK _32144_/D VGND VGND VPWR VPWR _32144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17078_ _17072_/X _17077_/X _16794_/X VGND VGND VPWR VPWR _17086_/C sky130_fd_sc_hd__o21ba_1
X_16029_ _16059_/A VGND VGND VPWR VPWR _17770_/A sky130_fd_sc_hd__buf_12
XFILLER_130_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32075_ _36172_/CLK _32075_/D VGND VGND VPWR VPWR _32075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35903_ _35903_/CLK _35903_/D VGND VGND VPWR VPWR _35903_/Q sky130_fd_sc_hd__dfxtp_1
X_31026_ _31026_/A VGND VGND VPWR VPWR _35735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35834_ _35834_/CLK _35834_/D VGND VGND VPWR VPWR _35834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19719_ _33012_/Q _32948_/Q _32884_/Q _32820_/Q _19642_/X _19643_/X VGND VGND VPWR
+ VPWR _19719_/X sky130_fd_sc_hd__mux4_1
XFILLER_211_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20991_ _32727_/Q _32663_/Q _32599_/Q _36055_/Q _20813_/X _20950_/X VGND VGND VPWR
+ VPWR _20991_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35765_ _35765_/CLK _35765_/D VGND VGND VPWR VPWR _35765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32977_ _36049_/CLK _32977_/D VGND VGND VPWR VPWR _32977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22730_ _22508_/X _22728_/X _22729_/X _22511_/X VGND VGND VPWR VPWR _22730_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34716_ _34782_/CLK _34716_/D VGND VGND VPWR VPWR _34716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31928_ _23313_/X _36163_/Q _31940_/S VGND VGND VPWR VPWR _31929_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35696_ _35951_/CLK _35696_/D VGND VGND VPWR VPWR _35696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22661_ _22460_/X _22659_/X _22660_/X _22465_/X VGND VGND VPWR VPWR _22661_/X sky130_fd_sc_hd__a22o_1
X_34647_ _36202_/CLK _34647_/D VGND VGND VPWR VPWR _34647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31859_ _23148_/X _36130_/Q _31877_/S VGND VGND VPWR VPWR _31860_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24400_ input46/X VGND VGND VPWR VPWR _24400_/X sky130_fd_sc_hd__buf_4
XFILLER_222_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21612_ _21401_/X _21610_/X _21611_/X _21406_/X VGND VGND VPWR VPWR _21612_/X sky130_fd_sc_hd__a22o_1
X_25380_ _25380_/A VGND VGND VPWR VPWR _33127_/D sky130_fd_sc_hd__clkbuf_1
X_22592_ _22305_/X _22590_/X _22591_/X _22308_/X VGND VGND VPWR VPWR _22592_/X sky130_fd_sc_hd__a22o_1
X_34578_ _34706_/CLK _34578_/D VGND VGND VPWR VPWR _34578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24331_ _24331_/A VGND VGND VPWR VPWR _32681_/D sky130_fd_sc_hd__clkbuf_1
X_33529_ _34298_/CLK _33529_/D VGND VGND VPWR VPWR _33529_/Q sky130_fd_sc_hd__dfxtp_1
X_21543_ _21539_/X _21542_/X _21408_/X VGND VGND VPWR VPWR _21544_/D sky130_fd_sc_hd__o21ba_1
XFILLER_107_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_38_CLK clkbuf_6_7__f_CLK/X VGND VGND VPWR VPWR _36121_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_166_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27050_ _26863_/X _33883_/Q _27062_/S VGND VGND VPWR VPWR _27051_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24262_ _32659_/Q _24261_/X _24274_/S VGND VGND VPWR VPWR _24263_/A sky130_fd_sc_hd__mux2_1
X_21474_ _34532_/Q _32420_/Q _34404_/Q _34340_/Q _21472_/X _21473_/X VGND VGND VPWR
+ VPWR _21474_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26001_ _25177_/X _33418_/Q _26007_/S VGND VGND VPWR VPWR _26002_/A sky130_fd_sc_hd__mux2_1
X_20425_ _33801_/Q _33737_/Q _33673_/Q _33609_/Q _20202_/X _20203_/X VGND VGND VPWR
+ VPWR _20425_/X sky130_fd_sc_hd__mux4_1
X_23213_ _32188_/Q _23175_/X _23235_/S VGND VGND VPWR VPWR _23214_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36179_ _36202_/CLK _36179_/D VGND VGND VPWR VPWR _36179_/Q sky130_fd_sc_hd__dfxtp_1
X_24193_ _24193_/A VGND VGND VPWR VPWR _32629_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20356_ _34822_/Q _34758_/Q _34694_/Q _34630_/Q _20294_/X _20295_/X VGND VGND VPWR
+ VPWR _20356_/X sky130_fd_sc_hd__mux4_1
XFILLER_218_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23144_ _23144_/A VGND VGND VPWR VPWR _32160_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27952_ _34310_/Q _24419_/X _27958_/S VGND VGND VPWR VPWR _27953_/A sky130_fd_sc_hd__mux2_1
X_23075_ _23074_/X _32077_/Q _23075_/S VGND VGND VPWR VPWR _23076_/A sky130_fd_sc_hd__mux2_1
XTAP_6215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20287_ _35844_/Q _32223_/Q _35716_/Q _35652_/Q _19966_/X _19967_/X VGND VGND VPWR
+ VPWR _20287_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26903_ input19/X VGND VGND VPWR VPWR _26903_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_66_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22026_ _35572_/Q _35508_/Q _35444_/Q _35380_/Q _21850_/X _21851_/X VGND VGND VPWR
+ VPWR _22026_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27883_ _34277_/Q _24317_/X _27895_/S VGND VGND VPWR VPWR _27884_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26834_ _26834_/A VGND VGND VPWR VPWR _33809_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29622_ _29622_/A VGND VGND VPWR VPWR _35070_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29553_ _29553_/A VGND VGND VPWR VPWR _35037_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26765_ _33779_/Q _24360_/X _26769_/S VGND VGND VPWR VPWR _26766_/A sky130_fd_sc_hd__mux2_1
X_23977_ _22883_/X _32527_/Q _23993_/S VGND VGND VPWR VPWR _23978_/A sky130_fd_sc_hd__mux2_1
XTAP_4879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28504_ _27014_/X _34572_/Q _28506_/S VGND VGND VPWR VPWR _28505_/A sky130_fd_sc_hd__mux2_1
X_25716_ _25716_/A VGND VGND VPWR VPWR _33283_/D sky130_fd_sc_hd__clkbuf_1
X_29484_ _23294_/X _35005_/Q _29488_/S VGND VGND VPWR VPWR _29485_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22928_ _22928_/A VGND VGND VPWR VPWR _32029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26696_ _33746_/Q _24258_/X _26706_/S VGND VGND VPWR VPWR _26697_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28435_ _26912_/X _34539_/Q _28435_/S VGND VGND VPWR VPWR _28436_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25647_ _25647_/A VGND VGND VPWR VPWR _33250_/D sky130_fd_sc_hd__clkbuf_1
X_22859_ _35853_/Q _32233_/Q _35725_/Q _35661_/Q _20589_/X _20591_/X VGND VGND VPWR
+ VPWR _22859_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28366_ _28366_/A VGND VGND VPWR VPWR _34506_/D sky130_fd_sc_hd__clkbuf_1
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16380_ _16380_/A _16380_/B _16380_/C _16380_/D VGND VGND VPWR VPWR _16381_/A sky130_fd_sc_hd__or4_4
X_25578_ _25578_/A VGND VGND VPWR VPWR _33219_/D sky130_fd_sc_hd__clkbuf_1
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27317_ _27317_/A VGND VGND VPWR VPWR _34009_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24529_ _24577_/S VGND VGND VPWR VPWR _24548_/S sky130_fd_sc_hd__buf_4
XFILLER_200_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28297_ _28297_/A VGND VGND VPWR VPWR _34473_/D sky130_fd_sc_hd__clkbuf_1
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_29_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _34202_/CLK sky130_fd_sc_hd__clkbuf_16
X_18050_ _35782_/Q _35142_/Q _34502_/Q _33862_/Q _17846_/X _17847_/X VGND VGND VPWR
+ VPWR _18050_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27248_ _26956_/X _33977_/Q _27260_/S VGND VGND VPWR VPWR _27249_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17001_ _33192_/Q _32552_/Q _35944_/Q _35880_/Q _16721_/X _16722_/X VGND VGND VPWR
+ VPWR _17001_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27179_ _26853_/X _33944_/Q _27197_/S VGND VGND VPWR VPWR _27180_/A sky130_fd_sc_hd__mux2_1
XANTENNA_7 _32114_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30190_ _35340_/Q _29243_/X _30192_/S VGND VGND VPWR VPWR _30191_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18952_ _34782_/Q _34718_/Q _34654_/Q _34590_/Q _18882_/X _18883_/X VGND VGND VPWR
+ VPWR _18952_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17903_ _17903_/A VGND VGND VPWR VPWR _17903_/X sky130_fd_sc_hd__buf_6
XFILLER_156_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18883_ _20295_/A VGND VGND VPWR VPWR _18883_/X sky130_fd_sc_hd__buf_4
XTAP_6760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32900_ _36103_/CLK _32900_/D VGND VGND VPWR VPWR _32900_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17834_ _17834_/A VGND VGND VPWR VPWR _17834_/X sky130_fd_sc_hd__buf_2
XFILLER_117_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33880_ _36185_/CLK _33880_/D VGND VGND VPWR VPWR _33880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32831_ _36033_/CLK _32831_/D VGND VGND VPWR VPWR _32831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17765_ _17770_/A VGND VGND VPWR VPWR _17765_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_66_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19504_ _34030_/Q _33966_/Q _33902_/Q _32238_/Q _19320_/X _19321_/X VGND VGND VPWR
+ VPWR _19504_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35550_ _35744_/CLK _35550_/D VGND VGND VPWR VPWR _35550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16716_ _16709_/X _16715_/X _16430_/X _16431_/X VGND VGND VPWR VPWR _16733_/B sky130_fd_sc_hd__o211a_2
XFILLER_78_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17696_ _17830_/A VGND VGND VPWR VPWR _17696_/X sky130_fd_sc_hd__clkbuf_4
X_32762_ _36090_/CLK _32762_/D VGND VGND VPWR VPWR _32762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34501_ _35845_/CLK _34501_/D VGND VGND VPWR VPWR _34501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16647_ _35550_/Q _35486_/Q _35422_/Q _35358_/Q _16544_/X _16545_/X VGND VGND VPWR
+ VPWR _16647_/X sky130_fd_sc_hd__mux4_1
X_19435_ _19363_/X _19433_/X _19434_/X _19367_/X VGND VGND VPWR VPWR _19435_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31713_ _36061_/Q input7/X _31721_/S VGND VGND VPWR VPWR _31714_/A sky130_fd_sc_hd__mux2_1
X_35481_ _35481_/CLK _35481_/D VGND VGND VPWR VPWR _35481_/Q sky130_fd_sc_hd__dfxtp_1
X_32693_ _36085_/CLK _32693_/D VGND VGND VPWR VPWR _32693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34432_ _35777_/CLK _34432_/D VGND VGND VPWR VPWR _34432_/Q sky130_fd_sc_hd__dfxtp_1
X_31644_ _31644_/A VGND VGND VPWR VPWR _36028_/D sky130_fd_sc_hd__clkbuf_1
X_16578_ _35548_/Q _35484_/Q _35420_/Q _35356_/Q _16544_/X _16545_/X VGND VGND VPWR
+ VPWR _16578_/X sky130_fd_sc_hd__mux4_1
X_19366_ _33002_/Q _32938_/Q _32874_/Q _32810_/Q _19289_/X _19290_/X VGND VGND VPWR
+ VPWR _19366_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18317_ _18359_/A VGND VGND VPWR VPWR _20062_/A sky130_fd_sc_hd__buf_12
X_34363_ _35579_/CLK _34363_/D VGND VGND VPWR VPWR _34363_/Q sky130_fd_sc_hd__dfxtp_1
X_31575_ _31575_/A VGND VGND VPWR VPWR _35995_/D sky130_fd_sc_hd__clkbuf_1
X_19297_ _20158_/A VGND VGND VPWR VPWR _19297_/X sky130_fd_sc_hd__buf_4
X_36102_ _36103_/CLK _36102_/D VGND VGND VPWR VPWR _36102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18248_ _33549_/Q _33485_/Q _33421_/Q _33357_/Q _16033_/X _16035_/X VGND VGND VPWR
+ VPWR _18248_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33314_ _33635_/CLK _33314_/D VGND VGND VPWR VPWR _33314_/Q sky130_fd_sc_hd__dfxtp_1
X_30526_ _30526_/A VGND VGND VPWR VPWR _35498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34294_ _34295_/CLK _34294_/D VGND VGND VPWR VPWR _34294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36033_ _36033_/CLK _36033_/D VGND VGND VPWR VPWR _36033_/Q sky130_fd_sc_hd__dfxtp_1
X_18179_ _34570_/Q _32458_/Q _34442_/Q _34378_/Q _17931_/X _17932_/X VGND VGND VPWR
+ VPWR _18179_/X sky130_fd_sc_hd__mux4_1
X_30457_ _23336_/X _35466_/Q _30463_/S VGND VGND VPWR VPWR _30458_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33245_ _34016_/CLK _33245_/D VGND VGND VPWR VPWR _33245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20210_ _34050_/Q _33986_/Q _33922_/Q _32258_/Q _20026_/X _20027_/X VGND VGND VPWR
+ VPWR _20210_/X sky130_fd_sc_hd__mux4_1
X_21190_ _21186_/X _21189_/X _21055_/X VGND VGND VPWR VPWR _21191_/D sky130_fd_sc_hd__o21ba_1
X_33176_ _35864_/CLK _33176_/D VGND VGND VPWR VPWR _33176_/Q sky130_fd_sc_hd__dfxtp_1
X_30388_ _23228_/X _35433_/Q _30392_/S VGND VGND VPWR VPWR _30389_/A sky130_fd_sc_hd__mux2_1
X_20141_ _20069_/X _20139_/X _20140_/X _20073_/X VGND VGND VPWR VPWR _20141_/X sky130_fd_sc_hd__a22o_1
X_32127_ _35949_/CLK _32127_/D VGND VGND VPWR VPWR _32127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20072_ _33022_/Q _32958_/Q _32894_/Q _32830_/Q _19995_/X _19996_/X VGND VGND VPWR
+ VPWR _20072_/X sky130_fd_sc_hd__mux4_1
X_32058_ _36027_/CLK _32058_/D VGND VGND VPWR VPWR _32058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31009_ _35727_/Q _29055_/X _31025_/S VGND VGND VPWR VPWR _31010_/A sky130_fd_sc_hd__mux2_1
XTAP_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23900_ _23900_/A VGND VGND VPWR VPWR _32491_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24880_ _24880_/A VGND VGND VPWR VPWR _32921_/D sky130_fd_sc_hd__clkbuf_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23831_ _23831_/A VGND VGND VPWR VPWR _32459_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35817_ _35818_/CLK _35817_/D VGND VGND VPWR VPWR _35817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_408 _36211_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26550_ _31815_/A _26685_/B VGND VGND VPWR VPWR _26683_/S sky130_fd_sc_hd__nand2_8
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35748_ _35748_/CLK _35748_/D VGND VGND VPWR VPWR _35748_/Q sky130_fd_sc_hd__dfxtp_1
X_23762_ _23762_/A VGND VGND VPWR VPWR _32426_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20974_ _35286_/Q _35222_/Q _35158_/Q _32278_/Q _20900_/X _20901_/X VGND VGND VPWR
+ VPWR _20974_/X sky130_fd_sc_hd__mux4_1
XANTENNA_419 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25501_ _33183_/Q _24298_/X _25505_/S VGND VGND VPWR VPWR _25502_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22713_ _33224_/Q _32584_/Q _35976_/Q _35912_/Q _20675_/X _20676_/X VGND VGND VPWR
+ VPWR _22713_/X sky130_fd_sc_hd__mux4_1
XFILLER_246_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26481_ _25088_/X _33645_/Q _26497_/S VGND VGND VPWR VPWR _26482_/A sky130_fd_sc_hd__mux2_1
X_23693_ _23693_/A VGND VGND VPWR VPWR _32395_/D sky130_fd_sc_hd__clkbuf_1
X_35679_ _35807_/CLK _35679_/D VGND VGND VPWR VPWR _35679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28220_ _26993_/X _34437_/Q _28228_/S VGND VGND VPWR VPWR _28221_/A sky130_fd_sc_hd__mux2_1
X_25432_ _25146_/X _33152_/Q _25450_/S VGND VGND VPWR VPWR _25433_/A sky130_fd_sc_hd__mux2_1
X_22644_ _22361_/X _22642_/X _22643_/X _22367_/X VGND VGND VPWR VPWR _22644_/X sky130_fd_sc_hd__a22o_1
XFILLER_224_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28151_ _26891_/X _34404_/Q _28165_/S VGND VGND VPWR VPWR _28152_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25363_ _25363_/A VGND VGND VPWR VPWR _33119_/D sky130_fd_sc_hd__clkbuf_1
X_22575_ _34052_/Q _33988_/Q _33924_/Q _32260_/Q _22326_/X _22327_/X VGND VGND VPWR
+ VPWR _22575_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_9__f_CLK clkbuf_5_4_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_9__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_178_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27102_ _26940_/X _33908_/Q _27104_/S VGND VGND VPWR VPWR _27103_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24314_ input15/X VGND VGND VPWR VPWR _24314_/X sky130_fd_sc_hd__buf_4
XFILLER_103_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28082_ _28082_/A VGND VGND VPWR VPWR _34371_/D sky130_fd_sc_hd__clkbuf_1
X_21526_ _21310_/X _21524_/X _21525_/X _21314_/X VGND VGND VPWR VPWR _21526_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25294_ _25294_/A VGND VGND VPWR VPWR _33087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27033_ _26838_/X _33875_/Q _27041_/S VGND VGND VPWR VPWR _27034_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24245_ input85/X input84/X _31680_/B VGND VGND VPWR VPWR _24401_/A sky130_fd_sc_hd__nor3_4
XFILLER_147_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21457_ _21302_/X _21455_/X _21456_/X _21308_/X VGND VGND VPWR VPWR _21457_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20408_ _20404_/X _20407_/X _20142_/X _20143_/X VGND VGND VPWR VPWR _20423_/B sky130_fd_sc_hd__o211a_1
XFILLER_218_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21388_ _22595_/A VGND VGND VPWR VPWR _21388_/X sky130_fd_sc_hd__clkbuf_4
X_24176_ _22976_/X _32621_/Q _24192_/S VGND VGND VPWR VPWR _24177_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23127_ input5/X VGND VGND VPWR VPWR _23127_/X sky130_fd_sc_hd__buf_6
X_20339_ _34054_/Q _33990_/Q _33926_/Q _32262_/Q _20026_/X _20027_/X VGND VGND VPWR
+ VPWR _20339_/X sky130_fd_sc_hd__mux4_1
XTAP_6001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28984_ _34799_/Q _24348_/X _28996_/S VGND VGND VPWR VPWR _28985_/A sky130_fd_sc_hd__mux2_1
XTAP_6023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23058_ _23058_/A VGND VGND VPWR VPWR _32071_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27935_ _34302_/Q _24394_/X _27937_/S VGND VGND VPWR VPWR _27936_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput99 _31968_/Q VGND VGND VPWR VPWR D1[18] sky130_fd_sc_hd__buf_2
XTAP_6067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22009_ _22362_/A VGND VGND VPWR VPWR _22009_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_102_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27866_ _34269_/Q _24292_/X _27874_/S VGND VGND VPWR VPWR _27867_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29605_ _35062_/Q _29175_/X _29623_/S VGND VGND VPWR VPWR _29606_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26817_ _33804_/Q _24437_/X _26819_/S VGND VGND VPWR VPWR _26818_/A sky130_fd_sc_hd__mux2_1
XTAP_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27797_ _27797_/A VGND VGND VPWR VPWR _34236_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17550_ _17903_/A VGND VGND VPWR VPWR _17550_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29536_ _29536_/A VGND VGND VPWR VPWR _35029_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26748_ _33771_/Q _24335_/X _26748_/S VGND VGND VPWR VPWR _26749_/A sky130_fd_sc_hd__mux2_1
XTAP_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_920 _27005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16501_ _16495_/X _16500_/X _16422_/X VGND VGND VPWR VPWR _16525_/A sky130_fd_sc_hd__o21ba_1
XFILLER_229_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_931 _29247_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17481_ _17834_/A VGND VGND VPWR VPWR _17481_/X sky130_fd_sc_hd__buf_2
XTAP_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_942 _29382_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29467_ _23267_/X _34997_/Q _29467_/S VGND VGND VPWR VPWR _29468_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26679_ _25180_/X _33739_/Q _26683_/S VGND VGND VPWR VPWR _26680_/A sky130_fd_sc_hd__mux2_1
XANTENNA_953 _29652_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_964 _30868_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16432_ _16426_/X _16429_/X _16430_/X _16431_/X VGND VGND VPWR VPWR _16457_/B sky130_fd_sc_hd__o211a_2
X_19220_ _32742_/Q _32678_/Q _32614_/Q _36070_/Q _19219_/X _19003_/X VGND VGND VPWR
+ VPWR _19220_/X sky130_fd_sc_hd__mux4_1
XANTENNA_975 _31948_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_986 _17796_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28418_ _28418_/A VGND VGND VPWR VPWR _34530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29398_ _23105_/X _34964_/Q _29404_/S VGND VGND VPWR VPWR _29399_/A sky130_fd_sc_hd__mux2_1
XANTENNA_997 _17956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_968 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19151_ _34020_/Q _33956_/Q _33892_/Q _32171_/Q _18967_/X _18968_/X VGND VGND VPWR
+ VPWR _19151_/X sky130_fd_sc_hd__mux4_1
X_28349_ _34498_/Q _24407_/X _28363_/S VGND VGND VPWR VPWR _28350_/A sky130_fd_sc_hd__mux2_1
X_16363_ _16356_/X _16362_/X _16040_/X _16042_/X VGND VGND VPWR VPWR _16380_/B sky130_fd_sc_hd__o211a_1
XFILLER_13_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18102_ _32776_/Q _32712_/Q _32648_/Q _36104_/Q _17978_/X _16873_/A VGND VGND VPWR
+ VPWR _18102_/X sky130_fd_sc_hd__mux4_1
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31360_ _31408_/S VGND VGND VPWR VPWR _31379_/S sky130_fd_sc_hd__buf_4
XFILLER_118_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19082_ _19010_/X _19080_/X _19081_/X _19014_/X VGND VGND VPWR VPWR _19082_/X sky130_fd_sc_hd__a22o_1
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16294_ _35540_/Q _35476_/Q _35412_/Q _35348_/Q _16191_/X _16192_/X VGND VGND VPWR
+ VPWR _16294_/X sky130_fd_sc_hd__mux4_1
XFILLER_199_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18033_ _18033_/A _18033_/B _18033_/C _18033_/D VGND VGND VPWR VPWR _18034_/A sky130_fd_sc_hd__or4_4
XFILLER_201_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30311_ _35397_/Q _29222_/X _30319_/S VGND VGND VPWR VPWR _30312_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31291_ _35861_/Q input62/X _31295_/S VGND VGND VPWR VPWR _31292_/A sky130_fd_sc_hd__mux2_1
X_33030_ _36039_/CLK _33030_/D VGND VGND VPWR VPWR _33030_/Q sky130_fd_sc_hd__dfxtp_1
X_30242_ _35364_/Q _29120_/X _30256_/S VGND VGND VPWR VPWR _30243_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30173_ _30173_/A VGND VGND VPWR VPWR _35331_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19984_ _33788_/Q _33724_/Q _33660_/Q _33596_/Q _19849_/X _19850_/X VGND VGND VPWR
+ VPWR _19984_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18935_ _32478_/Q _32350_/Q _32030_/Q _35998_/Q _18870_/X _18658_/X VGND VGND VPWR
+ VPWR _18935_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34981_ _35042_/CLK _34981_/D VGND VGND VPWR VPWR _34981_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1330 _20146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1341 _22557_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1352 _21759_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33932_ _34316_/CLK _33932_/D VGND VGND VPWR VPWR _33932_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1363 _24267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_9_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _35292_/CLK sky130_fd_sc_hd__clkbuf_16
X_18866_ _20278_/A VGND VGND VPWR VPWR _18866_/X sky130_fd_sc_hd__buf_6
XTAP_6590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1374 _26412_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1385 _31273_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1396 input89/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17817_ _34815_/Q _34751_/Q _34687_/Q _34623_/Q _17641_/X _17642_/X VGND VGND VPWR
+ VPWR _17817_/X sky130_fd_sc_hd__mux4_1
X_33863_ _35847_/CLK _33863_/D VGND VGND VPWR VPWR _33863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18797_ _33498_/Q _33434_/Q _33370_/Q _33306_/Q _18717_/X _18718_/X VGND VGND VPWR
+ VPWR _18797_/X sky130_fd_sc_hd__mux4_1
XFILLER_212_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35602_ _35666_/CLK _35602_/D VGND VGND VPWR VPWR _35602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32814_ _33007_/CLK _32814_/D VGND VGND VPWR VPWR _32814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17748_ _34557_/Q _32445_/Q _34429_/Q _34365_/Q _17578_/X _17579_/X VGND VGND VPWR
+ VPWR _17748_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33794_ _34306_/CLK _33794_/D VGND VGND VPWR VPWR _33794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35533_ _35597_/CLK _35533_/D VGND VGND VPWR VPWR _35533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32745_ _36137_/CLK _32745_/D VGND VGND VPWR VPWR _32745_/Q sky130_fd_sc_hd__dfxtp_1
X_17679_ _35067_/Q _35003_/Q _34939_/Q _34875_/Q _17509_/X _17510_/X VGND VGND VPWR
+ VPWR _17679_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19418_ _19418_/A _19418_/B _19418_/C _19418_/D VGND VGND VPWR VPWR _19419_/A sky130_fd_sc_hd__or4_4
XFILLER_223_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35464_ _35464_/CLK _35464_/D VGND VGND VPWR VPWR _35464_/Q sky130_fd_sc_hd__dfxtp_1
X_20690_ _21473_/A VGND VGND VPWR VPWR _20690_/X sky130_fd_sc_hd__buf_4
XFILLER_211_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32676_ _36132_/CLK _32676_/D VGND VGND VPWR VPWR _32676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34415_ _35052_/CLK _34415_/D VGND VGND VPWR VPWR _34415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31627_ _31627_/A VGND VGND VPWR VPWR _36020_/D sky130_fd_sc_hd__clkbuf_1
X_19349_ _34282_/Q _34218_/Q _34154_/Q _34090_/Q _19036_/X _19037_/X VGND VGND VPWR
+ VPWR _19349_/X sky130_fd_sc_hd__mux4_1
X_35395_ _35973_/CLK _35395_/D VGND VGND VPWR VPWR _35395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22360_ _22356_/X _22359_/X _22081_/X VGND VGND VPWR VPWR _22392_/A sky130_fd_sc_hd__o21ba_2
X_34346_ _35050_/CLK _34346_/D VGND VGND VPWR VPWR _34346_/Q sky130_fd_sc_hd__dfxtp_1
X_31558_ _31558_/A VGND VGND VPWR VPWR _35987_/D sky130_fd_sc_hd__clkbuf_1
X_21311_ _22370_/A VGND VGND VPWR VPWR _21311_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_163_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22291_ _32764_/Q _32700_/Q _32636_/Q _36092_/Q _22225_/X _22009_/X VGND VGND VPWR
+ VPWR _22291_/X sky130_fd_sc_hd__mux4_1
X_30509_ _23148_/X _35490_/Q _30527_/S VGND VGND VPWR VPWR _30510_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34277_ _34277_/CLK _34277_/D VGND VGND VPWR VPWR _34277_/Q sky130_fd_sc_hd__dfxtp_1
X_31489_ _23261_/X _35955_/Q _31493_/S VGND VGND VPWR VPWR _31490_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36016_ _36077_/CLK _36016_/D VGND VGND VPWR VPWR _36016_/Q sky130_fd_sc_hd__dfxtp_1
X_21242_ _35806_/Q _32181_/Q _35678_/Q _35614_/Q _21207_/X _21208_/X VGND VGND VPWR
+ VPWR _21242_/X sky130_fd_sc_hd__mux4_1
X_24030_ _24030_/A VGND VGND VPWR VPWR _32552_/D sky130_fd_sc_hd__clkbuf_1
X_33228_ _35978_/CLK _33228_/D VGND VGND VPWR VPWR _33228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21173_ _20957_/X _21171_/X _21172_/X _20961_/X VGND VGND VPWR VPWR _21173_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33159_ _36167_/CLK _33159_/D VGND VGND VPWR VPWR _33159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20124_ _20124_/A _20124_/B _20124_/C _20124_/D VGND VGND VPWR VPWR _20125_/A sky130_fd_sc_hd__or4_1
XFILLER_137_1258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25981_ _25146_/X _33408_/Q _25999_/S VGND VGND VPWR VPWR _25982_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27720_ _27831_/S VGND VGND VPWR VPWR _27739_/S sky130_fd_sc_hd__buf_4
X_20055_ _34302_/Q _34238_/Q _34174_/Q _34110_/Q _19742_/X _19743_/X VGND VGND VPWR
+ VPWR _20055_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24932_ _24932_/A VGND VGND VPWR VPWR _32946_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27651_ _34167_/Q _24373_/X _27667_/S VGND VGND VPWR VPWR _27652_/A sky130_fd_sc_hd__mux2_1
X_24863_ _24863_/A VGND VGND VPWR VPWR _32913_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26602_ _25066_/X _33702_/Q _26612_/S VGND VGND VPWR VPWR _26603_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23814_ _23044_/X _32451_/Q _23826_/S VGND VGND VPWR VPWR _23815_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27582_ _27582_/A VGND VGND VPWR VPWR _34134_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24794_ _22988_/X _32881_/Q _24802_/S VGND VGND VPWR VPWR _24795_/A sky130_fd_sc_hd__mux2_1
XANTENNA_216 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_227 _32136_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29321_ _29321_/A VGND VGND VPWR VPWR _34927_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26533_ _25165_/X _33670_/Q _26539_/S VGND VGND VPWR VPWR _26534_/A sky130_fd_sc_hd__mux2_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23745_ _22941_/X _32418_/Q _23763_/S VGND VGND VPWR VPWR _23746_/A sky130_fd_sc_hd__mux2_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ _22508_/A VGND VGND VPWR VPWR _20957_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_249 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29252_ _29252_/A VGND VGND VPWR VPWR _34894_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26464_ _25063_/X _33637_/Q _26476_/S VGND VGND VPWR VPWR _26465_/A sky130_fd_sc_hd__mux2_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23676_ _32387_/Q _23313_/X _23688_/S VGND VGND VPWR VPWR _23677_/A sky130_fd_sc_hd__mux2_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20888_ _22455_/A VGND VGND VPWR VPWR _20888_/X sky130_fd_sc_hd__buf_4
XFILLER_186_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28203_ _26968_/X _34429_/Q _28207_/S VGND VGND VPWR VPWR _28204_/A sky130_fd_sc_hd__mux2_1
X_25415_ _25122_/X _33144_/Q _25429_/S VGND VGND VPWR VPWR _25416_/A sky130_fd_sc_hd__mux2_1
X_22627_ _35333_/Q _35269_/Q _35205_/Q _32325_/Q _22312_/X _22313_/X VGND VGND VPWR
+ VPWR _22627_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29183_ _34872_/Q _29182_/X _29204_/S VGND VGND VPWR VPWR _29184_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26395_ _26395_/A VGND VGND VPWR VPWR _33604_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28134_ _26866_/X _34396_/Q _28144_/S VGND VGND VPWR VPWR _28135_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25346_ _25346_/A VGND VGND VPWR VPWR _33111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22558_ _35587_/Q _35523_/Q _35459_/Q _35395_/Q _22556_/X _22557_/X VGND VGND VPWR
+ VPWR _22558_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28065_ _28065_/A VGND VGND VPWR VPWR _34363_/D sky130_fd_sc_hd__clkbuf_1
X_21509_ _21505_/X _21508_/X _21408_/X VGND VGND VPWR VPWR _21510_/D sky130_fd_sc_hd__o21ba_1
X_25277_ _25119_/X _33079_/Q _25293_/S VGND VGND VPWR VPWR _25278_/A sky130_fd_sc_hd__mux2_1
X_22489_ _33217_/Q _32577_/Q _35969_/Q _35905_/Q _22380_/X _22381_/X VGND VGND VPWR
+ VPWR _22489_/X sky130_fd_sc_hd__mux4_1
X_27016_ _27016_/A VGND VGND VPWR VPWR _33868_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24228_ _23053_/X _32646_/Q _24234_/S VGND VGND VPWR VPWR _24229_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24159_ _22951_/X _32613_/Q _24171_/S VGND VGND VPWR VPWR _24160_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16981_ _33512_/Q _33448_/Q _33384_/Q _33320_/Q _16770_/X _16771_/X VGND VGND VPWR
+ VPWR _16981_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28967_ _34791_/Q _24323_/X _28975_/S VGND VGND VPWR VPWR _28968_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18720_ _34008_/Q _33944_/Q _33880_/Q _32152_/Q _18614_/X _18615_/X VGND VGND VPWR
+ VPWR _18720_/X sky130_fd_sc_hd__mux4_1
XTAP_5130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27918_ _27966_/S VGND VGND VPWR VPWR _27937_/S sky130_fd_sc_hd__buf_4
XTAP_5141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28898_ _28898_/A VGND VGND VPWR VPWR _34758_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18651_ _32726_/Q _32662_/Q _32598_/Q _36054_/Q _18513_/X _18650_/X VGND VGND VPWR
+ VPWR _18651_/X sky130_fd_sc_hd__mux4_1
XFILLER_237_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27849_ _34261_/Q _24267_/X _27853_/S VGND VGND VPWR VPWR _27850_/A sky130_fd_sc_hd__mux2_1
XTAP_5185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ _17347_/X _17600_/X _17601_/X _17350_/X VGND VGND VPWR VPWR _17602_/X sky130_fd_sc_hd__a22o_1
XFILLER_76_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30860_ _23333_/X _35657_/Q _30860_/S VGND VGND VPWR VPWR _30861_/A sky130_fd_sc_hd__mux2_1
XTAP_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18582_ _32468_/Q _32340_/Q _32020_/Q _35988_/Q _18517_/X _20163_/A VGND VGND VPWR
+ VPWR _18582_/X sky130_fd_sc_hd__mux4_1
XTAP_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29519_ _30059_/A _30600_/B VGND VGND VPWR VPWR _29652_/S sky130_fd_sc_hd__nor2_8
XTAP_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ _35767_/Q _35127_/Q _34487_/Q _33847_/Q _17493_/X _17494_/X VGND VGND VPWR
+ VPWR _17533_/X sky130_fd_sc_hd__mux4_1
XTAP_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30791_ _23223_/X _35624_/Q _30797_/S VGND VGND VPWR VPWR _30792_/A sky130_fd_sc_hd__mux2_1
XANTENNA_750 _22393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_761 _22500_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_260_CLK clkbuf_6_60__f_CLK/X VGND VGND VPWR VPWR _32965_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_166_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_772 _22538_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32530_ _36112_/CLK _32530_/D VGND VGND VPWR VPWR _32530_/Q sky130_fd_sc_hd__dfxtp_1
X_17464_ _34805_/Q _34741_/Q _34677_/Q _34613_/Q _17288_/X _17289_/X VGND VGND VPWR
+ VPWR _17464_/X sky130_fd_sc_hd__mux4_1
XANTENNA_783 _22633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_794 _22724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16415_ _34264_/Q _34200_/Q _34136_/Q _34072_/Q _16383_/X _16384_/X VGND VGND VPWR
+ VPWR _16415_/X sky130_fd_sc_hd__mux4_1
X_19203_ _34789_/Q _34725_/Q _34661_/Q _34597_/Q _18882_/X _18883_/X VGND VGND VPWR
+ VPWR _19203_/X sky130_fd_sc_hd__mux4_1
X_32461_ _35981_/CLK _32461_/D VGND VGND VPWR VPWR _32461_/Q sky130_fd_sc_hd__dfxtp_1
X_17395_ _34547_/Q _32435_/Q _34419_/Q _34355_/Q _17225_/X _17226_/X VGND VGND VPWR
+ VPWR _17395_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34200_ _35284_/CLK _34200_/D VGND VGND VPWR VPWR _34200_/Q sky130_fd_sc_hd__dfxtp_1
X_16346_ _34006_/Q _33942_/Q _33878_/Q _32150_/Q _16314_/X _16315_/X VGND VGND VPWR
+ VPWR _16346_/X sky130_fd_sc_hd__mux4_1
X_31412_ _23077_/X _35918_/Q _31430_/S VGND VGND VPWR VPWR _31413_/A sky130_fd_sc_hd__mux2_1
X_19134_ _35299_/Q _35235_/Q _35171_/Q _32291_/Q _18953_/X _18954_/X VGND VGND VPWR
+ VPWR _19134_/X sky130_fd_sc_hd__mux4_1
X_32392_ _35975_/CLK _32392_/D VGND VGND VPWR VPWR _32392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35180_ _35308_/CLK _35180_/D VGND VGND VPWR VPWR _35180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34131_ _34260_/CLK _34131_/D VGND VGND VPWR VPWR _34131_/Q sky130_fd_sc_hd__dfxtp_1
X_19065_ _19065_/A _19065_/B _19065_/C _19065_/D VGND VGND VPWR VPWR _19066_/A sky130_fd_sc_hd__or4_1
X_31343_ _31343_/A VGND VGND VPWR VPWR _35885_/D sky130_fd_sc_hd__clkbuf_1
X_16277_ _16143_/X _16275_/X _16276_/X _16146_/X VGND VGND VPWR VPWR _16277_/X sky130_fd_sc_hd__a22o_1
XFILLER_160_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18016_ _33029_/Q _32965_/Q _32901_/Q _32837_/Q _17695_/X _17696_/X VGND VGND VPWR
+ VPWR _18016_/X sky130_fd_sc_hd__mux4_1
X_34062_ _35021_/CLK _34062_/D VGND VGND VPWR VPWR _34062_/Q sky130_fd_sc_hd__dfxtp_1
X_31274_ _31274_/A VGND VGND VPWR VPWR _35853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_13_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_13_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_126_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30225_ _35356_/Q _29095_/X _30235_/S VGND VGND VPWR VPWR _30226_/A sky130_fd_sc_hd__mux2_1
X_33013_ _33013_/CLK _33013_/D VGND VGND VPWR VPWR _33013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30156_ _30156_/A VGND VGND VPWR VPWR _35323_/D sky130_fd_sc_hd__clkbuf_1
X_19967_ _20096_/A VGND VGND VPWR VPWR _19967_/X sky130_fd_sc_hd__buf_4
XFILLER_214_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18918_ _18743_/X _18916_/X _18917_/X _18746_/X VGND VGND VPWR VPWR _18918_/X sky130_fd_sc_hd__a22o_1
X_34964_ _35031_/CLK _34964_/D VGND VGND VPWR VPWR _34964_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_28_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_28_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_41_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30087_ _30087_/A VGND VGND VPWR VPWR _35290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1160 _22511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19898_ _19716_/X _19896_/X _19897_/X _19720_/X VGND VGND VPWR VPWR _19898_/X sky130_fd_sc_hd__a22o_1
XFILLER_67_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1171 _22447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1182 _21664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33915_ _36154_/CLK _33915_/D VGND VGND VPWR VPWR _33915_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1193 _22901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18849_ _18843_/X _18848_/X _18741_/X VGND VGND VPWR VPWR _18857_/C sky130_fd_sc_hd__o21ba_1
X_34895_ _35026_/CLK _34895_/D VGND VGND VPWR VPWR _34895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33846_ _35766_/CLK _33846_/D VGND VGND VPWR VPWR _33846_/Q sky130_fd_sc_hd__dfxtp_1
X_21860_ _35055_/Q _34991_/Q _34927_/Q _34863_/Q _21756_/X _21757_/X VGND VGND VPWR
+ VPWR _21860_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20811_ _20743_/X _20809_/X _20810_/X _20746_/X VGND VGND VPWR VPWR _20811_/X sky130_fd_sc_hd__a22o_1
X_21791_ _21754_/X _21789_/X _21790_/X _21759_/X VGND VGND VPWR VPWR _21791_/X sky130_fd_sc_hd__a22o_1
X_33777_ _33779_/CLK _33777_/D VGND VGND VPWR VPWR _33777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30989_ _35718_/Q _29225_/X _30995_/S VGND VGND VPWR VPWR _30990_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_251_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _33545_/CLK sky130_fd_sc_hd__clkbuf_16
X_23530_ _23031_/X _32319_/Q _23530_/S VGND VGND VPWR VPWR _23531_/A sky130_fd_sc_hd__mux2_1
X_35516_ _35517_/CLK _35516_/D VGND VGND VPWR VPWR _35516_/Q sky130_fd_sc_hd__dfxtp_1
X_20742_ _20736_/X _20739_/X _20740_/X _20741_/X VGND VGND VPWR VPWR _20742_/X sky130_fd_sc_hd__a22o_1
XFILLER_180_1407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32728_ _36123_/CLK _32728_/D VGND VGND VPWR VPWR _32728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23461_ _22929_/X _32286_/Q _23467_/S VGND VGND VPWR VPWR _23462_/A sky130_fd_sc_hd__mux2_1
X_35447_ _35638_/CLK _35447_/D VGND VGND VPWR VPWR _35447_/Q sky130_fd_sc_hd__dfxtp_1
X_20673_ _22361_/A VGND VGND VPWR VPWR _21749_/A sky130_fd_sc_hd__clkbuf_16
X_32659_ _36050_/CLK _32659_/D VGND VGND VPWR VPWR _32659_/Q sky130_fd_sc_hd__dfxtp_1
X_25200_ _25200_/A VGND VGND VPWR VPWR _33042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22412_ _22300_/X _22410_/X _22411_/X _22303_/X VGND VGND VPWR VPWR _22412_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26180_ _26180_/A VGND VGND VPWR VPWR _33502_/D sky130_fd_sc_hd__clkbuf_1
X_23392_ _32255_/Q _23300_/X _23392_/S VGND VGND VPWR VPWR _23393_/A sky130_fd_sc_hd__mux2_1
X_35378_ _35826_/CLK _35378_/D VGND VGND VPWR VPWR _35378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25131_ input40/X VGND VGND VPWR VPWR _25131_/X sky130_fd_sc_hd__buf_2
XFILLER_137_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22343_ _22305_/X _22341_/X _22342_/X _22308_/X VGND VGND VPWR VPWR _22343_/X sky130_fd_sc_hd__a22o_1
X_34329_ _35293_/CLK _34329_/D VGND VGND VPWR VPWR _34329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25062_ _25062_/A VGND VGND VPWR VPWR _32996_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22274_ _22270_/X _22273_/X _22100_/X VGND VGND VPWR VPWR _22282_/C sky130_fd_sc_hd__o21ba_1
XFILLER_163_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24013_ _24013_/A VGND VGND VPWR VPWR _32544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21225_ _33758_/Q _33694_/Q _33630_/Q _33566_/Q _21090_/X _21091_/X VGND VGND VPWR
+ VPWR _21225_/X sky130_fd_sc_hd__mux4_1
X_29870_ _35188_/Q _29169_/X _29872_/S VGND VGND VPWR VPWR _29871_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28821_ _28911_/S VGND VGND VPWR VPWR _28840_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_219_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21156_ _21152_/X _21155_/X _21055_/X VGND VGND VPWR VPWR _21157_/D sky130_fd_sc_hd__o21ba_1
XFILLER_63_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20107_ _33023_/Q _32959_/Q _32895_/Q _32831_/Q _19995_/X _19996_/X VGND VGND VPWR
+ VPWR _20107_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28752_ _26981_/X _34689_/Q _28768_/S VGND VGND VPWR VPWR _28753_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21087_ _21087_/A _21087_/B _21087_/C _21087_/D VGND VGND VPWR VPWR _21088_/A sky130_fd_sc_hd__or4_1
X_25964_ _25122_/X _33400_/Q _25978_/S VGND VGND VPWR VPWR _25965_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27703_ _27703_/A VGND VGND VPWR VPWR _34191_/D sky130_fd_sc_hd__clkbuf_1
X_20038_ _35837_/Q _32216_/Q _35709_/Q _35645_/Q _19966_/X _19967_/X VGND VGND VPWR
+ VPWR _20038_/X sky130_fd_sc_hd__mux4_1
XFILLER_115_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24915_ _24915_/A VGND VGND VPWR VPWR _32938_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25895_ _25895_/A VGND VGND VPWR VPWR _33367_/D sky130_fd_sc_hd__clkbuf_1
X_28683_ _28683_/A VGND VGND VPWR VPWR _34656_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_490_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _35807_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24846_ _23065_/X _32906_/Q _24852_/S VGND VGND VPWR VPWR _24847_/A sky130_fd_sc_hd__mux2_1
X_27634_ _34159_/Q _24348_/X _27646_/S VGND VGND VPWR VPWR _27635_/A sky130_fd_sc_hd__mux2_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27565_ _34126_/Q _24244_/X _27583_/S VGND VGND VPWR VPWR _27566_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24777_ _22963_/X _32873_/Q _24781_/S VGND VGND VPWR VPWR _24778_/A sky130_fd_sc_hd__mux2_1
X_21989_ _33203_/Q _32563_/Q _35955_/Q _35891_/Q _21674_/X _21675_/X VGND VGND VPWR
+ VPWR _21989_/X sky130_fd_sc_hd__mux4_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_242_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _34243_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26516_ _25140_/X _33662_/Q _26518_/S VGND VGND VPWR VPWR _26517_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29304_ _29304_/A VGND VGND VPWR VPWR _34919_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23728_ _22917_/X _32410_/Q _23742_/S VGND VGND VPWR VPWR _23729_/A sky130_fd_sc_hd__mux2_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27496_ _27496_/A VGND VGND VPWR VPWR _34094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29235_ _34889_/Q _29234_/X _29235_/S VGND VGND VPWR VPWR _29236_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26447_ _25038_/X _33629_/Q _26455_/S VGND VGND VPWR VPWR _26448_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23659_ _32379_/Q _23286_/X _23667_/S VGND VGND VPWR VPWR _23660_/A sky130_fd_sc_hd__mux2_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16200_ _34513_/Q _32401_/Q _34385_/Q _34321_/Q _16166_/X _16167_/X VGND VGND VPWR
+ VPWR _16200_/X sky130_fd_sc_hd__mux4_1
XFILLER_161_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17180_ _35757_/Q _35117_/Q _34477_/Q _33837_/Q _17140_/X _17141_/X VGND VGND VPWR
+ VPWR _17180_/X sky130_fd_sc_hd__mux4_1
X_29166_ input31/X VGND VGND VPWR VPWR _29166_/X sky130_fd_sc_hd__clkbuf_4
X_26378_ _26378_/A VGND VGND VPWR VPWR _33596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16131_ _35023_/Q _34959_/Q _34895_/Q _34831_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _16131_/X sky130_fd_sc_hd__mux4_1
XFILLER_183_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28117_ _26841_/X _34388_/Q _28123_/S VGND VGND VPWR VPWR _28118_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25329_ _24995_/X _33103_/Q _25345_/S VGND VGND VPWR VPWR _25330_/A sky130_fd_sc_hd__mux2_1
X_29097_ _29097_/A VGND VGND VPWR VPWR _34844_/D sky130_fd_sc_hd__clkbuf_1
X_28048_ _28048_/A VGND VGND VPWR VPWR _34355_/D sky130_fd_sc_hd__clkbuf_1
X_16062_ _17978_/A VGND VGND VPWR VPWR _17931_/A sky130_fd_sc_hd__buf_12
XFILLER_6_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30010_ _35254_/Q _29175_/X _30028_/S VGND VGND VPWR VPWR _30011_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19821_ _33527_/Q _33463_/Q _33399_/Q _33335_/Q _19776_/X _19777_/X VGND VGND VPWR
+ VPWR _19821_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29999_ _35249_/Q _29160_/X _30007_/S VGND VGND VPWR VPWR _30000_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19752_ _19708_/X _19750_/X _19751_/X _19714_/X VGND VGND VPWR VPWR _19752_/X sky130_fd_sc_hd__a22o_1
X_16964_ _16641_/X _16962_/X _16963_/X _16644_/X VGND VGND VPWR VPWR _16964_/X sky130_fd_sc_hd__a22o_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18703_ _18593_/X _18701_/X _18702_/X _18596_/X VGND VGND VPWR VPWR _18703_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31961_ _35036_/CLK _31961_/D VGND VGND VPWR VPWR _31961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19683_ _19363_/X _19681_/X _19682_/X _19367_/X VGND VGND VPWR VPWR _19683_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16895_ _35749_/Q _35109_/Q _34469_/Q _33829_/Q _16787_/X _16788_/X VGND VGND VPWR
+ VPWR _16895_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33700_ _33702_/CLK _33700_/D VGND VGND VPWR VPWR _33700_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_481_CLK clkbuf_6_3__f_CLK/X VGND VGND VPWR VPWR _35931_/CLK sky130_fd_sc_hd__clkbuf_16
X_18634_ _35285_/Q _35221_/Q _35157_/Q _32277_/Q _18600_/X _18601_/X VGND VGND VPWR
+ VPWR _18634_/X sky130_fd_sc_hd__mux4_1
X_30912_ _30912_/A VGND VGND VPWR VPWR _35681_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_209_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34680_ _35318_/CLK _34680_/D VGND VGND VPWR VPWR _34680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31892_ _23256_/X _36146_/Q _31898_/S VGND VGND VPWR VPWR _31893_/A sky130_fd_sc_hd__mux2_1
XTAP_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33631_ _34080_/CLK _33631_/D VGND VGND VPWR VPWR _33631_/Q sky130_fd_sc_hd__dfxtp_1
X_30843_ _30843_/A VGND VGND VPWR VPWR _35648_/D sky130_fd_sc_hd__clkbuf_1
X_18565_ _18374_/X _18563_/X _18564_/X _18384_/X VGND VGND VPWR VPWR _18565_/X sky130_fd_sc_hd__a22o_1
XTAP_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_233_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _34816_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_205_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17516_ _17516_/A _17516_/B _17516_/C _17516_/D VGND VGND VPWR VPWR _17517_/A sky130_fd_sc_hd__or4_1
X_33562_ _33692_/CLK _33562_/D VGND VGND VPWR VPWR _33562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18496_ _18490_/X _18495_/X _18371_/X VGND VGND VPWR VPWR _18504_/C sky130_fd_sc_hd__o21ba_1
X_30774_ _23142_/X _35616_/Q _30776_/S VGND VGND VPWR VPWR _30775_/A sky130_fd_sc_hd__mux2_1
XANTENNA_580 _20153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_591 _19457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35301_ _36005_/CLK _35301_/D VGND VGND VPWR VPWR _35301_/Q sky130_fd_sc_hd__dfxtp_1
X_32513_ _36033_/CLK _32513_/D VGND VGND VPWR VPWR _32513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17447_ _34037_/Q _33973_/Q _33909_/Q _32245_/Q _17373_/X _17374_/X VGND VGND VPWR
+ VPWR _17447_/X sky130_fd_sc_hd__mux4_1
X_33493_ _34006_/CLK _33493_/D VGND VGND VPWR VPWR _33493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35232_ _35294_/CLK _35232_/D VGND VGND VPWR VPWR _35232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32444_ _35580_/CLK _32444_/D VGND VGND VPWR VPWR _32444_/Q sky130_fd_sc_hd__dfxtp_1
X_17378_ _32755_/Q _32691_/Q _32627_/Q _36083_/Q _17272_/X _17056_/X VGND VGND VPWR
+ VPWR _17378_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19117_ _18796_/X _19115_/X _19116_/X _18799_/X VGND VGND VPWR VPWR _19117_/X sky130_fd_sc_hd__a22o_1
XFILLER_203_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16329_ _35541_/Q _35477_/Q _35413_/Q _35349_/Q _16191_/X _16192_/X VGND VGND VPWR
+ VPWR _16329_/X sky130_fd_sc_hd__mux4_1
X_35163_ _36201_/CLK _35163_/D VGND VGND VPWR VPWR _35163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32375_ _36023_/CLK _32375_/D VGND VGND VPWR VPWR _32375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34114_ _34243_/CLK _34114_/D VGND VGND VPWR VPWR _34114_/Q sky130_fd_sc_hd__dfxtp_1
X_31326_ _31326_/A VGND VGND VPWR VPWR _35877_/D sky130_fd_sc_hd__clkbuf_1
X_19048_ _32993_/Q _32929_/Q _32865_/Q _32801_/Q _18936_/X _18937_/X VGND VGND VPWR
+ VPWR _19048_/X sky130_fd_sc_hd__mux4_1
X_35094_ _35925_/CLK _35094_/D VGND VGND VPWR VPWR _35094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput201 _36226_/Q VGND VGND VPWR VPWR D2[52] sky130_fd_sc_hd__buf_2
Xoutput212 _36236_/Q VGND VGND VPWR VPWR D2[62] sky130_fd_sc_hd__buf_2
X_31257_ _35845_/Q input51/X _31265_/S VGND VGND VPWR VPWR _31258_/A sky130_fd_sc_hd__mux2_1
X_34045_ _36157_/CLK _34045_/D VGND VGND VPWR VPWR _34045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput223 _32092_/Q VGND VGND VPWR VPWR D3[14] sky130_fd_sc_hd__buf_2
XFILLER_86_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput234 _32102_/Q VGND VGND VPWR VPWR D3[24] sky130_fd_sc_hd__buf_2
Xoutput245 _32112_/Q VGND VGND VPWR VPWR D3[34] sky130_fd_sc_hd__buf_2
Xoutput256 _32122_/Q VGND VGND VPWR VPWR D3[44] sky130_fd_sc_hd__buf_2
X_21010_ _20687_/X _21008_/X _21009_/X _20697_/X VGND VGND VPWR VPWR _21010_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput267 _32132_/Q VGND VGND VPWR VPWR D3[54] sky130_fd_sc_hd__buf_2
X_30208_ _35348_/Q _29070_/X _30214_/S VGND VGND VPWR VPWR _30209_/A sky130_fd_sc_hd__mux2_1
X_31188_ _35812_/Q input15/X _31202_/S VGND VGND VPWR VPWR _31189_/A sky130_fd_sc_hd__mux2_1
Xoutput278 _32084_/Q VGND VGND VPWR VPWR D3[6] sky130_fd_sc_hd__buf_2
XFILLER_59_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30139_ _30139_/A VGND VGND VPWR VPWR _35315_/D sky130_fd_sc_hd__clkbuf_1
X_35996_ _36129_/CLK _35996_/D VGND VGND VPWR VPWR _35996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34947_ _34947_/CLK _34947_/D VGND VGND VPWR VPWR _34947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22961_ _22960_/X _32040_/Q _22970_/S VGND VGND VPWR VPWR _22962_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24700_ _24700_/A VGND VGND VPWR VPWR _32837_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_472_CLK clkbuf_6_8__f_CLK/X VGND VGND VPWR VPWR _35552_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_74_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21912_ _21908_/X _21911_/X _21736_/X _21737_/X VGND VGND VPWR VPWR _21929_/B sky130_fd_sc_hd__o211a_1
X_25680_ _25680_/A VGND VGND VPWR VPWR _33266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22892_ input45/X VGND VGND VPWR VPWR _22892_/X sky130_fd_sc_hd__clkbuf_4
X_34878_ _35326_/CLK _34878_/D VGND VGND VPWR VPWR _34878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24631_ _24631_/A VGND VGND VPWR VPWR _32804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33829_ _35941_/CLK _33829_/D VGND VGND VPWR VPWR _33829_/Q sky130_fd_sc_hd__dfxtp_1
X_21843_ _32495_/Q _32367_/Q _32047_/Q _36015_/Q _21523_/X _21664_/X VGND VGND VPWR
+ VPWR _21843_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_224_CLK clkbuf_6_54__f_CLK/X VGND VGND VPWR VPWR _35777_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27350_ _27350_/A VGND VGND VPWR VPWR _34025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1023 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24562_ _24562_/A VGND VGND VPWR VPWR _32773_/D sky130_fd_sc_hd__clkbuf_1
X_21774_ _21655_/X _21772_/X _21773_/X _21661_/X VGND VGND VPWR VPWR _21774_/X sky130_fd_sc_hd__a22o_1
XFILLER_212_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26301_ _26412_/S VGND VGND VPWR VPWR _26320_/S sky130_fd_sc_hd__buf_4
XFILLER_23_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23513_ _23513_/A VGND VGND VPWR VPWR _32310_/D sky130_fd_sc_hd__clkbuf_1
X_27281_ _27005_/X _33993_/Q _27281_/S VGND VGND VPWR VPWR _27282_/A sky130_fd_sc_hd__mux2_1
X_20725_ _20656_/X _20723_/X _20724_/X _20668_/X VGND VGND VPWR VPWR _20725_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24493_ _24493_/A VGND VGND VPWR VPWR _32740_/D sky130_fd_sc_hd__clkbuf_1
X_29020_ _34816_/Q _24400_/X _29038_/S VGND VGND VPWR VPWR _29021_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26232_ _25119_/X _33527_/Q _26248_/S VGND VGND VPWR VPWR _26233_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23444_ _22904_/X _32278_/Q _23446_/S VGND VGND VPWR VPWR _23445_/A sky130_fd_sc_hd__mux2_1
X_20656_ _22460_/A VGND VGND VPWR VPWR _20656_/X sky130_fd_sc_hd__buf_4
XFILLER_17_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26163_ _26163_/A VGND VGND VPWR VPWR _33494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23375_ _23375_/A VGND VGND VPWR VPWR _32246_/D sky130_fd_sc_hd__clkbuf_1
X_20587_ _22506_/A VGND VGND VPWR VPWR _20587_/X sky130_fd_sc_hd__buf_4
XFILLER_221_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25114_ _25114_/A VGND VGND VPWR VPWR _33013_/D sky130_fd_sc_hd__clkbuf_1
X_22326_ _22446_/A VGND VGND VPWR VPWR _22326_/X sky130_fd_sc_hd__buf_4
X_26094_ _26142_/S VGND VGND VPWR VPWR _26113_/S sky130_fd_sc_hd__buf_4
XFILLER_125_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1008 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29922_ _35213_/Q _29246_/X _29922_/S VGND VGND VPWR VPWR _29923_/A sky130_fd_sc_hd__mux2_1
X_25045_ _25044_/X _32991_/Q _25051_/S VGND VGND VPWR VPWR _25046_/A sky130_fd_sc_hd__mux2_1
X_22257_ _22155_/X _22255_/X _22256_/X _22158_/X VGND VGND VPWR VPWR _22257_/X sky130_fd_sc_hd__a22o_1
XFILLER_219_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_1163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21208_ _22396_/A VGND VGND VPWR VPWR _21208_/X sky130_fd_sc_hd__clkbuf_4
X_29853_ _29922_/S VGND VGND VPWR VPWR _29872_/S sky130_fd_sc_hd__buf_4
X_22188_ _22148_/X _22186_/X _22187_/X _22153_/X VGND VGND VPWR VPWR _22188_/X sky130_fd_sc_hd__a22o_1
XFILLER_152_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28804_ _28804_/A VGND VGND VPWR VPWR _34713_/D sky130_fd_sc_hd__clkbuf_1
X_21139_ _20957_/X _21137_/X _21138_/X _20961_/X VGND VGND VPWR VPWR _21139_/X sky130_fd_sc_hd__a22o_1
X_29784_ _29784_/A VGND VGND VPWR VPWR _35147_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26996_ input52/X VGND VGND VPWR VPWR _26996_/X sky130_fd_sc_hd__buf_4
XFILLER_48_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28735_ _26956_/X _34681_/Q _28747_/S VGND VGND VPWR VPWR _28736_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25947_ _25097_/X _33392_/Q _25957_/S VGND VGND VPWR VPWR _25948_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_463_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _35879_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16680_ _35743_/Q _35103_/Q _34463_/Q _33823_/Q _16434_/X _16435_/X VGND VGND VPWR
+ VPWR _16680_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25878_ _24995_/X _33359_/Q _25894_/S VGND VGND VPWR VPWR _25879_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28666_ _26853_/X _34648_/Q _28684_/S VGND VGND VPWR VPWR _28667_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24829_ _24829_/A VGND VGND VPWR VPWR _32897_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27617_ _34151_/Q _24323_/X _27625_/S VGND VGND VPWR VPWR _27618_/A sky130_fd_sc_hd__mux2_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28597_ _28597_/A VGND VGND VPWR VPWR _34615_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_215_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _35079_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18350_ _20062_/A VGND VGND VPWR VPWR _20295_/A sky130_fd_sc_hd__buf_12
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27548_ _27548_/A VGND VGND VPWR VPWR _34119_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _17195_/X _17299_/X _17300_/X _17200_/X VGND VGND VPWR VPWR _17301_/X sky130_fd_sc_hd__a22o_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18281_ input78/X VGND VGND VPWR VPWR _18359_/A sky130_fd_sc_hd__buf_6
XFILLER_163_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27479_ _27479_/A VGND VGND VPWR VPWR _34086_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29218_ _29218_/A VGND VGND VPWR VPWR _34883_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17232_ _17232_/A VGND VGND VPWR VPWR _31982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30490_ _23121_/X _35481_/Q _30506_/S VGND VGND VPWR VPWR _30491_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17163_ _17163_/A _17163_/B _17163_/C _17163_/D VGND VGND VPWR VPWR _17164_/A sky130_fd_sc_hd__or4_4
X_29149_ _34861_/Q _29148_/X _29173_/S VGND VGND VPWR VPWR _29150_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16114_ _33231_/Q _36111_/Q _33103_/Q _33039_/Q _16020_/X _16021_/X VGND VGND VPWR
+ VPWR _16114_/X sky130_fd_sc_hd__mux4_1
X_32160_ _34271_/CLK _32160_/D VGND VGND VPWR VPWR _32160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17094_ _34027_/Q _33963_/Q _33899_/Q _32235_/Q _17020_/X _17021_/X VGND VGND VPWR
+ VPWR _17094_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31111_ _31138_/S VGND VGND VPWR VPWR _31130_/S sky130_fd_sc_hd__buf_4
XFILLER_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16045_ _17795_/A VGND VGND VPWR VPWR _16045_/X sky130_fd_sc_hd__buf_8
XFILLER_157_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32091_ _35040_/CLK _32091_/D VGND VGND VPWR VPWR _32091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31042_ _35743_/Q _29104_/X _31046_/S VGND VGND VPWR VPWR _31043_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19804_ _35318_/Q _35254_/Q _35190_/Q _32310_/Q _19659_/X _19660_/X VGND VGND VPWR
+ VPWR _19804_/X sky130_fd_sc_hd__mux4_1
X_35850_ _35852_/CLK _35850_/D VGND VGND VPWR VPWR _35850_/Q sky130_fd_sc_hd__dfxtp_1
X_17996_ _34820_/Q _34756_/Q _34692_/Q _34628_/Q _17994_/X _17995_/X VGND VGND VPWR
+ VPWR _17996_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34801_ _35061_/CLK _34801_/D VGND VGND VPWR VPWR _34801_/Q sky130_fd_sc_hd__dfxtp_1
X_19735_ _34548_/Q _32436_/Q _34420_/Q _34356_/Q _19525_/X _19526_/X VGND VGND VPWR
+ VPWR _19735_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35781_ _35781_/CLK _35781_/D VGND VGND VPWR VPWR _35781_/Q sky130_fd_sc_hd__dfxtp_1
X_16947_ _34279_/Q _34215_/Q _34151_/Q _34087_/Q _16736_/X _16737_/X VGND VGND VPWR
+ VPWR _16947_/X sky130_fd_sc_hd__mux4_1
XFILLER_42_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32993_ _36065_/CLK _32993_/D VGND VGND VPWR VPWR _32993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_454_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _36005_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_226_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34732_ _35242_/CLK _34732_/D VGND VGND VPWR VPWR _34732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31944_ _23339_/X _36171_/Q _31948_/S VGND VGND VPWR VPWR _31945_/A sky130_fd_sc_hd__mux2_1
X_19666_ _19662_/X _19665_/X _19461_/X VGND VGND VPWR VPWR _19667_/D sky130_fd_sc_hd__o21ba_1
X_16878_ _16878_/A _16878_/B _16878_/C _16878_/D VGND VGND VPWR VPWR _16879_/A sky130_fd_sc_hd__or4_4
XFILLER_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18617_ _18443_/X _18613_/X _18616_/X _18446_/X VGND VGND VPWR VPWR _18617_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34663_ _36005_/CLK _34663_/D VGND VGND VPWR VPWR _34663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19597_ _19597_/A _19597_/B _19597_/C _19597_/D VGND VGND VPWR VPWR _19598_/A sky130_fd_sc_hd__or4_1
XFILLER_52_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31875_ _23231_/X _36138_/Q _31877_/S VGND VGND VPWR VPWR _31876_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_206_CLK clkbuf_6_52__f_CLK/X VGND VGND VPWR VPWR _36168_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_225_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33614_ _34256_/CLK _33614_/D VGND VGND VPWR VPWR _33614_/Q sky130_fd_sc_hd__dfxtp_1
X_18548_ _33235_/Q _36115_/Q _33107_/Q _33043_/Q _18320_/X _18321_/X VGND VGND VPWR
+ VPWR _18548_/X sky130_fd_sc_hd__mux4_1
X_30826_ _30826_/A VGND VGND VPWR VPWR _35640_/D sky130_fd_sc_hd__clkbuf_1
X_34594_ _35928_/CLK _34594_/D VGND VGND VPWR VPWR _34594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33545_ _33545_/CLK _33545_/D VGND VGND VPWR VPWR _33545_/Q sky130_fd_sc_hd__dfxtp_1
X_18479_ _18443_/X _18477_/X _18478_/X _18446_/X VGND VGND VPWR VPWR _18479_/X sky130_fd_sc_hd__a22o_1
X_30757_ _30868_/S VGND VGND VPWR VPWR _30776_/S sky130_fd_sc_hd__buf_4
XFILLER_33_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20510_ _35083_/Q _35019_/Q _34955_/Q _34891_/Q _18379_/X _18381_/X VGND VGND VPWR
+ VPWR _20510_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33476_ _33545_/CLK _33476_/D VGND VGND VPWR VPWR _33476_/Q sky130_fd_sc_hd__dfxtp_1
X_21490_ _32485_/Q _32357_/Q _32037_/Q _36005_/Q _21170_/X _21311_/X VGND VGND VPWR
+ VPWR _21490_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30688_ _35575_/Q _29179_/X _30704_/S VGND VGND VPWR VPWR _30689_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35215_ _35215_/CLK _35215_/D VGND VGND VPWR VPWR _35215_/Q sky130_fd_sc_hd__dfxtp_1
X_20441_ _18277_/X _20439_/X _20440_/X _18287_/X VGND VGND VPWR VPWR _20441_/X sky130_fd_sc_hd__a22o_1
X_32427_ _35179_/CLK _32427_/D VGND VGND VPWR VPWR _32427_/Q sky130_fd_sc_hd__dfxtp_1
X_36195_ _36196_/CLK _36195_/D VGND VGND VPWR VPWR _36195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35146_ _35788_/CLK _35146_/D VGND VGND VPWR VPWR _35146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23160_ _23346_/S VGND VGND VPWR VPWR _23182_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_118_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20372_ _32775_/Q _32711_/Q _32647_/Q _36103_/Q _20278_/X _20062_/X VGND VGND VPWR
+ VPWR _20372_/X sky130_fd_sc_hd__mux4_1
XFILLER_134_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32358_ _36005_/CLK _32358_/D VGND VGND VPWR VPWR _32358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22111_ _35062_/Q _34998_/Q _34934_/Q _34870_/Q _22109_/X _22110_/X VGND VGND VPWR
+ VPWR _22111_/X sky130_fd_sc_hd__mux4_1
XTAP_7109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31309_ _31309_/A VGND VGND VPWR VPWR _35869_/D sky130_fd_sc_hd__clkbuf_1
X_35077_ _35781_/CLK _35077_/D VGND VGND VPWR VPWR _35077_/Q sky130_fd_sc_hd__dfxtp_1
X_23091_ _32143_/Q _23090_/X _23115_/S VGND VGND VPWR VPWR _23092_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32289_ _35296_/CLK _32289_/D VGND VGND VPWR VPWR _32289_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22042_ _22556_/A VGND VGND VPWR VPWR _22042_/X sky130_fd_sc_hd__buf_4
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34028_ _35958_/CLK _34028_/D VGND VGND VPWR VPWR _34028_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26850_ input64/X VGND VGND VPWR VPWR _26850_/X sky130_fd_sc_hd__buf_4
XTAP_5729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25801_ _25081_/X _33323_/Q _25801_/S VGND VGND VPWR VPWR _25802_/A sky130_fd_sc_hd__mux2_1
X_26781_ _26781_/A VGND VGND VPWR VPWR _33786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35979_ _35979_/CLK _35979_/D VGND VGND VPWR VPWR _35979_/Q sky130_fd_sc_hd__dfxtp_1
X_23993_ _22907_/X _32535_/Q _23993_/S VGND VGND VPWR VPWR _23994_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_445_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _36132_/CLK sky130_fd_sc_hd__clkbuf_16
X_25732_ _25732_/A VGND VGND VPWR VPWR _33291_/D sky130_fd_sc_hd__clkbuf_1
X_28520_ _26838_/X _34579_/Q _28528_/S VGND VGND VPWR VPWR _28521_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22944_ _22944_/A VGND VGND VPWR VPWR _32034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_1356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28451_ _28451_/A VGND VGND VPWR VPWR _34546_/D sky130_fd_sc_hd__clkbuf_1
X_25663_ _25663_/A VGND VGND VPWR VPWR _33258_/D sky130_fd_sc_hd__clkbuf_1
X_22875_ input1/X VGND VGND VPWR VPWR _22875_/X sky130_fd_sc_hd__buf_4
XFILLER_216_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27402_ _34050_/Q _24407_/X _27416_/S VGND VGND VPWR VPWR _27403_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24614_ _24614_/A VGND VGND VPWR VPWR _32796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28382_ _28382_/A VGND VGND VPWR VPWR _34513_/D sky130_fd_sc_hd__clkbuf_1
X_21826_ _22532_/A VGND VGND VPWR VPWR _21826_/X sky130_fd_sc_hd__buf_4
X_25594_ _25594_/A VGND VGND VPWR VPWR _33227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27333_ _27333_/A VGND VGND VPWR VPWR _34017_/D sky130_fd_sc_hd__clkbuf_1
X_24545_ _24545_/A VGND VGND VPWR VPWR _32765_/D sky130_fd_sc_hd__clkbuf_1
X_21757_ _21757_/A VGND VGND VPWR VPWR _21757_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_169_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20708_ _22446_/A VGND VGND VPWR VPWR _20708_/X sky130_fd_sc_hd__buf_6
X_27264_ _27264_/A VGND VGND VPWR VPWR _33984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24476_ _24476_/A VGND VGND VPWR VPWR _32732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21688_ _33771_/Q _33707_/Q _33643_/Q _33579_/Q _21443_/X _21444_/X VGND VGND VPWR
+ VPWR _21688_/X sky130_fd_sc_hd__mux4_1
XFILLER_8_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26215_ _25094_/X _33519_/Q _26227_/S VGND VGND VPWR VPWR _26216_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29003_ _34808_/Q _24376_/X _29017_/S VGND VGND VPWR VPWR _29004_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23427_ _23559_/S VGND VGND VPWR VPWR _23446_/S sky130_fd_sc_hd__buf_6
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20639_ input75/X VGND VGND VPWR VPWR _22442_/A sky130_fd_sc_hd__buf_12
X_27195_ _26878_/X _33952_/Q _27197_/S VGND VGND VPWR VPWR _27196_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26146_ _24989_/X _33486_/Q _26164_/S VGND VGND VPWR VPWR _26147_/A sky130_fd_sc_hd__mux2_1
X_23358_ _23358_/A VGND VGND VPWR VPWR _32238_/D sky130_fd_sc_hd__clkbuf_1
X_22309_ _22305_/X _22306_/X _22307_/X _22308_/X VGND VGND VPWR VPWR _22309_/X sky130_fd_sc_hd__a22o_1
XFILLER_153_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26077_ _26077_/A VGND VGND VPWR VPWR _33453_/D sky130_fd_sc_hd__clkbuf_1
X_23289_ input41/X VGND VGND VPWR VPWR _23289_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_124_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29905_ _29905_/A VGND VGND VPWR VPWR _35204_/D sky130_fd_sc_hd__clkbuf_1
X_25028_ _25028_/A VGND VGND VPWR VPWR _32985_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17850_ _35584_/Q _35520_/Q _35456_/Q _35392_/Q _17603_/X _17604_/X VGND VGND VPWR
+ VPWR _17850_/X sky130_fd_sc_hd__mux4_1
X_29836_ _29836_/A VGND VGND VPWR VPWR _35171_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16801_ _17154_/A VGND VGND VPWR VPWR _16801_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29767_ _35139_/Q _29216_/X _29779_/S VGND VGND VPWR VPWR _29768_/A sky130_fd_sc_hd__mux2_1
X_17781_ _17932_/A VGND VGND VPWR VPWR _17781_/X sky130_fd_sc_hd__buf_4
X_26979_ _26977_/X _33856_/Q _27006_/S VGND VGND VPWR VPWR _26980_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_436_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _34153_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_208_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19520_ _19299_/X _19518_/X _19519_/X _19302_/X VGND VGND VPWR VPWR _19520_/X sky130_fd_sc_hd__a22o_1
XFILLER_8_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16732_ _16728_/X _16731_/X _16455_/X VGND VGND VPWR VPWR _16733_/D sky130_fd_sc_hd__o21ba_1
X_28718_ _26931_/X _34673_/Q _28726_/S VGND VGND VPWR VPWR _28719_/A sky130_fd_sc_hd__mux2_1
X_29698_ _35106_/Q _29113_/X _29716_/S VGND VGND VPWR VPWR _29699_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19451_ _35308_/Q _35244_/Q _35180_/Q _32300_/Q _19306_/X _19307_/X VGND VGND VPWR
+ VPWR _19451_/X sky130_fd_sc_hd__mux4_1
X_28649_ _26829_/X _34640_/Q _28663_/S VGND VGND VPWR VPWR _28650_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16663_ _33759_/Q _33695_/Q _33631_/Q _33567_/Q _16490_/X _16491_/X VGND VGND VPWR
+ VPWR _16663_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18402_ _18402_/A _18402_/B _18402_/C _18402_/D VGND VGND VPWR VPWR _18403_/A sky130_fd_sc_hd__or4_4
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31660_ _36036_/Q input50/X _31670_/S VGND VGND VPWR VPWR _31661_/A sky130_fd_sc_hd__mux2_1
X_19382_ _34538_/Q _32426_/Q _34410_/Q _34346_/Q _19172_/X _19173_/X VGND VGND VPWR
+ VPWR _19382_/X sky130_fd_sc_hd__mux4_1
X_16594_ _34269_/Q _34205_/Q _34141_/Q _34077_/Q _16383_/X _16384_/X VGND VGND VPWR
+ VPWR _16594_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30611_ _30611_/A VGND VGND VPWR VPWR _35538_/D sky130_fd_sc_hd__clkbuf_1
X_18333_ _20129_/A VGND VGND VPWR VPWR _18333_/X sky130_fd_sc_hd__buf_4
XFILLER_61_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31591_ _36003_/Q input14/X _31607_/S VGND VGND VPWR VPWR _31592_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33330_ _33775_/CLK _33330_/D VGND VGND VPWR VPWR _33330_/Q sky130_fd_sc_hd__dfxtp_1
X_18264_ _15997_/X _18262_/X _18263_/X _16003_/X VGND VGND VPWR VPWR _18264_/X sky130_fd_sc_hd__a22o_1
X_30542_ _23256_/X _35506_/Q _30548_/S VGND VGND VPWR VPWR _30543_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17215_ _35822_/Q _32199_/Q _35694_/Q _35630_/Q _16960_/X _16961_/X VGND VGND VPWR
+ VPWR _17215_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33261_ _36141_/CLK _33261_/D VGND VGND VPWR VPWR _33261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18195_ _32523_/Q _32395_/Q _32075_/Q _36043_/Q _17982_/X _17007_/A VGND VGND VPWR
+ VPWR _18195_/X sky130_fd_sc_hd__mux4_1
X_30473_ _23096_/X _35473_/Q _30485_/S VGND VGND VPWR VPWR _30474_/A sky130_fd_sc_hd__mux2_1
X_35000_ _35578_/CLK _35000_/D VGND VGND VPWR VPWR _35000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32212_ _35834_/CLK _32212_/D VGND VGND VPWR VPWR _32212_/Q sky130_fd_sc_hd__dfxtp_1
X_17146_ _16999_/X _17144_/X _17145_/X _17002_/X VGND VGND VPWR VPWR _17146_/X sky130_fd_sc_hd__a22o_1
X_33192_ _35944_/CLK _33192_/D VGND VGND VPWR VPWR _33192_/Q sky130_fd_sc_hd__dfxtp_1
X_32143_ _35664_/CLK _32143_/D VGND VGND VPWR VPWR _32143_/Q sky130_fd_sc_hd__dfxtp_1
X_17077_ _16999_/X _17073_/X _17076_/X _17002_/X VGND VGND VPWR VPWR _17077_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16028_ _17982_/A VGND VGND VPWR VPWR _16028_/X sky130_fd_sc_hd__buf_6
XFILLER_237_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32074_ _36170_/CLK _32074_/D VGND VGND VPWR VPWR _32074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35902_ _35903_/CLK _35902_/D VGND VGND VPWR VPWR _35902_/Q sky130_fd_sc_hd__dfxtp_1
X_31025_ _35735_/Q _29079_/X _31025_/S VGND VGND VPWR VPWR _31026_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35833_ _35833_/CLK _35833_/D VGND VGND VPWR VPWR _35833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17979_ _32772_/Q _32708_/Q _32644_/Q _36100_/Q _17978_/X _17762_/X VGND VGND VPWR
+ VPWR _17979_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_427_CLK clkbuf_6_36__f_CLK/X VGND VGND VPWR VPWR _36137_/CLK sky130_fd_sc_hd__clkbuf_16
X_19718_ _32500_/Q _32372_/Q _32052_/Q _36020_/Q _19576_/X _19717_/X VGND VGND VPWR
+ VPWR _19718_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35764_ _35828_/CLK _35764_/D VGND VGND VPWR VPWR _35764_/Q sky130_fd_sc_hd__dfxtp_1
X_20990_ _20986_/X _20989_/X _20611_/X VGND VGND VPWR VPWR _21012_/A sky130_fd_sc_hd__o21ba_1
X_32976_ _36049_/CLK _32976_/D VGND VGND VPWR VPWR _32976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34715_ _34779_/CLK _34715_/D VGND VGND VPWR VPWR _34715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31927_ _31927_/A VGND VGND VPWR VPWR _36162_/D sky130_fd_sc_hd__clkbuf_1
X_19649_ _35762_/Q _35122_/Q _34482_/Q _33842_/Q _19440_/X _19441_/X VGND VGND VPWR
+ VPWR _19649_/X sky130_fd_sc_hd__mux4_1
X_35695_ _35822_/CLK _35695_/D VGND VGND VPWR VPWR _35695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22660_ _35078_/Q _35014_/Q _34950_/Q _34886_/Q _22462_/X _22463_/X VGND VGND VPWR
+ VPWR _22660_/X sky130_fd_sc_hd__mux4_1
XFILLER_198_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34646_ _35286_/CLK _34646_/D VGND VGND VPWR VPWR _34646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31858_ _31948_/S VGND VGND VPWR VPWR _31877_/S sky130_fd_sc_hd__buf_4
XFILLER_240_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21611_ _35048_/Q _34984_/Q _34920_/Q _34856_/Q _21403_/X _21404_/X VGND VGND VPWR
+ VPWR _21611_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30809_ _30809_/A VGND VGND VPWR VPWR _35632_/D sky130_fd_sc_hd__clkbuf_1
X_34577_ _36216_/CLK _34577_/D VGND VGND VPWR VPWR _34577_/Q sky130_fd_sc_hd__dfxtp_1
X_22591_ _33220_/Q _32580_/Q _35972_/Q _35908_/Q _22380_/X _22381_/X VGND VGND VPWR
+ VPWR _22591_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31789_ _36097_/Q input47/X _31805_/S VGND VGND VPWR VPWR _31790_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_1075 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24330_ _32681_/Q _24329_/X _24336_/S VGND VGND VPWR VPWR _24331_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33528_ _34297_/CLK _33528_/D VGND VGND VPWR VPWR _33528_/Q sky130_fd_sc_hd__dfxtp_1
X_21542_ _21401_/X _21540_/X _21541_/X _21406_/X VGND VGND VPWR VPWR _21542_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24261_ input56/X VGND VGND VPWR VPWR _24261_/X sky130_fd_sc_hd__buf_6
X_21473_ _21473_/A VGND VGND VPWR VPWR _21473_/X sky130_fd_sc_hd__buf_4
X_33459_ _33779_/CLK _33459_/D VGND VGND VPWR VPWR _33459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26000_ _26000_/A VGND VGND VPWR VPWR _33417_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_51__f_CLK clkbuf_5_25_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_51__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_23212_ _23212_/A VGND VGND VPWR VPWR _32187_/D sky130_fd_sc_hd__clkbuf_1
X_20424_ _20424_/A VGND VGND VPWR VPWR _32136_/D sky130_fd_sc_hd__buf_4
XFILLER_193_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36178_ _36185_/CLK _36178_/D VGND VGND VPWR VPWR _36178_/Q sky130_fd_sc_hd__dfxtp_1
X_24192_ _23000_/X _32629_/Q _24192_/S VGND VGND VPWR VPWR _24193_/A sky130_fd_sc_hd__mux2_1
X_35129_ _35771_/CLK _35129_/D VGND VGND VPWR VPWR _35129_/Q sky130_fd_sc_hd__dfxtp_1
X_23143_ _32160_/Q _23142_/X _23146_/S VGND VGND VPWR VPWR _23144_/A sky130_fd_sc_hd__mux2_1
X_20355_ _20351_/X _20354_/X _20153_/X VGND VGND VPWR VPWR _20363_/C sky130_fd_sc_hd__o21ba_1
XFILLER_136_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27951_ _27951_/A VGND VGND VPWR VPWR _34309_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23074_ input60/X VGND VGND VPWR VPWR _23074_/X sky130_fd_sc_hd__buf_2
XFILLER_134_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20286_ _20281_/X _20285_/X _20142_/X _20143_/X VGND VGND VPWR VPWR _20303_/B sky130_fd_sc_hd__o211a_1
XFILLER_153_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26902_ _26902_/A VGND VGND VPWR VPWR _33831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22025_ _21947_/X _22023_/X _22024_/X _21950_/X VGND VGND VPWR VPWR _22025_/X sky130_fd_sc_hd__a22o_1
XFILLER_248_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27882_ _27882_/A VGND VGND VPWR VPWR _34276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29621_ _35070_/Q _29200_/X _29623_/S VGND VGND VPWR VPWR _29622_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26833_ _26832_/X _33809_/Q _26851_/S VGND VGND VPWR VPWR _26834_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_418_CLK clkbuf_6_35__f_CLK/X VGND VGND VPWR VPWR _35061_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29552_ _35037_/Q _29098_/X _29560_/S VGND VGND VPWR VPWR _29553_/A sky130_fd_sc_hd__mux2_1
X_23976_ _23976_/A VGND VGND VPWR VPWR _32526_/D sky130_fd_sc_hd__clkbuf_1
X_26764_ _26764_/A VGND VGND VPWR VPWR _33778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28503_ _28503_/A VGND VGND VPWR VPWR _34571_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25715_ _33283_/Q _24410_/X _25727_/S VGND VGND VPWR VPWR _25716_/A sky130_fd_sc_hd__mux2_1
X_22927_ _22926_/X _32029_/Q _22939_/S VGND VGND VPWR VPWR _22928_/A sky130_fd_sc_hd__mux2_1
X_26695_ _26695_/A VGND VGND VPWR VPWR _33745_/D sky130_fd_sc_hd__clkbuf_1
X_29483_ _29483_/A VGND VGND VPWR VPWR _35004_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28434_ _28434_/A VGND VGND VPWR VPWR _34538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22858_ _22854_/X _22857_/X _22442_/A _22443_/A VGND VGND VPWR VPWR _22873_/B sky130_fd_sc_hd__o211a_1
X_25646_ _33250_/Q _24307_/X _25664_/S VGND VGND VPWR VPWR _25647_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21809_ _33262_/Q _36142_/Q _33134_/Q _33070_/Q _21658_/X _21659_/X VGND VGND VPWR
+ VPWR _21809_/X sky130_fd_sc_hd__mux4_1
X_28365_ _34506_/Q _24431_/X _28371_/S VGND VGND VPWR VPWR _28366_/A sky130_fd_sc_hd__mux2_1
X_25577_ _33219_/Q _24410_/X _25589_/S VGND VGND VPWR VPWR _25578_/A sky130_fd_sc_hd__mux2_1
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22789_ _34059_/Q _33995_/Q _33931_/Q _32267_/Q _20658_/X _20660_/X VGND VGND VPWR
+ VPWR _22789_/X sky130_fd_sc_hd__mux4_1
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27316_ _34009_/Q _24280_/X _27332_/S VGND VGND VPWR VPWR _27317_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24528_ _24528_/A VGND VGND VPWR VPWR _32757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28296_ _34473_/Q _24329_/X _28300_/S VGND VGND VPWR VPWR _28297_/A sky130_fd_sc_hd__mux2_1
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24459_ _24459_/A VGND VGND VPWR VPWR _32724_/D sky130_fd_sc_hd__clkbuf_1
X_27247_ _27247_/A VGND VGND VPWR VPWR _33976_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17000_ _35560_/Q _35496_/Q _35432_/Q _35368_/Q _16897_/X _16898_/X VGND VGND VPWR
+ VPWR _17000_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27178_ _27289_/S VGND VGND VPWR VPWR _27197_/S sky130_fd_sc_hd__buf_6
XANTENNA_8 _32114_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26129_ _26129_/A VGND VGND VPWR VPWR _33478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18951_ _18945_/X _18950_/X _18741_/X VGND VGND VPWR VPWR _18961_/C sky130_fd_sc_hd__o21ba_1
XFILLER_10_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17902_ _17902_/A VGND VGND VPWR VPWR _17902_/X sky130_fd_sc_hd__buf_6
X_18882_ _20294_/A VGND VGND VPWR VPWR _18882_/X sky130_fd_sc_hd__buf_6
XTAP_6750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17833_ _17555_/X _17831_/X _17832_/X _17558_/X VGND VGND VPWR VPWR _17833_/X sky130_fd_sc_hd__a22o_1
X_29819_ _29819_/A VGND VGND VPWR VPWR _35163_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_409_CLK clkbuf_6_33__f_CLK/X VGND VGND VPWR VPWR _35050_/CLK sky130_fd_sc_hd__clkbuf_16
X_32830_ _32959_/CLK _32830_/D VGND VGND VPWR VPWR _32830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17764_ _17982_/A VGND VGND VPWR VPWR _17764_/X sky130_fd_sc_hd__buf_4
XFILLER_208_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19503_ _33518_/Q _33454_/Q _33390_/Q _33326_/Q _19423_/X _19424_/X VGND VGND VPWR
+ VPWR _19503_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16715_ _16710_/X _16712_/X _16713_/X _16714_/X VGND VGND VPWR VPWR _16715_/X sky130_fd_sc_hd__a22o_1
X_32761_ _36090_/CLK _32761_/D VGND VGND VPWR VPWR _32761_/Q sky130_fd_sc_hd__dfxtp_1
X_17695_ _17829_/A VGND VGND VPWR VPWR _17695_/X sky130_fd_sc_hd__buf_4
XFILLER_75_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34500_ _35780_/CLK _34500_/D VGND VGND VPWR VPWR _34500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19434_ _33004_/Q _32940_/Q _32876_/Q _32812_/Q _19289_/X _19290_/X VGND VGND VPWR
+ VPWR _19434_/X sky130_fd_sc_hd__mux4_1
X_31712_ _31712_/A VGND VGND VPWR VPWR _36060_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16646_ _17860_/A VGND VGND VPWR VPWR _16646_/X sky130_fd_sc_hd__clkbuf_4
X_35480_ _36001_/CLK _35480_/D VGND VGND VPWR VPWR _35480_/Q sky130_fd_sc_hd__dfxtp_1
X_32692_ _36149_/CLK _32692_/D VGND VGND VPWR VPWR _32692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34431_ _35710_/CLK _34431_/D VGND VGND VPWR VPWR _34431_/Q sky130_fd_sc_hd__dfxtp_1
X_31643_ _36028_/Q input41/X _31649_/S VGND VGND VPWR VPWR _31644_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19365_ _32490_/Q _32362_/Q _32042_/Q _36010_/Q _19223_/X _19364_/X VGND VGND VPWR
+ VPWR _19365_/X sky130_fd_sc_hd__mux4_1
X_16577_ _16288_/X _16575_/X _16576_/X _16291_/X VGND VGND VPWR VPWR _16577_/X sky130_fd_sc_hd__a22o_1
XFILLER_210_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18316_ _20278_/A VGND VGND VPWR VPWR _20162_/A sky130_fd_sc_hd__buf_12
XFILLER_231_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34362_ _34811_/CLK _34362_/D VGND VGND VPWR VPWR _34362_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31574_ _35995_/Q input5/X _31586_/S VGND VGND VPWR VPWR _31575_/A sky130_fd_sc_hd__mux2_1
X_19296_ _35752_/Q _35112_/Q _34472_/Q _33832_/Q _19087_/X _19088_/X VGND VGND VPWR
+ VPWR _19296_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36101_ _36167_/CLK _36101_/D VGND VGND VPWR VPWR _36101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33313_ _34266_/CLK _33313_/D VGND VGND VPWR VPWR _33313_/Q sky130_fd_sc_hd__dfxtp_1
X_18247_ _16014_/X _18245_/X _18246_/X _16023_/X VGND VGND VPWR VPWR _18247_/X sky130_fd_sc_hd__a22o_1
X_30525_ _23231_/X _35498_/Q _30527_/S VGND VGND VPWR VPWR _30526_/A sky130_fd_sc_hd__mux2_1
X_34293_ _34293_/CLK _34293_/D VGND VGND VPWR VPWR _34293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36032_ _36032_/CLK _36032_/D VGND VGND VPWR VPWR _36032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33244_ _33244_/CLK _33244_/D VGND VGND VPWR VPWR _33244_/Q sky130_fd_sc_hd__dfxtp_1
X_18178_ _16044_/X _18176_/X _18177_/X _16054_/X VGND VGND VPWR VPWR _18178_/X sky130_fd_sc_hd__a22o_1
X_30456_ _30456_/A VGND VGND VPWR VPWR _35465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17129_ _17122_/X _17127_/X _17128_/X VGND VGND VPWR VPWR _17163_/A sky130_fd_sc_hd__o21ba_1
X_33175_ _36118_/CLK _33175_/D VGND VGND VPWR VPWR _33175_/Q sky130_fd_sc_hd__dfxtp_1
X_30387_ _30387_/A VGND VGND VPWR VPWR _35432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20140_ _33024_/Q _32960_/Q _32896_/Q _32832_/Q _19995_/X _19996_/X VGND VGND VPWR
+ VPWR _20140_/X sky130_fd_sc_hd__mux4_1
X_32126_ _35562_/CLK _32126_/D VGND VGND VPWR VPWR _32126_/Q sky130_fd_sc_hd__dfxtp_1
X_20071_ _32510_/Q _32382_/Q _32062_/Q _36030_/Q _19929_/X _20070_/X VGND VGND VPWR
+ VPWR _20071_/X sky130_fd_sc_hd__mux4_1
X_32057_ _36025_/CLK _32057_/D VGND VGND VPWR VPWR _32057_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31008_ _31008_/A VGND VGND VPWR VPWR _35726_/D sky130_fd_sc_hd__clkbuf_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_930 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23830_ _23068_/X _32459_/Q _23834_/S VGND VGND VPWR VPWR _23831_/A sky130_fd_sc_hd__mux2_1
XTAP_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35816_ _35818_/CLK _35816_/D VGND VGND VPWR VPWR _35816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35747_ _35748_/CLK _35747_/D VGND VGND VPWR VPWR _35747_/Q sky130_fd_sc_hd__dfxtp_1
X_23761_ _22966_/X _32426_/Q _23763_/S VGND VGND VPWR VPWR _23762_/A sky130_fd_sc_hd__mux2_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_409 _36211_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32959_ _32959_/CLK _32959_/D VGND VGND VPWR VPWR _32959_/Q sky130_fd_sc_hd__dfxtp_1
X_20973_ _34774_/Q _34710_/Q _34646_/Q _34582_/Q _20829_/X _20830_/X VGND VGND VPWR
+ VPWR _20973_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22712_ _35592_/Q _35528_/Q _35464_/Q _35400_/Q _22556_/X _22557_/X VGND VGND VPWR
+ VPWR _22712_/X sky130_fd_sc_hd__mux4_1
XFILLER_26_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25500_ _25500_/A VGND VGND VPWR VPWR _33182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26480_ _26480_/A VGND VGND VPWR VPWR _33644_/D sky130_fd_sc_hd__clkbuf_1
X_23692_ _32395_/Q _23339_/X _23696_/S VGND VGND VPWR VPWR _23693_/A sky130_fd_sc_hd__mux2_1
X_35678_ _35807_/CLK _35678_/D VGND VGND VPWR VPWR _35678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25431_ _25458_/S VGND VGND VPWR VPWR _25450_/S sky130_fd_sc_hd__clkbuf_8
X_34629_ _35333_/CLK _34629_/D VGND VGND VPWR VPWR _34629_/Q sky130_fd_sc_hd__dfxtp_1
X_22643_ _33286_/Q _36166_/Q _33158_/Q _33094_/Q _22364_/X _22365_/X VGND VGND VPWR
+ VPWR _22643_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28150_ _28150_/A VGND VGND VPWR VPWR _34403_/D sky130_fd_sc_hd__clkbuf_1
X_25362_ _25044_/X _33119_/Q _25366_/S VGND VGND VPWR VPWR _25363_/A sky130_fd_sc_hd__mux2_1
X_22574_ _33540_/Q _33476_/Q _33412_/Q _33348_/Q _22429_/X _22430_/X VGND VGND VPWR
+ VPWR _22574_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27101_ _27101_/A VGND VGND VPWR VPWR _33907_/D sky130_fd_sc_hd__clkbuf_1
X_24313_ _24313_/A VGND VGND VPWR VPWR _32675_/D sky130_fd_sc_hd__clkbuf_1
X_28081_ _26987_/X _34371_/Q _28093_/S VGND VGND VPWR VPWR _28082_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21525_ _32998_/Q _32934_/Q _32870_/Q _32806_/Q _21236_/X _21237_/X VGND VGND VPWR
+ VPWR _21525_/X sky130_fd_sc_hd__mux4_1
X_25293_ _25143_/X _33087_/Q _25293_/S VGND VGND VPWR VPWR _25294_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27032_ _27032_/A VGND VGND VPWR VPWR _33874_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24244_ input1/X VGND VGND VPWR VPWR _24244_/X sky130_fd_sc_hd__buf_4
XFILLER_126_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21456_ _33252_/Q _36132_/Q _33124_/Q _33060_/Q _21305_/X _21306_/X VGND VGND VPWR
+ VPWR _21456_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20407_ _19454_/A _20405_/X _20406_/X _19459_/A VGND VGND VPWR VPWR _20407_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24175_ _24175_/A VGND VGND VPWR VPWR _32620_/D sky130_fd_sc_hd__clkbuf_1
X_21387_ _22594_/A VGND VGND VPWR VPWR _21387_/X sky130_fd_sc_hd__buf_6
XFILLER_108_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23126_ _23126_/A VGND VGND VPWR VPWR _32154_/D sky130_fd_sc_hd__clkbuf_1
X_20338_ _33542_/Q _33478_/Q _33414_/Q _33350_/Q _20129_/X _20130_/X VGND VGND VPWR
+ VPWR _20338_/X sky130_fd_sc_hd__mux4_1
X_28983_ _28983_/A VGND VGND VPWR VPWR _34798_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23057_ _23056_/X _32071_/Q _23063_/S VGND VGND VPWR VPWR _23058_/A sky130_fd_sc_hd__mux2_1
X_27934_ _27934_/A VGND VGND VPWR VPWR _34301_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20269_ _20269_/A _20269_/B _20269_/C _20269_/D VGND VGND VPWR VPWR _20270_/A sky130_fd_sc_hd__or4_4
XTAP_5301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22008_ _22501_/A VGND VGND VPWR VPWR _22008_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27865_ _27865_/A VGND VGND VPWR VPWR _34268_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29604_ _29652_/S VGND VGND VPWR VPWR _29623_/S sky130_fd_sc_hd__buf_4
X_26816_ _26816_/A VGND VGND VPWR VPWR _33803_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27796_ _34236_/Q _24388_/X _27802_/S VGND VGND VPWR VPWR _27797_/A sky130_fd_sc_hd__mux2_1
XTAP_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29535_ _35029_/Q _29073_/X _29539_/S VGND VGND VPWR VPWR _29536_/A sky130_fd_sc_hd__mux2_1
XTAP_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26747_ _26747_/A VGND VGND VPWR VPWR _33770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23959_ _23959_/A VGND VGND VPWR VPWR _32519_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1096 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_910 _27018_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_921 _27154_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16500_ _16496_/X _16497_/X _16498_/X _16499_/X VGND VGND VPWR VPWR _16500_/X sky130_fd_sc_hd__a22o_1
XTAP_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17480_ _17202_/X _17478_/X _17479_/X _17205_/X VGND VGND VPWR VPWR _17480_/X sky130_fd_sc_hd__a22o_1
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_932 _29247_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29466_ _29466_/A VGND VGND VPWR VPWR _34996_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26678_ _26678_/A VGND VGND VPWR VPWR _33738_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_943 _29382_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_954 _29787_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_965 _31138_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28417_ _26884_/X _34530_/Q _28435_/S VGND VGND VPWR VPWR _28418_/A sky130_fd_sc_hd__mux2_1
X_16431_ _17843_/A VGND VGND VPWR VPWR _16431_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_976 _31948_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25629_ _33242_/Q _24283_/X _25643_/S VGND VGND VPWR VPWR _25630_/A sky130_fd_sc_hd__mux2_1
X_29397_ _29397_/A VGND VGND VPWR VPWR _34963_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_987 _17796_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_998 _17957_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19150_ _33508_/Q _33444_/Q _33380_/Q _33316_/Q _19070_/X _19071_/X VGND VGND VPWR
+ VPWR _19150_/X sky130_fd_sc_hd__mux4_1
X_28348_ _28348_/A VGND VGND VPWR VPWR _34497_/D sky130_fd_sc_hd__clkbuf_1
X_16362_ _16357_/X _16359_/X _16360_/X _16361_/X VGND VGND VPWR VPWR _16362_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18101_ _18097_/X _18100_/X _17834_/X VGND VGND VPWR VPWR _18123_/A sky130_fd_sc_hd__o21ba_2
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16293_ _17860_/A VGND VGND VPWR VPWR _16293_/X sky130_fd_sc_hd__buf_4
XFILLER_9_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19081_ _32994_/Q _32930_/Q _32866_/Q _32802_/Q _18936_/X _18937_/X VGND VGND VPWR
+ VPWR _19081_/X sky130_fd_sc_hd__mux4_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28279_ _34465_/Q _24304_/X _28279_/S VGND VGND VPWR VPWR _28280_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18032_ _18028_/X _18031_/X _17867_/X VGND VGND VPWR VPWR _18033_/D sky130_fd_sc_hd__o21ba_1
X_30310_ _30310_/A VGND VGND VPWR VPWR _35396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31290_ _31290_/A VGND VGND VPWR VPWR _35860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_1265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30241_ _30241_/A VGND VGND VPWR VPWR _35363_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30172_ _35331_/Q _29216_/X _30184_/S VGND VGND VPWR VPWR _30173_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19983_ _19983_/A VGND VGND VPWR VPWR _32123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18934_ _18649_/X _18932_/X _18933_/X _18655_/X VGND VGND VPWR VPWR _18934_/X sky130_fd_sc_hd__a22o_1
X_34980_ _36004_/CLK _34980_/D VGND VGND VPWR VPWR _34980_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1320 input54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1331 _20147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33931_ _35273_/CLK _33931_/D VGND VGND VPWR VPWR _33931_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1342 _22434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18865_ _18861_/X _18864_/X _18722_/X VGND VGND VPWR VPWR _18891_/A sky130_fd_sc_hd__o21ba_1
XANTENNA_1353 _21191_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1364 _24273_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1375 _26497_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1386 _31408_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17816_ _17812_/X _17815_/X _17500_/X VGND VGND VPWR VPWR _17824_/C sky130_fd_sc_hd__o21ba_1
XFILLER_227_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33862_ _35784_/CLK _33862_/D VGND VGND VPWR VPWR _33862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18796_ _20208_/A VGND VGND VPWR VPWR _18796_/X sky130_fd_sc_hd__buf_4
XFILLER_227_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35601_ _35666_/CLK _35601_/D VGND VGND VPWR VPWR _35601_/Q sky130_fd_sc_hd__dfxtp_1
X_32813_ _36080_/CLK _32813_/D VGND VGND VPWR VPWR _32813_/Q sky130_fd_sc_hd__dfxtp_1
X_17747_ _17502_/X _17745_/X _17746_/X _17505_/X VGND VGND VPWR VPWR _17747_/X sky130_fd_sc_hd__a22o_1
XFILLER_54_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33793_ _33793_/CLK _33793_/D VGND VGND VPWR VPWR _33793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_894 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35532_ _35532_/CLK _35532_/D VGND VGND VPWR VPWR _35532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32744_ _36137_/CLK _32744_/D VGND VGND VPWR VPWR _32744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17678_ _34555_/Q _32443_/Q _34427_/Q _34363_/Q _17578_/X _17579_/X VGND VGND VPWR
+ VPWR _17678_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19417_ _19413_/X _19416_/X _19108_/X VGND VGND VPWR VPWR _19418_/D sky130_fd_sc_hd__o21ba_1
X_35463_ _35590_/CLK _35463_/D VGND VGND VPWR VPWR _35463_/Q sky130_fd_sc_hd__dfxtp_1
X_16629_ _34014_/Q _33950_/Q _33886_/Q _32158_/Q _16314_/X _16315_/X VGND VGND VPWR
+ VPWR _16629_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32675_ _36132_/CLK _32675_/D VGND VGND VPWR VPWR _32675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34414_ _35052_/CLK _34414_/D VGND VGND VPWR VPWR _34414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19348_ _33770_/Q _33706_/Q _33642_/Q _33578_/Q _19143_/X _19144_/X VGND VGND VPWR
+ VPWR _19348_/X sky130_fd_sc_hd__mux4_1
X_31626_ _36020_/Q input32/X _31628_/S VGND VGND VPWR VPWR _31627_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35394_ _35909_/CLK _35394_/D VGND VGND VPWR VPWR _35394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34345_ _35944_/CLK _34345_/D VGND VGND VPWR VPWR _34345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31557_ _35987_/Q input56/X _31565_/S VGND VGND VPWR VPWR _31558_/A sky130_fd_sc_hd__mux2_1
X_19279_ _34280_/Q _34216_/Q _34152_/Q _34088_/Q _19036_/X _19037_/X VGND VGND VPWR
+ VPWR _19279_/X sky130_fd_sc_hd__mux4_1
XFILLER_202_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21310_ _22508_/A VGND VGND VPWR VPWR _21310_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_108_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30508_ _30598_/S VGND VGND VPWR VPWR _30527_/S sky130_fd_sc_hd__buf_6
X_22290_ _22286_/X _22289_/X _22081_/X VGND VGND VPWR VPWR _22320_/A sky130_fd_sc_hd__o21ba_1
X_34276_ _34276_/CLK _34276_/D VGND VGND VPWR VPWR _34276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31488_ _31488_/A VGND VGND VPWR VPWR _35954_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36015_ _36015_/CLK _36015_/D VGND VGND VPWR VPWR _36015_/Q sky130_fd_sc_hd__dfxtp_1
X_33227_ _34251_/CLK _33227_/D VGND VGND VPWR VPWR _33227_/Q sky130_fd_sc_hd__dfxtp_1
X_21241_ _22455_/A VGND VGND VPWR VPWR _21241_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_89_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30439_ _23307_/X _35457_/Q _30455_/S VGND VGND VPWR VPWR _30440_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33158_ _36166_/CLK _33158_/D VGND VGND VPWR VPWR _33158_/Q sky130_fd_sc_hd__dfxtp_1
X_21172_ _32988_/Q _32924_/Q _32860_/Q _32796_/Q _20883_/X _20884_/X VGND VGND VPWR
+ VPWR _21172_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20123_ _20119_/X _20122_/X _19814_/X VGND VGND VPWR VPWR _20124_/D sky130_fd_sc_hd__o21ba_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32109_ _35552_/CLK _32109_/D VGND VGND VPWR VPWR _32109_/Q sky130_fd_sc_hd__dfxtp_1
X_25980_ _26007_/S VGND VGND VPWR VPWR _25999_/S sky130_fd_sc_hd__buf_4
X_33089_ _36161_/CLK _33089_/D VGND VGND VPWR VPWR _33089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20054_ _33790_/Q _33726_/Q _33662_/Q _33598_/Q _19849_/X _19850_/X VGND VGND VPWR
+ VPWR _20054_/X sky130_fd_sc_hd__mux4_1
X_24931_ _22991_/X _32946_/Q _24937_/S VGND VGND VPWR VPWR _24932_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27650_ _27650_/A VGND VGND VPWR VPWR _34166_/D sky130_fd_sc_hd__clkbuf_1
X_24862_ _22889_/X _32913_/Q _24874_/S VGND VGND VPWR VPWR _24863_/A sky130_fd_sc_hd__mux2_1
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26601_ _26601_/A VGND VGND VPWR VPWR _33701_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23813_ _23813_/A VGND VGND VPWR VPWR _32450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27581_ _34134_/Q _24270_/X _27583_/S VGND VGND VPWR VPWR _27582_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24793_ _24793_/A VGND VGND VPWR VPWR _32880_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29320_ _23247_/X _34927_/Q _29332_/S VGND VGND VPWR VPWR _29321_/A sky130_fd_sc_hd__mux2_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26532_ _26532_/A VGND VGND VPWR VPWR _33669_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_228 _32136_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23744_ _23834_/S VGND VGND VPWR VPWR _23763_/S sky130_fd_sc_hd__buf_6
XANTENNA_239 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20956_ _20949_/X _20951_/X _20954_/X _20955_/X VGND VGND VPWR VPWR _20956_/X sky130_fd_sc_hd__a22o_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29251_ _23077_/X _34894_/Q _29269_/S VGND VGND VPWR VPWR _29252_/A sky130_fd_sc_hd__mux2_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23675_ _23675_/A VGND VGND VPWR VPWR _32386_/D sky130_fd_sc_hd__clkbuf_1
X_26463_ _26463_/A VGND VGND VPWR VPWR _33636_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20887_ _20881_/X _20886_/X _20640_/X _20642_/X VGND VGND VPWR VPWR _20908_/B sky130_fd_sc_hd__o211a_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28202_ _28202_/A VGND VGND VPWR VPWR _34428_/D sky130_fd_sc_hd__clkbuf_1
X_22626_ _34821_/Q _34757_/Q _34693_/Q _34629_/Q _22594_/X _22595_/X VGND VGND VPWR
+ VPWR _22626_/X sky130_fd_sc_hd__mux4_1
XFILLER_241_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25414_ _25414_/A VGND VGND VPWR VPWR _33143_/D sky130_fd_sc_hd__clkbuf_1
X_26394_ _25159_/X _33604_/Q _26404_/S VGND VGND VPWR VPWR _26395_/A sky130_fd_sc_hd__mux2_1
X_29182_ input37/X VGND VGND VPWR VPWR _29182_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25345_ _25019_/X _33111_/Q _25345_/S VGND VGND VPWR VPWR _25346_/A sky130_fd_sc_hd__mux2_1
X_28133_ _28133_/A VGND VGND VPWR VPWR _34395_/D sky130_fd_sc_hd__clkbuf_1
X_22557_ _22557_/A VGND VGND VPWR VPWR _22557_/X sky130_fd_sc_hd__buf_4
XFILLER_155_805 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21508_ _21401_/X _21506_/X _21507_/X _21406_/X VGND VGND VPWR VPWR _21508_/X sky130_fd_sc_hd__a22o_1
XFILLER_181_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28064_ _26962_/X _34363_/Q _28072_/S VGND VGND VPWR VPWR _28065_/A sky130_fd_sc_hd__mux2_1
X_25276_ _25276_/A VGND VGND VPWR VPWR _33078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22488_ _35585_/Q _35521_/Q _35457_/Q _35393_/Q _22203_/X _22204_/X VGND VGND VPWR
+ VPWR _22488_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27015_ _27014_/X _33868_/Q _27018_/S VGND VGND VPWR VPWR _27016_/A sky130_fd_sc_hd__mux2_1
X_24227_ _24227_/A VGND VGND VPWR VPWR _32645_/D sky130_fd_sc_hd__clkbuf_1
X_21439_ _21435_/X _21438_/X _21408_/X VGND VGND VPWR VPWR _21440_/D sky130_fd_sc_hd__o21ba_1
XFILLER_182_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24158_ _24158_/A VGND VGND VPWR VPWR _32612_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23109_ _32149_/Q _23108_/X _23115_/S VGND VGND VPWR VPWR _23110_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24089_ _24089_/A VGND VGND VPWR VPWR _32580_/D sky130_fd_sc_hd__clkbuf_1
X_28966_ _28966_/A VGND VGND VPWR VPWR _34790_/D sky130_fd_sc_hd__clkbuf_1
X_16980_ _16842_/X _16978_/X _16979_/X _16847_/X VGND VGND VPWR VPWR _16980_/X sky130_fd_sc_hd__a22o_1
XFILLER_1_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27917_ _27917_/A VGND VGND VPWR VPWR _34293_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28897_ _26996_/X _34758_/Q _28903_/S VGND VGND VPWR VPWR _28898_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18650_ _20062_/A VGND VGND VPWR VPWR _18650_/X sky130_fd_sc_hd__buf_4
X_27848_ _27848_/A VGND VGND VPWR VPWR _34260_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17601_ _35769_/Q _35129_/Q _34489_/Q _33849_/Q _17493_/X _17494_/X VGND VGND VPWR
+ VPWR _17601_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18581_ _18314_/X _18579_/X _18580_/X _18323_/X VGND VGND VPWR VPWR _18581_/X sky130_fd_sc_hd__a22o_1
XFILLER_236_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27779_ _34228_/Q _24363_/X _27781_/S VGND VGND VPWR VPWR _27780_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29518_ _29518_/A VGND VGND VPWR VPWR _35021_/D sky130_fd_sc_hd__clkbuf_1
X_17532_ _35831_/Q _32209_/Q _35703_/Q _35639_/Q _17313_/X _17314_/X VGND VGND VPWR
+ VPWR _17532_/X sky130_fd_sc_hd__mux4_1
XTAP_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30790_ _30790_/A VGND VGND VPWR VPWR _35623_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_740 _21690_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_751 _22393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_762 _22500_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29449_ _23237_/X _34988_/Q _29467_/S VGND VGND VPWR VPWR _29450_/A sky130_fd_sc_hd__mux2_1
X_17463_ _17459_/X _17462_/X _17147_/X VGND VGND VPWR VPWR _17471_/C sky130_fd_sc_hd__o21ba_1
XFILLER_233_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_773 _22538_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_784 _22634_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_795 _22784_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19202_ _19196_/X _19201_/X _19094_/X VGND VGND VPWR VPWR _19210_/C sky130_fd_sc_hd__o21ba_1
XFILLER_232_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16414_ _33752_/Q _33688_/Q _33624_/Q _33560_/Q _16137_/X _16138_/X VGND VGND VPWR
+ VPWR _16414_/X sky130_fd_sc_hd__mux4_1
X_32460_ _35789_/CLK _32460_/D VGND VGND VPWR VPWR _32460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17394_ _17149_/X _17392_/X _17393_/X _17152_/X VGND VGND VPWR VPWR _17394_/X sky130_fd_sc_hd__a22o_1
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31411_ _31543_/S VGND VGND VPWR VPWR _31430_/S sky130_fd_sc_hd__buf_4
X_19133_ _34787_/Q _34723_/Q _34659_/Q _34595_/Q _18882_/X _18883_/X VGND VGND VPWR
+ VPWR _19133_/X sky130_fd_sc_hd__mux4_1
X_16345_ _33494_/Q _33430_/Q _33366_/Q _33302_/Q _15998_/X _15999_/X VGND VGND VPWR
+ VPWR _16345_/X sky130_fd_sc_hd__mux4_1
X_32391_ _32901_/CLK _32391_/D VGND VGND VPWR VPWR _32391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34130_ _34256_/CLK _34130_/D VGND VGND VPWR VPWR _34130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19064_ _19060_/X _19063_/X _18755_/X VGND VGND VPWR VPWR _19065_/D sky130_fd_sc_hd__o21ba_1
XFILLER_12_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31342_ _35885_/Q input25/X _31358_/S VGND VGND VPWR VPWR _31343_/A sky130_fd_sc_hd__mux2_1
X_16276_ _34004_/Q _33940_/Q _33876_/Q _32148_/Q _16108_/X _16109_/X VGND VGND VPWR
+ VPWR _16276_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18015_ _32517_/Q _32389_/Q _32069_/Q _36037_/Q _17982_/X _17770_/X VGND VGND VPWR
+ VPWR _18015_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34061_ _34316_/CLK _34061_/D VGND VGND VPWR VPWR _34061_/Q sky130_fd_sc_hd__dfxtp_1
X_31273_ _35853_/Q input60/X _31273_/S VGND VGND VPWR VPWR _31274_/A sky130_fd_sc_hd__mux2_1
X_33012_ _33013_/CLK _33012_/D VGND VGND VPWR VPWR _33012_/Q sky130_fd_sc_hd__dfxtp_1
X_30224_ _30224_/A VGND VGND VPWR VPWR _35355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19966_ _20095_/A VGND VGND VPWR VPWR _19966_/X sky130_fd_sc_hd__buf_6
X_30155_ _35323_/Q _29191_/X _30163_/S VGND VGND VPWR VPWR _30156_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18917_ _35293_/Q _35229_/Q _35165_/Q _32285_/Q _18600_/X _18601_/X VGND VGND VPWR
+ VPWR _18917_/X sky130_fd_sc_hd__mux4_1
X_34963_ _36204_/CLK _34963_/D VGND VGND VPWR VPWR _34963_/Q sky130_fd_sc_hd__dfxtp_1
X_19897_ _33017_/Q _32953_/Q _32889_/Q _32825_/Q _19642_/X _19643_/X VGND VGND VPWR
+ VPWR _19897_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1150 _19597_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30086_ _35290_/Q _29089_/X _30100_/S VGND VGND VPWR VPWR _30087_/A sky130_fd_sc_hd__mux2_1
XANTENNA_1161 _22557_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1172 _20660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1183 _22217_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33914_ _36154_/CLK _33914_/D VGND VGND VPWR VPWR _33914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18848_ _18593_/X _18846_/X _18847_/X _18596_/X VGND VGND VPWR VPWR _18848_/X sky130_fd_sc_hd__a22o_1
X_34894_ _35026_/CLK _34894_/D VGND VGND VPWR VPWR _34894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1194 _22914_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33845_ _35828_/CLK _33845_/D VGND VGND VPWR VPWR _33845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18779_ _18775_/X _18778_/X _18741_/X VGND VGND VPWR VPWR _18787_/C sky130_fd_sc_hd__o21ba_1
XFILLER_212_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20810_ _34002_/Q _33938_/Q _33874_/Q _32146_/Q _20708_/X _20709_/X VGND VGND VPWR
+ VPWR _20810_/X sky130_fd_sc_hd__mux4_1
X_21790_ _35053_/Q _34989_/Q _34925_/Q _34861_/Q _21756_/X _21757_/X VGND VGND VPWR
+ VPWR _21790_/X sky130_fd_sc_hd__mux4_1
X_33776_ _34289_/CLK _33776_/D VGND VGND VPWR VPWR _33776_/Q sky130_fd_sc_hd__dfxtp_1
X_30988_ _30988_/A VGND VGND VPWR VPWR _35717_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35515_ _35515_/CLK _35515_/D VGND VGND VPWR VPWR _35515_/Q sky130_fd_sc_hd__dfxtp_1
X_20741_ _22458_/A VGND VGND VPWR VPWR _20741_/X sky130_fd_sc_hd__buf_4
X_32727_ _36055_/CLK _32727_/D VGND VGND VPWR VPWR _32727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23460_ _23460_/A VGND VGND VPWR VPWR _32285_/D sky130_fd_sc_hd__clkbuf_1
X_35446_ _35956_/CLK _35446_/D VGND VGND VPWR VPWR _35446_/Q sky130_fd_sc_hd__dfxtp_1
X_20672_ _20655_/X _20669_/X _20671_/X VGND VGND VPWR VPWR _20702_/C sky130_fd_sc_hd__o21ba_1
X_32658_ _36050_/CLK _32658_/D VGND VGND VPWR VPWR _32658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22411_ _35775_/Q _35135_/Q _34495_/Q _33855_/Q _22093_/X _22094_/X VGND VGND VPWR
+ VPWR _22411_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31609_ _31678_/S VGND VGND VPWR VPWR _31628_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_104_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23391_ _23391_/A VGND VGND VPWR VPWR _32254_/D sky130_fd_sc_hd__clkbuf_1
X_35377_ _35953_/CLK _35377_/D VGND VGND VPWR VPWR _35377_/Q sky130_fd_sc_hd__dfxtp_1
X_32589_ _35917_/CLK _32589_/D VGND VGND VPWR VPWR _32589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25130_ _25130_/A VGND VGND VPWR VPWR _33018_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22342_ _33213_/Q _32573_/Q _35965_/Q _35901_/Q _22027_/X _22028_/X VGND VGND VPWR
+ VPWR _22342_/X sky130_fd_sc_hd__mux4_1
X_34328_ _35292_/CLK _34328_/D VGND VGND VPWR VPWR _34328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25061_ _25060_/X _32996_/Q _25082_/S VGND VGND VPWR VPWR _25062_/A sky130_fd_sc_hd__mux2_1
X_34259_ _34259_/CLK _34259_/D VGND VGND VPWR VPWR _34259_/Q sky130_fd_sc_hd__dfxtp_1
X_22273_ _21952_/X _22271_/X _22272_/X _21955_/X VGND VGND VPWR VPWR _22273_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24012_ _22935_/X _32544_/Q _24014_/S VGND VGND VPWR VPWR _24013_/A sky130_fd_sc_hd__mux2_1
X_21224_ _21224_/A VGND VGND VPWR VPWR _36189_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28820_ _28820_/A VGND VGND VPWR VPWR _34721_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21155_ _21048_/X _21153_/X _21154_/X _21053_/X VGND VGND VPWR VPWR _21155_/X sky130_fd_sc_hd__a22o_1
X_20106_ _32511_/Q _32383_/Q _32063_/Q _36031_/Q _19929_/X _20070_/X VGND VGND VPWR
+ VPWR _20106_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28751_ _28751_/A VGND VGND VPWR VPWR _34688_/D sky130_fd_sc_hd__clkbuf_1
X_25963_ _25963_/A VGND VGND VPWR VPWR _33399_/D sky130_fd_sc_hd__clkbuf_1
X_21086_ _21082_/X _21085_/X _21055_/X VGND VGND VPWR VPWR _21087_/D sky130_fd_sc_hd__o21ba_1
X_27702_ _34191_/Q _24249_/X _27718_/S VGND VGND VPWR VPWR _27703_/A sky130_fd_sc_hd__mux2_1
X_20037_ _20033_/X _20036_/X _19789_/X _19790_/X VGND VGND VPWR VPWR _20052_/B sky130_fd_sc_hd__o211a_1
XFILLER_24_1248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24914_ _22966_/X _32938_/Q _24916_/S VGND VGND VPWR VPWR _24915_/A sky130_fd_sc_hd__mux2_1
X_28682_ _26878_/X _34656_/Q _28684_/S VGND VGND VPWR VPWR _28683_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25894_ _25019_/X _33367_/Q _25894_/S VGND VGND VPWR VPWR _25895_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27633_ _27633_/A VGND VGND VPWR VPWR _34158_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24845_ _24845_/A VGND VGND VPWR VPWR _32905_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27564_ _27696_/S VGND VGND VPWR VPWR _27583_/S sky130_fd_sc_hd__buf_6
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21988_ _35571_/Q _35507_/Q _35443_/Q _35379_/Q _21850_/X _21851_/X VGND VGND VPWR
+ VPWR _21988_/X sky130_fd_sc_hd__mux4_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24776_ _24776_/A VGND VGND VPWR VPWR _32872_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29303_ _23220_/X _34919_/Q _29311_/S VGND VGND VPWR VPWR _29304_/A sky130_fd_sc_hd__mux2_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26515_ _26515_/A VGND VGND VPWR VPWR _33661_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20939_ _20935_/X _20938_/X _20700_/X VGND VGND VPWR VPWR _20940_/D sky130_fd_sc_hd__o21ba_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23727_ _23727_/A VGND VGND VPWR VPWR _32409_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27495_ _26922_/X _34094_/Q _27509_/S VGND VGND VPWR VPWR _27496_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29234_ input55/X VGND VGND VPWR VPWR _29234_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_186_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26446_ _26446_/A VGND VGND VPWR VPWR _33628_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23658_ _23658_/A VGND VGND VPWR VPWR _32378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22609_ _34053_/Q _33989_/Q _33925_/Q _32261_/Q _22326_/X _22327_/X VGND VGND VPWR
+ VPWR _22609_/X sky130_fd_sc_hd__mux4_1
X_29165_ _29165_/A VGND VGND VPWR VPWR _34866_/D sky130_fd_sc_hd__clkbuf_1
X_26377_ _25134_/X _33596_/Q _26383_/S VGND VGND VPWR VPWR _26378_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23589_ _23589_/A VGND VGND VPWR VPWR _32345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16130_ _34511_/Q _32399_/Q _34383_/Q _34319_/Q _16088_/X _16090_/X VGND VGND VPWR
+ VPWR _16130_/X sky130_fd_sc_hd__mux4_1
X_28116_ _28116_/A VGND VGND VPWR VPWR _34387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25328_ _25328_/A VGND VGND VPWR VPWR _33102_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29096_ _34844_/Q _29095_/X _29111_/S VGND VGND VPWR VPWR _29097_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16061_ _35534_/Q _35470_/Q _35406_/Q _35342_/Q _16058_/X _16060_/X VGND VGND VPWR
+ VPWR _16061_/X sky130_fd_sc_hd__mux4_1
X_28047_ _26937_/X _34355_/Q _28051_/S VGND VGND VPWR VPWR _28048_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25259_ _25259_/A VGND VGND VPWR VPWR _33070_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19820_ _19495_/X _19818_/X _19819_/X _19500_/X VGND VGND VPWR VPWR _19820_/X sky130_fd_sc_hd__a22o_1
X_29998_ _29998_/A VGND VGND VPWR VPWR _35248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19751_ _33269_/Q _36149_/Q _33141_/Q _33077_/Q _19711_/X _19712_/X VGND VGND VPWR
+ VPWR _19751_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16963_ _35751_/Q _35111_/Q _34471_/Q _33831_/Q _16787_/X _16788_/X VGND VGND VPWR
+ VPWR _16963_/X sky130_fd_sc_hd__mux4_1
X_28949_ _28949_/A VGND VGND VPWR VPWR _34782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18702_ _33175_/Q _32535_/Q _35927_/Q _35863_/Q _18668_/X _18669_/X VGND VGND VPWR
+ VPWR _18702_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_28__f_CLK clkbuf_5_14_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_28__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_133_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31960_ _35036_/CLK _31960_/D VGND VGND VPWR VPWR _31960_/Q sky130_fd_sc_hd__dfxtp_1
X_19682_ _33011_/Q _32947_/Q _32883_/Q _32819_/Q _19642_/X _19643_/X VGND VGND VPWR
+ VPWR _19682_/X sky130_fd_sc_hd__mux4_1
X_16894_ _35813_/Q _32189_/Q _35685_/Q _35621_/Q _16607_/X _16608_/X VGND VGND VPWR
+ VPWR _16894_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18633_ _34773_/Q _34709_/Q _34645_/Q _34581_/Q _18529_/X _18530_/X VGND VGND VPWR
+ VPWR _18633_/X sky130_fd_sc_hd__mux4_1
X_30911_ _35681_/Q _29110_/X _30911_/S VGND VGND VPWR VPWR _30912_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31891_ _31891_/A VGND VGND VPWR VPWR _36145_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33630_ _34142_/CLK _33630_/D VGND VGND VPWR VPWR _33630_/Q sky130_fd_sc_hd__dfxtp_1
X_30842_ _23303_/X _35648_/Q _30860_/S VGND VGND VPWR VPWR _30843_/A sky130_fd_sc_hd__mux2_1
X_18564_ _35283_/Q _35219_/Q _35155_/Q _32275_/Q _18379_/X _18381_/X VGND VGND VPWR
+ VPWR _18564_/X sky130_fd_sc_hd__mux4_1
XTAP_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17515_ _17506_/X _17513_/X _17514_/X VGND VGND VPWR VPWR _17516_/D sky130_fd_sc_hd__o21ba_1
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33561_ _35671_/CLK _33561_/D VGND VGND VPWR VPWR _33561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18495_ _18356_/X _18493_/X _18494_/X _18368_/X VGND VGND VPWR VPWR _18495_/X sky130_fd_sc_hd__a22o_1
X_30773_ _30773_/A VGND VGND VPWR VPWR _35615_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_570 _20147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35300_ _35300_/CLK _35300_/D VGND VGND VPWR VPWR _35300_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32512_ _36032_/CLK _32512_/D VGND VGND VPWR VPWR _32512_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_581 _19449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_592 _19459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17446_ _33525_/Q _33461_/Q _33397_/Q _33333_/Q _17123_/X _17124_/X VGND VGND VPWR
+ VPWR _17446_/X sky130_fd_sc_hd__mux4_1
X_33492_ _33940_/CLK _33492_/D VGND VGND VPWR VPWR _33492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35231_ _35296_/CLK _35231_/D VGND VGND VPWR VPWR _35231_/Q sky130_fd_sc_hd__dfxtp_1
X_32443_ _35579_/CLK _32443_/D VGND VGND VPWR VPWR _32443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17377_ _17371_/X _17376_/X _17128_/X VGND VGND VPWR VPWR _17399_/A sky130_fd_sc_hd__o21ba_1
XFILLER_207_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19116_ _34019_/Q _33955_/Q _33891_/Q _32163_/Q _18967_/X _18968_/X VGND VGND VPWR
+ VPWR _19116_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16328_ _16288_/X _16326_/X _16327_/X _16291_/X VGND VGND VPWR VPWR _16328_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35162_ _35164_/CLK _35162_/D VGND VGND VPWR VPWR _35162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32374_ _36022_/CLK _32374_/D VGND VGND VPWR VPWR _32374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34113_ _36165_/CLK _34113_/D VGND VGND VPWR VPWR _34113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31325_ _35877_/Q input16/X _31337_/S VGND VGND VPWR VPWR _31326_/A sky130_fd_sc_hd__mux2_1
X_19047_ _32481_/Q _32353_/Q _32033_/Q _36001_/Q _18870_/X _19011_/X VGND VGND VPWR
+ VPWR _19047_/X sky130_fd_sc_hd__mux4_1
X_35093_ _35730_/CLK _35093_/D VGND VGND VPWR VPWR _35093_/Q sky130_fd_sc_hd__dfxtp_1
X_16259_ _35539_/Q _35475_/Q _35411_/Q _35347_/Q _16191_/X _16192_/X VGND VGND VPWR
+ VPWR _16259_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput202 _36227_/Q VGND VGND VPWR VPWR D2[53] sky130_fd_sc_hd__buf_2
Xoutput213 _36237_/Q VGND VGND VPWR VPWR D2[63] sky130_fd_sc_hd__buf_2
XFILLER_161_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34044_ _34044_/CLK _34044_/D VGND VGND VPWR VPWR _34044_/Q sky130_fd_sc_hd__dfxtp_1
X_31256_ _31256_/A VGND VGND VPWR VPWR _35844_/D sky130_fd_sc_hd__clkbuf_1
Xoutput224 _32093_/Q VGND VGND VPWR VPWR D3[15] sky130_fd_sc_hd__buf_2
XFILLER_173_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput235 _32103_/Q VGND VGND VPWR VPWR D3[25] sky130_fd_sc_hd__buf_2
XFILLER_177_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput246 _32113_/Q VGND VGND VPWR VPWR D3[35] sky130_fd_sc_hd__buf_2
X_30207_ _30207_/A VGND VGND VPWR VPWR _35347_/D sky130_fd_sc_hd__clkbuf_1
Xoutput257 _32123_/Q VGND VGND VPWR VPWR D3[45] sky130_fd_sc_hd__buf_2
Xoutput268 _32133_/Q VGND VGND VPWR VPWR D3[55] sky130_fd_sc_hd__buf_2
Xoutput279 _32085_/Q VGND VGND VPWR VPWR D3[7] sky130_fd_sc_hd__buf_2
X_31187_ _31187_/A VGND VGND VPWR VPWR _35811_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30138_ _35315_/Q _29166_/X _30142_/S VGND VGND VPWR VPWR _30139_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19949_ _19945_/X _19948_/X _19814_/X VGND VGND VPWR VPWR _19950_/D sky130_fd_sc_hd__o21ba_1
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35995_ _35995_/CLK _35995_/D VGND VGND VPWR VPWR _35995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22960_ input19/X VGND VGND VPWR VPWR _22960_/X sky130_fd_sc_hd__clkbuf_4
X_34946_ _34947_/CLK _34946_/D VGND VGND VPWR VPWR _34946_/Q sky130_fd_sc_hd__dfxtp_1
X_30069_ _35282_/Q _29064_/X _30079_/S VGND VGND VPWR VPWR _30070_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21911_ _21663_/X _21909_/X _21910_/X _21667_/X VGND VGND VPWR VPWR _21911_/X sky130_fd_sc_hd__a22o_1
XFILLER_228_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22891_ _22891_/A VGND VGND VPWR VPWR _32017_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34877_ _35989_/CLK _34877_/D VGND VGND VPWR VPWR _34877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21842_ _21655_/X _21840_/X _21841_/X _21661_/X VGND VGND VPWR VPWR _21842_/X sky130_fd_sc_hd__a22o_1
X_24630_ _22948_/X _32804_/Q _24644_/S VGND VGND VPWR VPWR _24631_/A sky130_fd_sc_hd__mux2_1
X_33828_ _35941_/CLK _33828_/D VGND VGND VPWR VPWR _33828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24561_ _23050_/X _32773_/Q _24569_/S VGND VGND VPWR VPWR _24562_/A sky130_fd_sc_hd__mux2_1
X_21773_ _33261_/Q _36141_/Q _33133_/Q _33069_/Q _21658_/X _21659_/X VGND VGND VPWR
+ VPWR _21773_/X sky130_fd_sc_hd__mux4_1
X_33759_ _34271_/CLK _33759_/D VGND VGND VPWR VPWR _33759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26300_ _26300_/A VGND VGND VPWR VPWR _33559_/D sky130_fd_sc_hd__clkbuf_1
X_20724_ _33167_/Q _32527_/Q _35919_/Q _35855_/Q _20663_/X _20665_/X VGND VGND VPWR
+ VPWR _20724_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23512_ _23003_/X _32310_/Q _23530_/S VGND VGND VPWR VPWR _23513_/A sky130_fd_sc_hd__mux2_1
X_27280_ _27280_/A VGND VGND VPWR VPWR _33992_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24492_ _22948_/X _32740_/Q _24506_/S VGND VGND VPWR VPWR _24493_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23443_ _23443_/A VGND VGND VPWR VPWR _32277_/D sky130_fd_sc_hd__clkbuf_1
X_26231_ _26231_/A VGND VGND VPWR VPWR _33526_/D sky130_fd_sc_hd__clkbuf_1
X_20655_ _20644_/X _20647_/X _20652_/X _20654_/X VGND VGND VPWR VPWR _20655_/X sky130_fd_sc_hd__a22o_1
X_35429_ _35749_/CLK _35429_/D VGND VGND VPWR VPWR _35429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26162_ _25016_/X _33494_/Q _26164_/S VGND VGND VPWR VPWR _26163_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23374_ _32246_/Q _23270_/X _23392_/S VGND VGND VPWR VPWR _23375_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20586_ _22367_/A VGND VGND VPWR VPWR _22506_/A sky130_fd_sc_hd__buf_12
XFILLER_143_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22325_ _33533_/Q _33469_/Q _33405_/Q _33341_/Q _22076_/X _22077_/X VGND VGND VPWR
+ VPWR _22325_/X sky130_fd_sc_hd__mux4_1
X_25113_ _25112_/X _33013_/Q _25113_/S VGND VGND VPWR VPWR _25114_/A sky130_fd_sc_hd__mux2_1
X_26093_ _26093_/A VGND VGND VPWR VPWR _33461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29921_ _29921_/A VGND VGND VPWR VPWR _35212_/D sky130_fd_sc_hd__clkbuf_1
X_25044_ input9/X VGND VGND VPWR VPWR _25044_/X sky130_fd_sc_hd__clkbuf_4
X_22256_ _34043_/Q _33979_/Q _33915_/Q _32251_/Q _21973_/X _21974_/X VGND VGND VPWR
+ VPWR _22256_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21207_ _22395_/A VGND VGND VPWR VPWR _21207_/X sky130_fd_sc_hd__buf_4
X_29852_ _29852_/A VGND VGND VPWR VPWR _35179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_160_CLK clkbuf_6_30__f_CLK/X VGND VGND VPWR VPWR _35464_/CLK sky130_fd_sc_hd__clkbuf_16
X_22187_ _34297_/Q _34233_/Q _34169_/Q _34105_/Q _22042_/X _22043_/X VGND VGND VPWR
+ VPWR _22187_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_1348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28803_ _26857_/X _34713_/Q _28819_/S VGND VGND VPWR VPWR _28804_/A sky130_fd_sc_hd__mux2_1
X_21138_ _32987_/Q _32923_/Q _32859_/Q _32795_/Q _20883_/X _20884_/X VGND VGND VPWR
+ VPWR _21138_/X sky130_fd_sc_hd__mux4_1
X_29783_ _35147_/Q _29240_/X _29787_/S VGND VGND VPWR VPWR _29784_/A sky130_fd_sc_hd__mux2_1
X_26995_ _26995_/A VGND VGND VPWR VPWR _33861_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28734_ _28734_/A VGND VGND VPWR VPWR _34680_/D sky130_fd_sc_hd__clkbuf_1
X_21069_ _32473_/Q _32345_/Q _32025_/Q _35993_/Q _20817_/X _20958_/X VGND VGND VPWR
+ VPWR _21069_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25946_ _25946_/A VGND VGND VPWR VPWR _33391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28665_ _28776_/S VGND VGND VPWR VPWR _28684_/S sky130_fd_sc_hd__buf_4
X_25877_ _25877_/A VGND VGND VPWR VPWR _33358_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27616_ _27616_/A VGND VGND VPWR VPWR _34150_/D sky130_fd_sc_hd__clkbuf_1
X_24828_ _23038_/X _32897_/Q _24844_/S VGND VGND VPWR VPWR _24829_/A sky130_fd_sc_hd__mux2_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28596_ _26950_/X _34615_/Q _28612_/S VGND VGND VPWR VPWR _28597_/A sky130_fd_sc_hd__mux2_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_12_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_12_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27547_ _26999_/X _34119_/Q _27551_/S VGND VGND VPWR VPWR _27548_/A sky130_fd_sc_hd__mux2_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24759_ _24759_/A VGND VGND VPWR VPWR _32864_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _34289_/Q _34225_/Q _34161_/Q _34097_/Q _17089_/X _17090_/X VGND VGND VPWR
+ VPWR _17300_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18280_ _20202_/A VGND VGND VPWR VPWR _18280_/X sky130_fd_sc_hd__buf_8
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27478_ _26897_/X _34086_/Q _27488_/S VGND VGND VPWR VPWR _27479_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29217_ _34883_/Q _29216_/X _29235_/S VGND VGND VPWR VPWR _29218_/A sky130_fd_sc_hd__mux2_1
X_17231_ _17231_/A _17231_/B _17231_/C _17231_/D VGND VGND VPWR VPWR _17232_/A sky130_fd_sc_hd__or4_4
XFILLER_35_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26429_ _26429_/A VGND VGND VPWR VPWR _33620_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_27_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_27_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_204_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29148_ input25/X VGND VGND VPWR VPWR _29148_/X sky130_fd_sc_hd__clkbuf_4
X_17162_ _17153_/X _17160_/X _17161_/X VGND VGND VPWR VPWR _17163_/D sky130_fd_sc_hd__o21ba_1
XFILLER_183_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16113_ _32719_/Q _32655_/Q _32591_/Q _36047_/Q _17862_/A _17713_/A VGND VGND VPWR
+ VPWR _16113_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29079_ input64/X VGND VGND VPWR VPWR _29079_/X sky130_fd_sc_hd__buf_4
X_17093_ _33515_/Q _33451_/Q _33387_/Q _33323_/Q _16770_/X _16771_/X VGND VGND VPWR
+ VPWR _17093_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31110_ _31110_/A VGND VGND VPWR VPWR _35775_/D sky130_fd_sc_hd__clkbuf_1
X_16044_ _17855_/A VGND VGND VPWR VPWR _16044_/X sky130_fd_sc_hd__buf_4
XFILLER_196_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32090_ _35040_/CLK _32090_/D VGND VGND VPWR VPWR _32090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31041_ _31041_/A VGND VGND VPWR VPWR _35742_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_151_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _35147_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_237_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19803_ _34806_/Q _34742_/Q _34678_/Q _34614_/Q _19588_/X _19589_/X VGND VGND VPWR
+ VPWR _19803_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17995_ _17995_/A VGND VGND VPWR VPWR _17995_/X sky130_fd_sc_hd__buf_4
XFILLER_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34800_ _35061_/CLK _34800_/D VGND VGND VPWR VPWR _34800_/Q sky130_fd_sc_hd__dfxtp_1
X_16946_ _33767_/Q _33703_/Q _33639_/Q _33575_/Q _16843_/X _16844_/X VGND VGND VPWR
+ VPWR _16946_/X sky130_fd_sc_hd__mux4_1
X_19734_ _19449_/X _19732_/X _19733_/X _19452_/X VGND VGND VPWR VPWR _19734_/X sky130_fd_sc_hd__a22o_1
X_35780_ _35780_/CLK _35780_/D VGND VGND VPWR VPWR _35780_/Q sky130_fd_sc_hd__dfxtp_1
X_32992_ _36065_/CLK _32992_/D VGND VGND VPWR VPWR _32992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31943_ _31943_/A VGND VGND VPWR VPWR _36170_/D sky130_fd_sc_hd__clkbuf_1
X_34731_ _34986_/CLK _34731_/D VGND VGND VPWR VPWR _34731_/Q sky130_fd_sc_hd__dfxtp_1
X_19665_ _19454_/X _19663_/X _19664_/X _19459_/X VGND VGND VPWR VPWR _19665_/X sky130_fd_sc_hd__a22o_1
XFILLER_49_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16877_ _16871_/X _16876_/X _16808_/X VGND VGND VPWR VPWR _16878_/D sky130_fd_sc_hd__o21ba_1
XFILLER_225_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18616_ _34005_/Q _33941_/Q _33877_/Q _32149_/Q _18614_/X _18615_/X VGND VGND VPWR
+ VPWR _18616_/X sky130_fd_sc_hd__mux4_1
XTAP_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34662_ _35303_/CLK _34662_/D VGND VGND VPWR VPWR _34662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19596_ _19592_/X _19595_/X _19461_/X VGND VGND VPWR VPWR _19597_/D sky130_fd_sc_hd__o21ba_1
X_31874_ _31874_/A VGND VGND VPWR VPWR _36137_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33613_ _34124_/CLK _33613_/D VGND VGND VPWR VPWR _33613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18547_ _32723_/Q _32659_/Q _32595_/Q _36051_/Q _18513_/X _20013_/A VGND VGND VPWR
+ VPWR _18547_/X sky130_fd_sc_hd__mux4_1
X_30825_ _23277_/X _35640_/Q _30839_/S VGND VGND VPWR VPWR _30826_/A sky130_fd_sc_hd__mux2_1
XFILLER_234_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34593_ _35098_/CLK _34593_/D VGND VGND VPWR VPWR _34593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33544_ _33544_/CLK _33544_/D VGND VGND VPWR VPWR _33544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18478_ _34001_/Q _33937_/Q _33873_/Q _32145_/Q _18408_/X _18409_/X VGND VGND VPWR
+ VPWR _18478_/X sky130_fd_sc_hd__mux4_1
XFILLER_205_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30756_ _30756_/A VGND VGND VPWR VPWR _35607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17429_ _33204_/Q _32564_/Q _35956_/Q _35892_/Q _17427_/X _17428_/X VGND VGND VPWR
+ VPWR _17429_/X sky130_fd_sc_hd__mux4_1
X_33475_ _34050_/CLK _33475_/D VGND VGND VPWR VPWR _33475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30687_ _30687_/A VGND VGND VPWR VPWR _35574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_1099 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35214_ _36216_/CLK _35214_/D VGND VGND VPWR VPWR _35214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20440_ _35785_/Q _35145_/Q _34505_/Q _33865_/Q _20146_/X _20147_/X VGND VGND VPWR
+ VPWR _20440_/X sky130_fd_sc_hd__mux4_1
X_32426_ _35179_/CLK _32426_/D VGND VGND VPWR VPWR _32426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36194_ _36194_/CLK _36194_/D VGND VGND VPWR VPWR _36194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35145_ _35845_/CLK _35145_/D VGND VGND VPWR VPWR _35145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20371_ _20367_/X _20370_/X _20134_/X VGND VGND VPWR VPWR _20393_/A sky130_fd_sc_hd__o21ba_2
X_32357_ _36005_/CLK _32357_/D VGND VGND VPWR VPWR _32357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_390_CLK clkbuf_6_35__f_CLK/X VGND VGND VPWR VPWR _35313_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_162_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22110_ _22463_/A VGND VGND VPWR VPWR _22110_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_134_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31308_ _35869_/Q input7/X _31316_/S VGND VGND VPWR VPWR _31309_/A sky130_fd_sc_hd__mux2_1
X_35076_ _35779_/CLK _35076_/D VGND VGND VPWR VPWR _35076_/Q sky130_fd_sc_hd__dfxtp_1
X_23090_ input12/X VGND VGND VPWR VPWR _23090_/X sky130_fd_sc_hd__buf_4
XFILLER_115_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32288_ _35294_/CLK _32288_/D VGND VGND VPWR VPWR _32288_/Q sky130_fd_sc_hd__dfxtp_1
X_34027_ _36136_/CLK _34027_/D VGND VGND VPWR VPWR _34027_/Q sky130_fd_sc_hd__dfxtp_1
X_22041_ _33781_/Q _33717_/Q _33653_/Q _33589_/Q _21796_/X _21797_/X VGND VGND VPWR
+ VPWR _22041_/X sky130_fd_sc_hd__mux4_1
XTAP_6409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_142_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _35852_/CLK sky130_fd_sc_hd__clkbuf_16
X_31239_ _31239_/A VGND VGND VPWR VPWR _35836_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25800_ _25800_/A VGND VGND VPWR VPWR _33322_/D sky130_fd_sc_hd__clkbuf_1
X_26780_ _33786_/Q _24382_/X _26790_/S VGND VGND VPWR VPWR _26781_/A sky130_fd_sc_hd__mux2_1
X_35978_ _35978_/CLK _35978_/D VGND VGND VPWR VPWR _35978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23992_ _23992_/A VGND VGND VPWR VPWR _32534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25731_ _33291_/Q _24434_/X _25735_/S VGND VGND VPWR VPWR _25732_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_11__f_CLK clkbuf_5_5_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_11__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_34929_ _35954_/CLK _34929_/D VGND VGND VPWR VPWR _34929_/Q sky130_fd_sc_hd__dfxtp_1
X_22943_ _22941_/X _32034_/Q _22970_/S VGND VGND VPWR VPWR _22944_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28450_ _26934_/X _34546_/Q _28456_/S VGND VGND VPWR VPWR _28451_/A sky130_fd_sc_hd__mux2_1
X_25662_ _33258_/Q _24332_/X _25664_/S VGND VGND VPWR VPWR _25663_/A sky130_fd_sc_hd__mux2_1
X_22874_ _22874_/A VGND VGND VPWR VPWR _36237_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27401_ _27401_/A VGND VGND VPWR VPWR _34049_/D sky130_fd_sc_hd__clkbuf_1
X_24613_ _22923_/X _32796_/Q _24623_/S VGND VGND VPWR VPWR _24614_/A sky130_fd_sc_hd__mux2_1
X_28381_ _26832_/X _34513_/Q _28393_/S VGND VGND VPWR VPWR _28382_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21825_ _22531_/A VGND VGND VPWR VPWR _21825_/X sky130_fd_sc_hd__buf_6
X_25593_ _33227_/Q _24434_/X _25597_/S VGND VGND VPWR VPWR _25594_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27332_ _34017_/Q _24304_/X _27332_/S VGND VGND VPWR VPWR _27333_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_1013 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24544_ _23025_/X _32765_/Q _24548_/S VGND VGND VPWR VPWR _24545_/A sky130_fd_sc_hd__mux2_1
X_21756_ _22462_/A VGND VGND VPWR VPWR _21756_/X sky130_fd_sc_hd__buf_4
XFILLER_93_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20707_ _33487_/Q _33423_/Q _33359_/Q _33295_/Q _20598_/X _20599_/X VGND VGND VPWR
+ VPWR _20707_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27263_ _26977_/X _33984_/Q _27281_/S VGND VGND VPWR VPWR _27264_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21687_ _21687_/A VGND VGND VPWR VPWR _36202_/D sky130_fd_sc_hd__clkbuf_1
X_24475_ _22923_/X _32732_/Q _24485_/S VGND VGND VPWR VPWR _24476_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29002_ _29002_/A VGND VGND VPWR VPWR _34807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26214_ _26214_/A VGND VGND VPWR VPWR _33518_/D sky130_fd_sc_hd__clkbuf_1
X_23426_ _29384_/A _30735_/B VGND VGND VPWR VPWR _23559_/S sky130_fd_sc_hd__nand2_8
X_20638_ _20626_/X _20631_/X _20636_/X _20637_/X VGND VGND VPWR VPWR _20638_/X sky130_fd_sc_hd__a22o_1
XFILLER_109_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27194_ _27194_/A VGND VGND VPWR VPWR _33951_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26145_ _26277_/S VGND VGND VPWR VPWR _26164_/S sky130_fd_sc_hd__buf_4
X_23357_ _32238_/Q _23244_/X _23371_/S VGND VGND VPWR VPWR _23358_/A sky130_fd_sc_hd__mux2_1
X_20569_ _34573_/Q _32461_/Q _34445_/Q _34381_/Q _18363_/X _18365_/X VGND VGND VPWR
+ VPWR _20569_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_381_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _35953_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_165_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22308_ _22465_/A VGND VGND VPWR VPWR _22308_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_153_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23288_ _23288_/A VGND VGND VPWR VPWR _32213_/D sky130_fd_sc_hd__clkbuf_1
X_26076_ _25088_/X _33453_/Q _26092_/S VGND VGND VPWR VPWR _26077_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29904_ _35204_/Q _29219_/X _29914_/S VGND VGND VPWR VPWR _29905_/A sky130_fd_sc_hd__mux2_1
X_22239_ _21952_/X _22237_/X _22238_/X _21955_/X VGND VGND VPWR VPWR _22239_/X sky130_fd_sc_hd__a22o_1
X_25027_ _25026_/X _32985_/Q _25051_/S VGND VGND VPWR VPWR _25028_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_133_CLK clkbuf_6_23__f_CLK/X VGND VGND VPWR VPWR _34262_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29835_ _35171_/Q _29117_/X _29851_/S VGND VGND VPWR VPWR _29836_/A sky130_fd_sc_hd__mux2_1
XTAP_6943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16800_ _16796_/X _16797_/X _16798_/X _16799_/X VGND VGND VPWR VPWR _16800_/X sky130_fd_sc_hd__a22o_1
XTAP_6987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29766_ _29766_/A VGND VGND VPWR VPWR _35138_/D sky130_fd_sc_hd__clkbuf_1
X_17780_ _17931_/A VGND VGND VPWR VPWR _17780_/X sky130_fd_sc_hd__buf_6
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26978_ _27018_/S VGND VGND VPWR VPWR _27006_/S sky130_fd_sc_hd__buf_4
XFILLER_93_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16731_ _16448_/X _16729_/X _16730_/X _16453_/X VGND VGND VPWR VPWR _16731_/X sky130_fd_sc_hd__a22o_1
X_28717_ _28717_/A VGND VGND VPWR VPWR _34672_/D sky130_fd_sc_hd__clkbuf_1
X_25929_ _25929_/A VGND VGND VPWR VPWR _33383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29697_ _29787_/S VGND VGND VPWR VPWR _29716_/S sky130_fd_sc_hd__buf_4
XFILLER_234_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19450_ _34796_/Q _34732_/Q _34668_/Q _34604_/Q _19235_/X _19236_/X VGND VGND VPWR
+ VPWR _19450_/X sky130_fd_sc_hd__mux4_1
XFILLER_207_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28648_ _28648_/A VGND VGND VPWR VPWR _34639_/D sky130_fd_sc_hd__clkbuf_1
X_16662_ _16662_/A VGND VGND VPWR VPWR _31966_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18401_ _18385_/X _18398_/X _18400_/X VGND VGND VPWR VPWR _18402_/D sky130_fd_sc_hd__o21ba_1
XFILLER_34_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19381_ _19096_/X _19379_/X _19380_/X _19099_/X VGND VGND VPWR VPWR _19381_/X sky130_fd_sc_hd__a22o_1
XFILLER_216_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28579_ _26925_/X _34607_/Q _28591_/S VGND VGND VPWR VPWR _28580_/A sky130_fd_sc_hd__mux2_1
X_16593_ _33757_/Q _33693_/Q _33629_/Q _33565_/Q _16490_/X _16491_/X VGND VGND VPWR
+ VPWR _16593_/X sky130_fd_sc_hd__mux4_1
X_30610_ _35538_/Q _29064_/X _30620_/S VGND VGND VPWR VPWR _30611_/A sky130_fd_sc_hd__mux2_1
X_18332_ _18357_/A VGND VGND VPWR VPWR _20129_/A sky130_fd_sc_hd__buf_12
XFILLER_91_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31590_ _31590_/A VGND VGND VPWR VPWR _36002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18263_ _33229_/Q _32589_/Q _35981_/Q _35917_/Q _16075_/X _16076_/X VGND VGND VPWR
+ VPWR _18263_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30541_ _30541_/A VGND VGND VPWR VPWR _35505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17214_ _17210_/X _17213_/X _17136_/X _17137_/X VGND VGND VPWR VPWR _17231_/B sky130_fd_sc_hd__o211a_1
XFILLER_147_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33260_ _36146_/CLK _33260_/D VGND VGND VPWR VPWR _33260_/Q sky130_fd_sc_hd__dfxtp_1
X_18194_ _17149_/A _18192_/X _18193_/X _17152_/A VGND VGND VPWR VPWR _18194_/X sky130_fd_sc_hd__a22o_1
X_30472_ _30472_/A VGND VGND VPWR VPWR _35472_/D sky130_fd_sc_hd__clkbuf_1
X_32211_ _35833_/CLK _32211_/D VGND VGND VPWR VPWR _32211_/Q sky130_fd_sc_hd__dfxtp_1
X_17145_ _33196_/Q _32556_/Q _35948_/Q _35884_/Q _17074_/X _17075_/X VGND VGND VPWR
+ VPWR _17145_/X sky130_fd_sc_hd__mux4_1
X_33191_ _35943_/CLK _33191_/D VGND VGND VPWR VPWR _33191_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_372_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _36080_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32142_ _35664_/CLK _32142_/D VGND VGND VPWR VPWR _32142_/Q sky130_fd_sc_hd__dfxtp_1
X_17076_ _33194_/Q _32554_/Q _35946_/Q _35882_/Q _17074_/X _17075_/X VGND VGND VPWR
+ VPWR _17076_/X sky130_fd_sc_hd__mux4_1
XFILLER_171_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16027_ _16057_/A VGND VGND VPWR VPWR _17982_/A sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_124_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _33490_/CLK sky130_fd_sc_hd__clkbuf_16
X_32073_ _36041_/CLK _32073_/D VGND VGND VPWR VPWR _32073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31024_ _31024_/A VGND VGND VPWR VPWR _35734_/D sky130_fd_sc_hd__clkbuf_1
X_35901_ _35965_/CLK _35901_/D VGND VGND VPWR VPWR _35901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35832_ _35833_/CLK _35832_/D VGND VGND VPWR VPWR _35832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17978_ _17978_/A VGND VGND VPWR VPWR _17978_/X sky130_fd_sc_hd__buf_6
X_16929_ _35750_/Q _35110_/Q _34470_/Q _33830_/Q _16787_/X _16788_/X VGND VGND VPWR
+ VPWR _16929_/X sky130_fd_sc_hd__mux4_1
X_19717_ _20070_/A VGND VGND VPWR VPWR _19717_/X sky130_fd_sc_hd__clkbuf_4
X_32975_ _35984_/CLK _32975_/D VGND VGND VPWR VPWR _32975_/Q sky130_fd_sc_hd__dfxtp_1
X_35763_ _35765_/CLK _35763_/D VGND VGND VPWR VPWR _35763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34714_ _34779_/CLK _34714_/D VGND VGND VPWR VPWR _34714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31926_ _23310_/X _36162_/Q _31940_/S VGND VGND VPWR VPWR _31927_/A sky130_fd_sc_hd__mux2_1
X_19648_ _35826_/Q _32203_/Q _35698_/Q _35634_/Q _19613_/X _19614_/X VGND VGND VPWR
+ VPWR _19648_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35694_ _35822_/CLK _35694_/D VGND VGND VPWR VPWR _35694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34645_ _36189_/CLK _34645_/D VGND VGND VPWR VPWR _34645_/Q sky130_fd_sc_hd__dfxtp_1
X_19579_ _19363_/X _19577_/X _19578_/X _19367_/X VGND VGND VPWR VPWR _19579_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31857_ _31857_/A VGND VGND VPWR VPWR _36129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21610_ _34536_/Q _32424_/Q _34408_/Q _34344_/Q _21472_/X _21473_/X VGND VGND VPWR
+ VPWR _21610_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30808_ _23250_/X _35632_/Q _30818_/S VGND VGND VPWR VPWR _30809_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22590_ _35588_/Q _35524_/Q _35460_/Q _35396_/Q _22556_/X _22557_/X VGND VGND VPWR
+ VPWR _22590_/X sky130_fd_sc_hd__mux4_1
X_34576_ _35280_/CLK _34576_/D VGND VGND VPWR VPWR _34576_/Q sky130_fd_sc_hd__dfxtp_1
X_31788_ _31788_/A VGND VGND VPWR VPWR _36096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21541_ _35046_/Q _34982_/Q _34918_/Q _34854_/Q _21403_/X _21404_/X VGND VGND VPWR
+ VPWR _21541_/X sky130_fd_sc_hd__mux4_1
XFILLER_244_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30739_ _23090_/X _35599_/Q _30755_/S VGND VGND VPWR VPWR _30740_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33527_ _34039_/CLK _33527_/D VGND VGND VPWR VPWR _33527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24260_ _24260_/A VGND VGND VPWR VPWR _32658_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21472_ _22312_/A VGND VGND VPWR VPWR _21472_/X sky130_fd_sc_hd__buf_6
X_33458_ _33775_/CLK _33458_/D VGND VGND VPWR VPWR _33458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23211_ _32187_/Q _23152_/X _23235_/S VGND VGND VPWR VPWR _23212_/A sky130_fd_sc_hd__mux2_1
X_20423_ _20423_/A _20423_/B _20423_/C _20423_/D VGND VGND VPWR VPWR _20424_/A sky130_fd_sc_hd__or4_1
X_32409_ _35293_/CLK _32409_/D VGND VGND VPWR VPWR _32409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24191_ _24191_/A VGND VGND VPWR VPWR _32628_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36177_ _36185_/CLK _36177_/D VGND VGND VPWR VPWR _36177_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_363_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _33775_/CLK sky130_fd_sc_hd__clkbuf_16
X_33389_ _34292_/CLK _33389_/D VGND VGND VPWR VPWR _33389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23142_ input10/X VGND VGND VPWR VPWR _23142_/X sky130_fd_sc_hd__buf_4
X_20354_ _18297_/X _20352_/X _20353_/X _18303_/X VGND VGND VPWR VPWR _20354_/X sky130_fd_sc_hd__a22o_1
X_35128_ _35766_/CLK _35128_/D VGND VGND VPWR VPWR _35128_/Q sky130_fd_sc_hd__dfxtp_1
X_27950_ _34309_/Q _24416_/X _27958_/S VGND VGND VPWR VPWR _27951_/A sky130_fd_sc_hd__mux2_1
X_23073_ _23073_/A VGND VGND VPWR VPWR _32076_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_115_CLK clkbuf_6_20__f_CLK/X VGND VGND VPWR VPWR _36216_/CLK sky130_fd_sc_hd__clkbuf_16
X_35059_ _35827_/CLK _35059_/D VGND VGND VPWR VPWR _35059_/Q sky130_fd_sc_hd__dfxtp_1
X_20285_ _20069_/X _20283_/X _20284_/X _20073_/X VGND VGND VPWR VPWR _20285_/X sky130_fd_sc_hd__a22o_1
XTAP_6206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26901_ _26900_/X _33831_/Q _26913_/S VGND VGND VPWR VPWR _26902_/A sky130_fd_sc_hd__mux2_1
X_22024_ _35764_/Q _35124_/Q _34484_/Q _33844_/Q _21740_/X _21741_/X VGND VGND VPWR
+ VPWR _22024_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27881_ _34276_/Q _24314_/X _27895_/S VGND VGND VPWR VPWR _27882_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29620_ _29620_/A VGND VGND VPWR VPWR _35069_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26832_ input34/X VGND VGND VPWR VPWR _26832_/X sky130_fd_sc_hd__buf_4
XTAP_5549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29551_ _29551_/A VGND VGND VPWR VPWR _35036_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26763_ _33778_/Q _24357_/X _26769_/S VGND VGND VPWR VPWR _26764_/A sky130_fd_sc_hd__mux2_1
X_23975_ _22875_/X _32526_/Q _23993_/S VGND VGND VPWR VPWR _23976_/A sky130_fd_sc_hd__mux2_1
XTAP_4859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28502_ _27011_/X _34571_/Q _28506_/S VGND VGND VPWR VPWR _28503_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25714_ _25714_/A VGND VGND VPWR VPWR _33282_/D sky130_fd_sc_hd__clkbuf_1
X_29482_ _23289_/X _35004_/Q _29488_/S VGND VGND VPWR VPWR _29483_/A sky130_fd_sc_hd__mux2_1
X_22926_ input7/X VGND VGND VPWR VPWR _22926_/X sky130_fd_sc_hd__buf_6
XFILLER_17_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26694_ _33745_/Q _24255_/X _26706_/S VGND VGND VPWR VPWR _26695_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28433_ _26909_/X _34538_/Q _28435_/S VGND VGND VPWR VPWR _28434_/A sky130_fd_sc_hd__mux2_1
X_25645_ _25735_/S VGND VGND VPWR VPWR _25664_/S sky130_fd_sc_hd__buf_4
XFILLER_231_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22857_ _21754_/A _22855_/X _22856_/X _21759_/A VGND VGND VPWR VPWR _22857_/X sky130_fd_sc_hd__a22o_1
XFILLER_232_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28364_ _28364_/A VGND VGND VPWR VPWR _34505_/D sky130_fd_sc_hd__clkbuf_1
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21808_ _32750_/Q _32686_/Q _32622_/Q _36078_/Q _21519_/X _21656_/X VGND VGND VPWR
+ VPWR _21808_/X sky130_fd_sc_hd__mux4_1
X_25576_ _25576_/A VGND VGND VPWR VPWR _33218_/D sky130_fd_sc_hd__clkbuf_1
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22788_ _33547_/Q _33483_/Q _33419_/Q _33355_/Q _20633_/X _20635_/X VGND VGND VPWR
+ VPWR _22788_/X sky130_fd_sc_hd__mux4_2
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27315_ _27315_/A VGND VGND VPWR VPWR _34008_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24527_ _23000_/X _32757_/Q _24527_/S VGND VGND VPWR VPWR _24528_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28295_ _28295_/A VGND VGND VPWR VPWR _34472_/D sky130_fd_sc_hd__clkbuf_1
X_21739_ _35820_/Q _32197_/Q _35692_/Q _35628_/Q _21560_/X _21561_/X VGND VGND VPWR
+ VPWR _21739_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27246_ _26953_/X _33976_/Q _27260_/S VGND VGND VPWR VPWR _27247_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24458_ _22898_/X _32724_/Q _24464_/S VGND VGND VPWR VPWR _24459_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23409_ _32263_/Q _23327_/X _23413_/S VGND VGND VPWR VPWR _23410_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27177_ _27177_/A VGND VGND VPWR VPWR _33943_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_354_CLK clkbuf_6_44__f_CLK/X VGND VGND VPWR VPWR _35765_/CLK sky130_fd_sc_hd__clkbuf_16
X_24389_ _32700_/Q _24388_/X _24398_/S VGND VGND VPWR VPWR _24390_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_9 _32114_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26128_ _25165_/X _33478_/Q _26134_/S VGND VGND VPWR VPWR _26129_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_106_CLK clkbuf_6_22__f_CLK/X VGND VGND VPWR VPWR _35793_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_158_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26059_ _25063_/X _33445_/Q _26071_/S VGND VGND VPWR VPWR _26060_/A sky130_fd_sc_hd__mux2_1
X_18950_ _18946_/X _18947_/X _18948_/X _18949_/X VGND VGND VPWR VPWR _18950_/X sky130_fd_sc_hd__a22o_1
X_17901_ _17901_/A VGND VGND VPWR VPWR _17901_/X sky130_fd_sc_hd__buf_4
XFILLER_152_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18881_ _18877_/X _18880_/X _18741_/X VGND VGND VPWR VPWR _18891_/C sky130_fd_sc_hd__o21ba_1
XTAP_6740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17832_ _34048_/Q _33984_/Q _33920_/Q _32256_/Q _17726_/X _17727_/X VGND VGND VPWR
+ VPWR _17832_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29818_ _35163_/Q _29092_/X _29830_/S VGND VGND VPWR VPWR _29819_/A sky130_fd_sc_hd__mux2_1
XTAP_6784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17763_ _32766_/Q _32702_/Q _32638_/Q _36094_/Q _17625_/X _17762_/X VGND VGND VPWR
+ VPWR _17763_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29749_ _29749_/A VGND VGND VPWR VPWR _35130_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16714_ _17911_/A VGND VGND VPWR VPWR _16714_/X sky130_fd_sc_hd__clkbuf_4
X_19502_ _20208_/A VGND VGND VPWR VPWR _19502_/X sky130_fd_sc_hd__clkbuf_4
X_32760_ _36089_/CLK _32760_/D VGND VGND VPWR VPWR _32760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17694_ _32508_/Q _32380_/Q _32060_/Q _36028_/Q _17629_/X _17417_/X VGND VGND VPWR
+ VPWR _17694_/X sky130_fd_sc_hd__mux4_1
XFILLER_207_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19433_ _32492_/Q _32364_/Q _32044_/Q _36012_/Q _19223_/X _19364_/X VGND VGND VPWR
+ VPWR _19433_/X sky130_fd_sc_hd__mux4_1
X_31711_ _36060_/Q input6/X _31721_/S VGND VGND VPWR VPWR _31712_/A sky130_fd_sc_hd__mux2_1
X_16645_ _16641_/X _16642_/X _16643_/X _16644_/X VGND VGND VPWR VPWR _16645_/X sky130_fd_sc_hd__a22o_1
XFILLER_35_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32691_ _34032_/CLK _32691_/D VGND VGND VPWR VPWR _32691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34430_ _35581_/CLK _34430_/D VGND VGND VPWR VPWR _34430_/Q sky130_fd_sc_hd__dfxtp_1
X_31642_ _31642_/A VGND VGND VPWR VPWR _36027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19364_ _20070_/A VGND VGND VPWR VPWR _19364_/X sky130_fd_sc_hd__clkbuf_8
X_16576_ _35740_/Q _35100_/Q _34460_/Q _33820_/Q _16434_/X _16435_/X VGND VGND VPWR
+ VPWR _16576_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18315_ _18357_/A VGND VGND VPWR VPWR _20278_/A sky130_fd_sc_hd__buf_12
XFILLER_128_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34361_ _35577_/CLK _34361_/D VGND VGND VPWR VPWR _34361_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19295_ _35816_/Q _32192_/Q _35688_/Q _35624_/Q _19260_/X _19261_/X VGND VGND VPWR
+ VPWR _19295_/X sky130_fd_sc_hd__mux4_1
X_31573_ _31573_/A VGND VGND VPWR VPWR _35994_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_1358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36100_ _36100_/CLK _36100_/D VGND VGND VPWR VPWR _36100_/Q sky130_fd_sc_hd__dfxtp_1
X_33312_ _33692_/CLK _33312_/D VGND VGND VPWR VPWR _33312_/Q sky130_fd_sc_hd__dfxtp_1
X_18246_ _34317_/Q _34253_/Q _34189_/Q _34125_/Q _16045_/X _16046_/X VGND VGND VPWR
+ VPWR _18246_/X sky130_fd_sc_hd__mux4_1
X_30524_ _30524_/A VGND VGND VPWR VPWR _35497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34292_ _34292_/CLK _34292_/D VGND VGND VPWR VPWR _34292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36031_ _36031_/CLK _36031_/D VGND VGND VPWR VPWR _36031_/Q sky130_fd_sc_hd__dfxtp_1
X_33243_ _34265_/CLK _33243_/D VGND VGND VPWR VPWR _33243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18177_ _35338_/Q _35274_/Q _35210_/Q _32330_/Q _16088_/X _16090_/X VGND VGND VPWR
+ VPWR _18177_/X sky130_fd_sc_hd__mux4_1
X_30455_ _23333_/X _35465_/Q _30455_/S VGND VGND VPWR VPWR _30456_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_345_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _34292_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17128_ _17834_/A VGND VGND VPWR VPWR _17128_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_237_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33174_ _36117_/CLK _33174_/D VGND VGND VPWR VPWR _33174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30386_ _23223_/X _35432_/Q _30392_/S VGND VGND VPWR VPWR _30387_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32125_ _35562_/CLK _32125_/D VGND VGND VPWR VPWR _32125_/Q sky130_fd_sc_hd__dfxtp_1
X_17059_ _17770_/A VGND VGND VPWR VPWR _17059_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_217_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20070_ _20070_/A VGND VGND VPWR VPWR _20070_/X sky130_fd_sc_hd__clkbuf_4
X_32056_ _36024_/CLK _32056_/D VGND VGND VPWR VPWR _32056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31007_ _35726_/Q _29048_/X _31025_/S VGND VGND VPWR VPWR _31008_/A sky130_fd_sc_hd__mux2_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1059 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35815_ _35815_/CLK _35815_/D VGND VGND VPWR VPWR _35815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20972_ _20966_/X _20971_/X _20671_/X VGND VGND VPWR VPWR _20980_/C sky130_fd_sc_hd__o21ba_1
X_35746_ _35941_/CLK _35746_/D VGND VGND VPWR VPWR _35746_/Q sky130_fd_sc_hd__dfxtp_1
X_23760_ _23760_/A VGND VGND VPWR VPWR _32425_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32958_ _36095_/CLK _32958_/D VGND VGND VPWR VPWR _32958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22711_ _20577_/X _22709_/X _22710_/X _20587_/X VGND VGND VPWR VPWR _22711_/X sky130_fd_sc_hd__a22o_1
XFILLER_183_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31909_ _23283_/X _36154_/Q _31919_/S VGND VGND VPWR VPWR _31910_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23691_ _23691_/A VGND VGND VPWR VPWR _32394_/D sky130_fd_sc_hd__clkbuf_1
X_35677_ _35807_/CLK _35677_/D VGND VGND VPWR VPWR _35677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32889_ _32954_/CLK _32889_/D VGND VGND VPWR VPWR _32889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25430_ _25430_/A VGND VGND VPWR VPWR _33151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34628_ _35332_/CLK _34628_/D VGND VGND VPWR VPWR _34628_/Q sky130_fd_sc_hd__dfxtp_1
X_22642_ _32774_/Q _32710_/Q _32646_/Q _36102_/Q _22578_/X _22362_/X VGND VGND VPWR
+ VPWR _22642_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22573_ _22501_/X _22571_/X _22572_/X _22506_/X VGND VGND VPWR VPWR _22573_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25361_ _25361_/A VGND VGND VPWR VPWR _33118_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34559_ _35710_/CLK _34559_/D VGND VGND VPWR VPWR _34559_/Q sky130_fd_sc_hd__dfxtp_1
X_27100_ _26937_/X _33907_/Q _27104_/S VGND VGND VPWR VPWR _27101_/A sky130_fd_sc_hd__mux2_1
X_24312_ _32675_/Q _24311_/X _24336_/S VGND VGND VPWR VPWR _24313_/A sky130_fd_sc_hd__mux2_1
X_28080_ _28080_/A VGND VGND VPWR VPWR _34370_/D sky130_fd_sc_hd__clkbuf_1
X_21524_ _32486_/Q _32358_/Q _32038_/Q _36006_/Q _21523_/X _21311_/X VGND VGND VPWR
+ VPWR _21524_/X sky130_fd_sc_hd__mux4_1
X_25292_ _25292_/A VGND VGND VPWR VPWR _33086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27031_ _26835_/X _33874_/Q _27041_/S VGND VGND VPWR VPWR _27032_/A sky130_fd_sc_hd__mux2_1
X_36229_ _36232_/CLK _36229_/D VGND VGND VPWR VPWR _36229_/Q sky130_fd_sc_hd__dfxtp_1
X_24243_ _24243_/A VGND VGND VPWR VPWR _32653_/D sky130_fd_sc_hd__clkbuf_1
X_21455_ _32740_/Q _32676_/Q _32612_/Q _36068_/Q _21166_/X _21303_/X VGND VGND VPWR
+ VPWR _21455_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_336_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _36087_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_135_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20406_ _33032_/Q _32968_/Q _32904_/Q _32840_/Q _18280_/X _18283_/X VGND VGND VPWR
+ VPWR _20406_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24174_ _22972_/X _32620_/Q _24192_/S VGND VGND VPWR VPWR _24175_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21386_ _35810_/Q _32186_/Q _35682_/Q _35618_/Q _21207_/X _21208_/X VGND VGND VPWR
+ VPWR _21386_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20337_ _20201_/X _20335_/X _20336_/X _20206_/X VGND VGND VPWR VPWR _20337_/X sky130_fd_sc_hd__a22o_1
XFILLER_123_928 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23125_ _32154_/Q _23124_/X _23146_/S VGND VGND VPWR VPWR _23126_/A sky130_fd_sc_hd__mux2_1
X_28982_ _34798_/Q _24345_/X _28996_/S VGND VGND VPWR VPWR _28983_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23056_ input53/X VGND VGND VPWR VPWR _23056_/X sky130_fd_sc_hd__buf_4
X_27933_ _34301_/Q _24391_/X _27937_/S VGND VGND VPWR VPWR _27934_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20268_ _20264_/X _20267_/X _20167_/X VGND VGND VPWR VPWR _20269_/D sky130_fd_sc_hd__o21ba_1
XTAP_6025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22007_ _22003_/X _22006_/X _21728_/X VGND VGND VPWR VPWR _22039_/A sky130_fd_sc_hd__o21ba_1
XTAP_6069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27864_ _34268_/Q _24289_/X _27874_/S VGND VGND VPWR VPWR _27865_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20199_ _20199_/A _20199_/B _20199_/C _20199_/D VGND VGND VPWR VPWR _20200_/A sky130_fd_sc_hd__or4_1
XTAP_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26815_ _33803_/Q _24434_/X _26819_/S VGND VGND VPWR VPWR _26816_/A sky130_fd_sc_hd__mux2_1
XTAP_5368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29603_ _29603_/A VGND VGND VPWR VPWR _35061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27795_ _27795_/A VGND VGND VPWR VPWR _34235_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29534_ _29534_/A VGND VGND VPWR VPWR _35028_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26746_ _33770_/Q _24332_/X _26748_/S VGND VGND VPWR VPWR _26747_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23958_ _23056_/X _32519_/Q _23962_/S VGND VGND VPWR VPWR _23959_/A sky130_fd_sc_hd__mux2_1
XTAP_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_900 _26007_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_911 _27018_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_922 _27154_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22909_ _22909_/A VGND VGND VPWR VPWR _32023_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29465_ _23264_/X _34996_/Q _29467_/S VGND VGND VPWR VPWR _29466_/A sky130_fd_sc_hd__mux2_1
X_26677_ _25177_/X _33738_/Q _26683_/S VGND VGND VPWR VPWR _26678_/A sky130_fd_sc_hd__mux2_1
XTAP_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_933 _29247_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_944 _29517_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23889_ _22954_/X _32486_/Q _23899_/S VGND VGND VPWR VPWR _23890_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_955 _29787_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28416_ _28506_/S VGND VGND VPWR VPWR _28435_/S sky130_fd_sc_hd__clkbuf_8
X_16430_ _17842_/A VGND VGND VPWR VPWR _16430_/X sky130_fd_sc_hd__clkbuf_4
X_25628_ _25628_/A VGND VGND VPWR VPWR _33241_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_966 _31138_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29396_ _23102_/X _34963_/Q _29404_/S VGND VGND VPWR VPWR _29397_/A sky130_fd_sc_hd__mux2_1
XANTENNA_977 _17855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_988 _17796_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_999 _17957_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28347_ _34497_/Q _24404_/X _28363_/S VGND VGND VPWR VPWR _28348_/A sky130_fd_sc_hd__mux2_1
X_16361_ _17911_/A VGND VGND VPWR VPWR _16361_/X sky130_fd_sc_hd__buf_4
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25559_ _25559_/A VGND VGND VPWR VPWR _33210_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18100_ _17908_/X _18098_/X _18099_/X _17911_/X VGND VGND VPWR VPWR _18100_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19080_ _32482_/Q _32354_/Q _32034_/Q _36002_/Q _18870_/X _19011_/X VGND VGND VPWR
+ VPWR _19080_/X sky130_fd_sc_hd__mux4_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ _16288_/X _16289_/X _16290_/X _16291_/X VGND VGND VPWR VPWR _16292_/X sky130_fd_sc_hd__a22o_1
XFILLER_13_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28278_ _28278_/A VGND VGND VPWR VPWR _34464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18031_ _17860_/X _18029_/X _18030_/X _17865_/X VGND VGND VPWR VPWR _18031_/X sky130_fd_sc_hd__a22o_1
XFILLER_199_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27229_ _26928_/X _33968_/Q _27239_/S VGND VGND VPWR VPWR _27230_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_327_CLK clkbuf_6_44__f_CLK/X VGND VGND VPWR VPWR _35958_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_185_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30240_ _35363_/Q _29117_/X _30256_/S VGND VGND VPWR VPWR _30241_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30171_ _30171_/A VGND VGND VPWR VPWR _35330_/D sky130_fd_sc_hd__clkbuf_1
X_19982_ _19982_/A _19982_/B _19982_/C _19982_/D VGND VGND VPWR VPWR _19983_/A sky130_fd_sc_hd__or4_4
XFILLER_193_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18933_ _33246_/Q _36126_/Q _33118_/Q _33054_/Q _18652_/X _18653_/X VGND VGND VPWR
+ VPWR _18933_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1310 _17125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1321 input54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1332 _18360_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33930_ _35273_/CLK _33930_/D VGND VGND VPWR VPWR _33930_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1343 _22434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_1248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1354 _21728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18864_ _18796_/X _18862_/X _18863_/X _18799_/X VGND VGND VPWR VPWR _18864_/X sky130_fd_sc_hd__a22o_1
XTAP_6570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1365 _24304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1376 _26863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1387 _31408_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17815_ _17705_/X _17813_/X _17814_/X _17708_/X VGND VGND VPWR VPWR _17815_/X sky130_fd_sc_hd__a22o_1
X_33861_ _35780_/CLK _33861_/D VGND VGND VPWR VPWR _33861_/Q sky130_fd_sc_hd__dfxtp_1
X_18795_ _18789_/X _18792_/X _18793_/X _18794_/X VGND VGND VPWR VPWR _18795_/X sky130_fd_sc_hd__a22o_1
XTAP_5880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35600_ _35664_/CLK _35600_/D VGND VGND VPWR VPWR _35600_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17746_ _35325_/Q _35261_/Q _35197_/Q _32317_/Q _17712_/X _17713_/X VGND VGND VPWR
+ VPWR _17746_/X sky130_fd_sc_hd__mux4_1
X_32812_ _36080_/CLK _32812_/D VGND VGND VPWR VPWR _32812_/Q sky130_fd_sc_hd__dfxtp_1
X_33792_ _33793_/CLK _33792_/D VGND VGND VPWR VPWR _33792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35531_ _35979_/CLK _35531_/D VGND VGND VPWR VPWR _35531_/Q sky130_fd_sc_hd__dfxtp_1
X_17677_ _17502_/X _17675_/X _17676_/X _17505_/X VGND VGND VPWR VPWR _17677_/X sky130_fd_sc_hd__a22o_1
XFILLER_36_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32743_ _36072_/CLK _32743_/D VGND VGND VPWR VPWR _32743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19416_ _19101_/X _19414_/X _19415_/X _19106_/X VGND VGND VPWR VPWR _19416_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16628_ _33502_/Q _33438_/Q _33374_/Q _33310_/Q _16417_/X _16418_/X VGND VGND VPWR
+ VPWR _16628_/X sky130_fd_sc_hd__mux4_1
X_35462_ _35975_/CLK _35462_/D VGND VGND VPWR VPWR _35462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32674_ _36132_/CLK _32674_/D VGND VGND VPWR VPWR _32674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34413_ _35307_/CLK _34413_/D VGND VGND VPWR VPWR _34413_/Q sky130_fd_sc_hd__dfxtp_1
X_31625_ _31625_/A VGND VGND VPWR VPWR _36019_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19347_ _19347_/A VGND VGND VPWR VPWR _32105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16559_ _33756_/Q _33692_/Q _33628_/Q _33564_/Q _16490_/X _16491_/X VGND VGND VPWR
+ VPWR _16559_/X sky130_fd_sc_hd__mux4_1
X_35393_ _35909_/CLK _35393_/D VGND VGND VPWR VPWR _35393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31556_ _31556_/A VGND VGND VPWR VPWR _35986_/D sky130_fd_sc_hd__clkbuf_1
X_19278_ _33768_/Q _33704_/Q _33640_/Q _33576_/Q _19143_/X _19144_/X VGND VGND VPWR
+ VPWR _19278_/X sky130_fd_sc_hd__mux4_1
X_34344_ _34922_/CLK _34344_/D VGND VGND VPWR VPWR _34344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18229_ _35852_/Q _32232_/Q _35724_/Q _35660_/Q _15989_/X _15991_/X VGND VGND VPWR
+ VPWR _18229_/X sky130_fd_sc_hd__mux4_1
X_30507_ _30507_/A VGND VGND VPWR VPWR _35489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34275_ _34276_/CLK _34275_/D VGND VGND VPWR VPWR _34275_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_318_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _35831_/CLK sky130_fd_sc_hd__clkbuf_16
X_31487_ _23256_/X _35954_/Q _31493_/S VGND VGND VPWR VPWR _31488_/A sky130_fd_sc_hd__mux2_1
X_33226_ _35978_/CLK _33226_/D VGND VGND VPWR VPWR _33226_/Q sky130_fd_sc_hd__dfxtp_1
X_36014_ _36015_/CLK _36014_/D VGND VGND VPWR VPWR _36014_/Q sky130_fd_sc_hd__dfxtp_1
X_21240_ _21234_/X _21239_/X _21030_/X _21031_/X VGND VGND VPWR VPWR _21261_/B sky130_fd_sc_hd__o211a_1
X_30438_ _30438_/A VGND VGND VPWR VPWR _35456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33157_ _36100_/CLK _33157_/D VGND VGND VPWR VPWR _33157_/Q sky130_fd_sc_hd__dfxtp_1
X_21171_ _32476_/Q _32348_/Q _32028_/Q _35996_/Q _21170_/X _20958_/X VGND VGND VPWR
+ VPWR _21171_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30369_ _23142_/X _35424_/Q _30371_/S VGND VGND VPWR VPWR _30370_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20122_ _19807_/X _20120_/X _20121_/X _19812_/X VGND VGND VPWR VPWR _20122_/X sky130_fd_sc_hd__a22o_1
X_32108_ _35552_/CLK _32108_/D VGND VGND VPWR VPWR _32108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33088_ _36160_/CLK _33088_/D VGND VGND VPWR VPWR _33088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24930_ _24930_/A VGND VGND VPWR VPWR _32945_/D sky130_fd_sc_hd__clkbuf_1
X_20053_ _20053_/A VGND VGND VPWR VPWR _32125_/D sky130_fd_sc_hd__clkbuf_1
X_32039_ _35303_/CLK _32039_/D VGND VGND VPWR VPWR _32039_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24861_ _24861_/A VGND VGND VPWR VPWR _32912_/D sky130_fd_sc_hd__clkbuf_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26600_ _25063_/X _33701_/Q _26612_/S VGND VGND VPWR VPWR _26601_/A sky130_fd_sc_hd__mux2_1
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23812_ _23041_/X _32450_/Q _23826_/S VGND VGND VPWR VPWR _23813_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27580_ _27580_/A VGND VGND VPWR VPWR _34133_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24792_ _22985_/X _32880_/Q _24802_/S VGND VGND VPWR VPWR _24793_/A sky130_fd_sc_hd__mux2_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_207 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26531_ _25162_/X _33669_/Q _26539_/S VGND VGND VPWR VPWR _26532_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_218 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35729_ _35729_/CLK _35729_/D VGND VGND VPWR VPWR _35729_/Q sky130_fd_sc_hd__dfxtp_1
X_23743_ _23743_/A VGND VGND VPWR VPWR _32417_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20955_ _22506_/A VGND VGND VPWR VPWR _20955_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_229 _32136_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29250_ _29382_/S VGND VGND VPWR VPWR _29269_/S sky130_fd_sc_hd__buf_4
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26462_ _25060_/X _33636_/Q _26476_/S VGND VGND VPWR VPWR _26463_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23674_ _32386_/Q _23310_/X _23688_/S VGND VGND VPWR VPWR _23675_/A sky130_fd_sc_hd__mux2_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ _20626_/X _20882_/X _20885_/X _20637_/X VGND VGND VPWR VPWR _20886_/X sky130_fd_sc_hd__a22o_1
XFILLER_214_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28201_ _26965_/X _34428_/Q _28207_/S VGND VGND VPWR VPWR _28202_/A sky130_fd_sc_hd__mux2_1
X_25413_ _25119_/X _33143_/Q _25429_/S VGND VGND VPWR VPWR _25414_/A sky130_fd_sc_hd__mux2_1
X_22625_ _22621_/X _22624_/X _22453_/X VGND VGND VPWR VPWR _22633_/C sky130_fd_sc_hd__o21ba_1
XFILLER_201_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29181_ _29181_/A VGND VGND VPWR VPWR _34871_/D sky130_fd_sc_hd__clkbuf_1
X_26393_ _26393_/A VGND VGND VPWR VPWR _33603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28132_ _26863_/X _34395_/Q _28144_/S VGND VGND VPWR VPWR _28133_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25344_ _25344_/A VGND VGND VPWR VPWR _33110_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22556_ _22556_/A VGND VGND VPWR VPWR _22556_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_224_1288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28063_ _28063_/A VGND VGND VPWR VPWR _34362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21507_ _35045_/Q _34981_/Q _34917_/Q _34853_/Q _21403_/X _21404_/X VGND VGND VPWR
+ VPWR _21507_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_309_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _35257_/CLK sky130_fd_sc_hd__clkbuf_16
X_25275_ _25115_/X _33078_/Q _25293_/S VGND VGND VPWR VPWR _25276_/A sky130_fd_sc_hd__mux2_1
X_22487_ _22300_/X _22485_/X _22486_/X _22303_/X VGND VGND VPWR VPWR _22487_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27014_ input59/X VGND VGND VPWR VPWR _27014_/X sky130_fd_sc_hd__clkbuf_4
X_24226_ _23050_/X _32645_/Q _24234_/S VGND VGND VPWR VPWR _24227_/A sky130_fd_sc_hd__mux2_1
X_21438_ _21401_/X _21436_/X _21437_/X _21406_/X VGND VGND VPWR VPWR _21438_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24157_ _22948_/X _32612_/Q _24171_/S VGND VGND VPWR VPWR _24158_/A sky130_fd_sc_hd__mux2_1
X_21369_ _21089_/X _21367_/X _21368_/X _21094_/X VGND VGND VPWR VPWR _21369_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23108_ input62/X VGND VGND VPWR VPWR _23108_/X sky130_fd_sc_hd__buf_4
X_24088_ _23047_/X _32580_/Q _24098_/S VGND VGND VPWR VPWR _24089_/A sky130_fd_sc_hd__mux2_1
X_28965_ _34790_/Q _24320_/X _28975_/S VGND VGND VPWR VPWR _28966_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23039_ _23038_/X _32065_/Q _23063_/S VGND VGND VPWR VPWR _23040_/A sky130_fd_sc_hd__mux2_1
XTAP_5110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27916_ _34293_/Q _24366_/X _27916_/S VGND VGND VPWR VPWR _27917_/A sky130_fd_sc_hd__mux2_1
X_28896_ _28896_/A VGND VGND VPWR VPWR _34757_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27847_ _34260_/Q _24264_/X _27853_/S VGND VGND VPWR VPWR _27848_/A sky130_fd_sc_hd__mux2_1
XTAP_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _35833_/Q _32211_/Q _35705_/Q _35641_/Q _17313_/X _17314_/X VGND VGND VPWR
+ VPWR _17600_/X sky130_fd_sc_hd__mux4_1
XTAP_5198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18580_ _33236_/Q _36116_/Q _33108_/Q _33044_/Q _18320_/X _18321_/X VGND VGND VPWR
+ VPWR _18580_/X sky130_fd_sc_hd__mux4_1
XTAP_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27778_ _27778_/A VGND VGND VPWR VPWR _34227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _17527_/X _17530_/X _17489_/X _17490_/X VGND VGND VPWR VPWR _17546_/B sky130_fd_sc_hd__o211a_1
X_29517_ _23345_/X _35021_/Q _29517_/S VGND VGND VPWR VPWR _29518_/A sky130_fd_sc_hd__mux2_1
XTAP_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26729_ _26819_/S VGND VGND VPWR VPWR _26748_/S sky130_fd_sc_hd__buf_4
XTAP_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_730 _20980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_741 _21719_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_752 _22425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29448_ _29517_/S VGND VGND VPWR VPWR _29467_/S sky130_fd_sc_hd__buf_4
X_17462_ _17352_/X _17460_/X _17461_/X _17355_/X VGND VGND VPWR VPWR _17462_/X sky130_fd_sc_hd__a22o_1
XFILLER_229_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_763 _22500_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_774 _22538_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_785 _22634_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19201_ _18946_/X _19199_/X _19200_/X _18949_/X VGND VGND VPWR VPWR _19201_/X sky130_fd_sc_hd__a22o_1
X_16413_ _16413_/A VGND VGND VPWR VPWR _31959_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_796 _22844_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29379_ _29379_/A VGND VGND VPWR VPWR _34955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1041 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17393_ _35315_/Q _35251_/Q _35187_/Q _32307_/Q _17359_/X _17360_/X VGND VGND VPWR
+ VPWR _17393_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31410_ _31410_/A _31410_/B VGND VGND VPWR VPWR _31543_/S sky130_fd_sc_hd__nand2_8
XFILLER_198_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19132_ _19128_/X _19131_/X _19094_/X VGND VGND VPWR VPWR _19140_/C sky130_fd_sc_hd__o21ba_1
X_16344_ _16136_/X _16342_/X _16343_/X _16141_/X VGND VGND VPWR VPWR _16344_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32390_ _32518_/CLK _32390_/D VGND VGND VPWR VPWR _32390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19063_ _18748_/X _19061_/X _19062_/X _18753_/X VGND VGND VPWR VPWR _19063_/X sky130_fd_sc_hd__a22o_1
X_31341_ _31341_/A VGND VGND VPWR VPWR _35884_/D sky130_fd_sc_hd__clkbuf_1
X_16275_ _33492_/Q _33428_/Q _33364_/Q _33300_/Q _15998_/X _15999_/X VGND VGND VPWR
+ VPWR _16275_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18014_ _17761_/X _18012_/X _18013_/X _17767_/X VGND VGND VPWR VPWR _18014_/X sky130_fd_sc_hd__a22o_1
XFILLER_199_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34060_ _34060_/CLK _34060_/D VGND VGND VPWR VPWR _34060_/Q sky130_fd_sc_hd__dfxtp_1
X_31272_ _31272_/A VGND VGND VPWR VPWR _35852_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33011_ _35765_/CLK _33011_/D VGND VGND VPWR VPWR _33011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30223_ _35355_/Q _29092_/X _30235_/S VGND VGND VPWR VPWR _30224_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_1468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30154_ _30154_/A VGND VGND VPWR VPWR _35322_/D sky130_fd_sc_hd__clkbuf_1
X_19965_ _19961_/X _19964_/X _19789_/X _19790_/X VGND VGND VPWR VPWR _19982_/B sky130_fd_sc_hd__o211a_1
XFILLER_114_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18916_ _34781_/Q _34717_/Q _34653_/Q _34589_/Q _18882_/X _18883_/X VGND VGND VPWR
+ VPWR _18916_/X sky130_fd_sc_hd__mux4_1
XTAP_7090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34962_ _35026_/CLK _34962_/D VGND VGND VPWR VPWR _34962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30085_ _30085_/A VGND VGND VPWR VPWR _35289_/D sky130_fd_sc_hd__clkbuf_1
X_19896_ _32505_/Q _32377_/Q _32057_/Q _36025_/Q _19576_/X _19717_/X VGND VGND VPWR
+ VPWR _19896_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1140 _20201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1151 _20203_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1162 _22501_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_1468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33913_ _36154_/CLK _33913_/D VGND VGND VPWR VPWR _33913_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1173 _22453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18847_ _33179_/Q _32539_/Q _35931_/Q _35867_/Q _18668_/X _18669_/X VGND VGND VPWR
+ VPWR _18847_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34893_ _35021_/CLK _34893_/D VGND VGND VPWR VPWR _34893_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1184 _22217_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1195 _22932_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33844_ _35700_/CLK _33844_/D VGND VGND VPWR VPWR _33844_/Q sky130_fd_sc_hd__dfxtp_1
X_18778_ _18593_/X _18776_/X _18777_/X _18596_/X VGND VGND VPWR VPWR _18778_/X sky130_fd_sc_hd__a22o_1
XFILLER_227_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17729_ _17555_/X _17725_/X _17728_/X _17558_/X VGND VGND VPWR VPWR _17729_/X sky130_fd_sc_hd__a22o_1
X_30987_ _35717_/Q _29222_/X _30995_/S VGND VGND VPWR VPWR _30988_/A sky130_fd_sc_hd__mux2_1
X_33775_ _33775_/CLK _33775_/D VGND VGND VPWR VPWR _33775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35514_ _35578_/CLK _35514_/D VGND VGND VPWR VPWR _35514_/Q sky130_fd_sc_hd__dfxtp_1
X_20740_ _34256_/Q _34192_/Q _34128_/Q _34064_/Q _20605_/X _20607_/X VGND VGND VPWR
+ VPWR _20740_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32726_ _36055_/CLK _32726_/D VGND VGND VPWR VPWR _32726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20671_ _22453_/A VGND VGND VPWR VPWR _20671_/X sky130_fd_sc_hd__buf_2
XFILLER_23_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35445_ _36021_/CLK _35445_/D VGND VGND VPWR VPWR _35445_/Q sky130_fd_sc_hd__dfxtp_1
X_32657_ _36050_/CLK _32657_/D VGND VGND VPWR VPWR _32657_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_95_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _34775_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22410_ _35839_/Q _32218_/Q _35711_/Q _35647_/Q _22266_/X _22267_/X VGND VGND VPWR
+ VPWR _22410_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31608_ _31608_/A VGND VGND VPWR VPWR _36011_/D sky130_fd_sc_hd__clkbuf_1
X_32588_ _35532_/CLK _32588_/D VGND VGND VPWR VPWR _32588_/Q sky130_fd_sc_hd__dfxtp_1
X_23390_ _32254_/Q _23297_/X _23392_/S VGND VGND VPWR VPWR _23391_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35376_ _35952_/CLK _35376_/D VGND VGND VPWR VPWR _35376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34327_ _36196_/CLK _34327_/D VGND VGND VPWR VPWR _34327_/Q sky130_fd_sc_hd__dfxtp_1
X_22341_ _35581_/Q _35517_/Q _35453_/Q _35389_/Q _22203_/X _22204_/X VGND VGND VPWR
+ VPWR _22341_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31539_ _23339_/X _35979_/Q _31543_/S VGND VGND VPWR VPWR _31540_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22272_ _33211_/Q _32571_/Q _35963_/Q _35899_/Q _22027_/X _22028_/X VGND VGND VPWR
+ VPWR _22272_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_1445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25060_ input15/X VGND VGND VPWR VPWR _25060_/X sky130_fd_sc_hd__buf_2
X_34258_ _35789_/CLK _34258_/D VGND VGND VPWR VPWR _34258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24011_ _24011_/A VGND VGND VPWR VPWR _32543_/D sky130_fd_sc_hd__clkbuf_1
X_21223_ _21223_/A _21223_/B _21223_/C _21223_/D VGND VGND VPWR VPWR _21224_/A sky130_fd_sc_hd__or4_2
X_33209_ _36027_/CLK _33209_/D VGND VGND VPWR VPWR _33209_/Q sky130_fd_sc_hd__dfxtp_1
X_34189_ _34317_/CLK _34189_/D VGND VGND VPWR VPWR _34189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21154_ _35035_/Q _34971_/Q _34907_/Q _34843_/Q _21050_/X _21051_/X VGND VGND VPWR
+ VPWR _21154_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20105_ _20061_/X _20103_/X _20104_/X _20067_/X VGND VGND VPWR VPWR _20105_/X sky130_fd_sc_hd__a22o_1
X_28750_ _26977_/X _34688_/Q _28768_/S VGND VGND VPWR VPWR _28751_/A sky130_fd_sc_hd__mux2_1
X_25962_ _25119_/X _33399_/Q _25978_/S VGND VGND VPWR VPWR _25963_/A sky130_fd_sc_hd__mux2_1
X_21085_ _21048_/X _21083_/X _21084_/X _21053_/X VGND VGND VPWR VPWR _21085_/X sky130_fd_sc_hd__a22o_1
XFILLER_154_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27701_ _27701_/A VGND VGND VPWR VPWR _34190_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20036_ _19716_/X _20034_/X _20035_/X _19720_/X VGND VGND VPWR VPWR _20036_/X sky130_fd_sc_hd__a22o_1
XFILLER_63_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24913_ _24913_/A VGND VGND VPWR VPWR _32937_/D sky130_fd_sc_hd__clkbuf_1
X_28681_ _28681_/A VGND VGND VPWR VPWR _34655_/D sky130_fd_sc_hd__clkbuf_1
X_25893_ _25893_/A VGND VGND VPWR VPWR _33366_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27632_ _34158_/Q _24345_/X _27646_/S VGND VGND VPWR VPWR _27633_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24844_ _23062_/X _32905_/Q _24844_/S VGND VGND VPWR VPWR _24845_/A sky130_fd_sc_hd__mux2_1
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27563_ _27833_/A _30870_/B VGND VGND VPWR VPWR _27696_/S sky130_fd_sc_hd__nor2_8
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24775_ _22960_/X _32872_/Q _24781_/S VGND VGND VPWR VPWR _24776_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21987_ _21947_/X _21985_/X _21986_/X _21950_/X VGND VGND VPWR VPWR _21987_/X sky130_fd_sc_hd__a22o_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29302_ _29302_/A VGND VGND VPWR VPWR _34918_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26514_ _25137_/X _33661_/Q _26518_/S VGND VGND VPWR VPWR _26515_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23726_ _22914_/X _32409_/Q _23742_/S VGND VGND VPWR VPWR _23727_/A sky130_fd_sc_hd__mux2_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20938_ _20687_/X _20936_/X _20937_/X _20697_/X VGND VGND VPWR VPWR _20938_/X sky130_fd_sc_hd__a22o_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_892 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27494_ _27494_/A VGND VGND VPWR VPWR _34093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29233_ _29233_/A VGND VGND VPWR VPWR _34888_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26445_ _25035_/X _33628_/Q _26455_/S VGND VGND VPWR VPWR _26446_/A sky130_fd_sc_hd__mux2_1
X_23657_ _32378_/Q _23283_/X _23667_/S VGND VGND VPWR VPWR _23658_/A sky130_fd_sc_hd__mux2_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20869_ _20865_/X _20868_/X _20700_/X VGND VGND VPWR VPWR _20870_/D sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_86_CLK clkbuf_leaf_87_CLK/A VGND VGND VPWR VPWR _35799_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22608_ _33541_/Q _33477_/Q _33413_/Q _33349_/Q _22429_/X _22430_/X VGND VGND VPWR
+ VPWR _22608_/X sky130_fd_sc_hd__mux4_1
XFILLER_161_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29164_ _34866_/Q _29163_/X _29173_/S VGND VGND VPWR VPWR _29165_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26376_ _26376_/A VGND VGND VPWR VPWR _33595_/D sky130_fd_sc_hd__clkbuf_1
X_23588_ _32345_/Q _23121_/X _23604_/S VGND VGND VPWR VPWR _23589_/A sky130_fd_sc_hd__mux2_1
X_28115_ _26838_/X _34387_/Q _28123_/S VGND VGND VPWR VPWR _28116_/A sky130_fd_sc_hd__mux2_1
X_25327_ _24989_/X _33102_/Q _25345_/S VGND VGND VPWR VPWR _25328_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22539_ _33795_/Q _33731_/Q _33667_/Q _33603_/Q _22502_/X _22503_/X VGND VGND VPWR
+ VPWR _22539_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29095_ input6/X VGND VGND VPWR VPWR _29095_/X sky130_fd_sc_hd__buf_4
XFILLER_185_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16060_ _17847_/A VGND VGND VPWR VPWR _16060_/X sky130_fd_sc_hd__buf_6
XFILLER_194_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28046_ _28046_/A VGND VGND VPWR VPWR _34354_/D sky130_fd_sc_hd__clkbuf_1
X_25258_ _25091_/X _33070_/Q _25272_/S VGND VGND VPWR VPWR _25259_/A sky130_fd_sc_hd__mux2_1
X_24209_ _23025_/X _32637_/Q _24213_/S VGND VGND VPWR VPWR _24210_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25189_ _30735_/B _31815_/B VGND VGND VPWR VPWR _25322_/S sky130_fd_sc_hd__nand2_8
XFILLER_185_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29997_ _35248_/Q _29157_/X _30007_/S VGND VGND VPWR VPWR _29998_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19750_ _32757_/Q _32693_/Q _32629_/Q _36085_/Q _19572_/X _19709_/X VGND VGND VPWR
+ VPWR _19750_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16962_ _35815_/Q _32191_/Q _35687_/Q _35623_/Q _16960_/X _16961_/X VGND VGND VPWR
+ VPWR _16962_/X sky130_fd_sc_hd__mux4_1
X_28948_ _34782_/Q _24295_/X _28954_/S VGND VGND VPWR VPWR _28949_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _35098_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_46_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18701_ _35543_/Q _35479_/Q _35415_/Q _35351_/Q _18491_/X _18492_/X VGND VGND VPWR
+ VPWR _18701_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19681_ _32499_/Q _32371_/Q _32051_/Q _36019_/Q _19576_/X _19364_/X VGND VGND VPWR
+ VPWR _19681_/X sky130_fd_sc_hd__mux4_1
X_16893_ _16889_/X _16892_/X _16783_/X _16784_/X VGND VGND VPWR VPWR _16910_/B sky130_fd_sc_hd__o211a_1
XFILLER_77_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28879_ _28879_/A VGND VGND VPWR VPWR _34749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18632_ _18628_/X _18631_/X _18371_/X VGND VGND VPWR VPWR _18640_/C sky130_fd_sc_hd__o21ba_1
X_30910_ _30910_/A VGND VGND VPWR VPWR _35680_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31890_ _23253_/X _36145_/Q _31898_/S VGND VGND VPWR VPWR _31891_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30841_ _30868_/S VGND VGND VPWR VPWR _30860_/S sky130_fd_sc_hd__buf_4
XTAP_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18563_ _34771_/Q _34707_/Q _34643_/Q _34579_/Q _18529_/X _18530_/X VGND VGND VPWR
+ VPWR _18563_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17514_ _17867_/A VGND VGND VPWR VPWR _17514_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18494_ _33169_/Q _32529_/Q _35921_/Q _35857_/Q _18363_/X _18365_/X VGND VGND VPWR
+ VPWR _18494_/X sky130_fd_sc_hd__mux4_1
X_33560_ _35671_/CLK _33560_/D VGND VGND VPWR VPWR _33560_/Q sky130_fd_sc_hd__dfxtp_1
X_30772_ _23139_/X _35615_/Q _30776_/S VGND VGND VPWR VPWR _30773_/A sky130_fd_sc_hd__mux2_1
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_560 _20146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_571 _20147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32511_ _36033_/CLK _32511_/D VGND VGND VPWR VPWR _32511_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_582 _19449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17445_ _17195_/X _17441_/X _17444_/X _17200_/X VGND VGND VPWR VPWR _17445_/X sky130_fd_sc_hd__a22o_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33491_ _36237_/CLK _33491_/D VGND VGND VPWR VPWR _33491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_593 _19459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_77_CLK clkbuf_leaf_80_CLK/A VGND VGND VPWR VPWR _35921_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_60_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32442_ _35771_/CLK _32442_/D VGND VGND VPWR VPWR _32442_/Q sky130_fd_sc_hd__dfxtp_1
X_35230_ _35294_/CLK _35230_/D VGND VGND VPWR VPWR _35230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17376_ _17202_/X _17372_/X _17375_/X _17205_/X VGND VGND VPWR VPWR _17376_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16327_ _35733_/Q _35093_/Q _34453_/Q _33813_/Q _16049_/X _16051_/X VGND VGND VPWR
+ VPWR _16327_/X sky130_fd_sc_hd__mux4_1
X_19115_ _33507_/Q _33443_/Q _33379_/Q _33315_/Q _19070_/X _19071_/X VGND VGND VPWR
+ VPWR _19115_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35161_ _36201_/CLK _35161_/D VGND VGND VPWR VPWR _35161_/Q sky130_fd_sc_hd__dfxtp_1
X_32373_ _36085_/CLK _32373_/D VGND VGND VPWR VPWR _32373_/Q sky130_fd_sc_hd__dfxtp_1
X_34112_ _36165_/CLK _34112_/D VGND VGND VPWR VPWR _34112_/Q sky130_fd_sc_hd__dfxtp_1
X_31324_ _31324_/A VGND VGND VPWR VPWR _35876_/D sky130_fd_sc_hd__clkbuf_1
X_19046_ _19002_/X _19044_/X _19045_/X _19008_/X VGND VGND VPWR VPWR _19046_/X sky130_fd_sc_hd__a22o_1
X_16258_ _16044_/X _16256_/X _16257_/X _16054_/X VGND VGND VPWR VPWR _16258_/X sky130_fd_sc_hd__a22o_1
X_35092_ _35730_/CLK _35092_/D VGND VGND VPWR VPWR _35092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput203 _36228_/Q VGND VGND VPWR VPWR D2[54] sky130_fd_sc_hd__buf_2
XFILLER_86_1221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31255_ _35844_/Q input50/X _31265_/S VGND VGND VPWR VPWR _31256_/A sky130_fd_sc_hd__mux2_1
X_34043_ _34171_/CLK _34043_/D VGND VGND VPWR VPWR _34043_/Q sky130_fd_sc_hd__dfxtp_1
X_16189_ _35729_/Q _35089_/Q _34449_/Q _33809_/Q _16049_/X _16051_/X VGND VGND VPWR
+ VPWR _16189_/X sky130_fd_sc_hd__mux4_1
Xoutput214 _36180_/Q VGND VGND VPWR VPWR D2[6] sky130_fd_sc_hd__buf_2
Xoutput225 _32094_/Q VGND VGND VPWR VPWR D3[16] sky130_fd_sc_hd__buf_2
Xoutput236 _32104_/Q VGND VGND VPWR VPWR D3[26] sky130_fd_sc_hd__buf_2
X_30206_ _35347_/Q _29067_/X _30214_/S VGND VGND VPWR VPWR _30207_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput247 _32114_/Q VGND VGND VPWR VPWR D3[36] sky130_fd_sc_hd__buf_2
XFILLER_177_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput258 _32124_/Q VGND VGND VPWR VPWR D3[46] sky130_fd_sc_hd__buf_2
X_31186_ _35811_/Q input14/X _31202_/S VGND VGND VPWR VPWR _31187_/A sky130_fd_sc_hd__mux2_1
Xoutput269 _32134_/Q VGND VGND VPWR VPWR D3[56] sky130_fd_sc_hd__buf_2
XFILLER_138_1377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30137_ _30137_/A VGND VGND VPWR VPWR _35314_/D sky130_fd_sc_hd__clkbuf_1
X_19948_ _19807_/X _19946_/X _19947_/X _19812_/X VGND VGND VPWR VPWR _19948_/X sky130_fd_sc_hd__a22o_1
X_35994_ _35994_/CLK _35994_/D VGND VGND VPWR VPWR _35994_/Q sky130_fd_sc_hd__dfxtp_1
X_34945_ _35075_/CLK _34945_/D VGND VGND VPWR VPWR _34945_/Q sky130_fd_sc_hd__dfxtp_1
X_30068_ _30068_/A VGND VGND VPWR VPWR _35281_/D sky130_fd_sc_hd__clkbuf_1
X_19879_ _20232_/A VGND VGND VPWR VPWR _19879_/X sky130_fd_sc_hd__buf_4
XFILLER_67_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21910_ _33009_/Q _32945_/Q _32881_/Q _32817_/Q _21589_/X _21590_/X VGND VGND VPWR
+ VPWR _21910_/X sky130_fd_sc_hd__mux4_1
XFILLER_244_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22890_ _22889_/X _32017_/Q _22908_/S VGND VGND VPWR VPWR _22891_/A sky130_fd_sc_hd__mux2_1
X_34876_ _35515_/CLK _34876_/D VGND VGND VPWR VPWR _34876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21841_ _33263_/Q _36143_/Q _33135_/Q _33071_/Q _21658_/X _21659_/X VGND VGND VPWR
+ VPWR _21841_/X sky130_fd_sc_hd__mux4_1
X_33827_ _35876_/CLK _33827_/D VGND VGND VPWR VPWR _33827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24560_ _24560_/A VGND VGND VPWR VPWR _32772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21772_ _32749_/Q _32685_/Q _32621_/Q _36077_/Q _21519_/X _21656_/X VGND VGND VPWR
+ VPWR _21772_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33758_ _34080_/CLK _33758_/D VGND VGND VPWR VPWR _33758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23511_ _23559_/S VGND VGND VPWR VPWR _23530_/S sky130_fd_sc_hd__buf_4
XFILLER_93_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20723_ _35535_/Q _35471_/Q _35407_/Q _35343_/Q _20658_/X _20660_/X VGND VGND VPWR
+ VPWR _20723_/X sky130_fd_sc_hd__mux4_1
X_32709_ _36100_/CLK _32709_/D VGND VGND VPWR VPWR _32709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24491_ _24491_/A VGND VGND VPWR VPWR _32739_/D sky130_fd_sc_hd__clkbuf_1
X_33689_ _35799_/CLK _33689_/D VGND VGND VPWR VPWR _33689_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_68_CLK clkbuf_leaf_73_CLK/A VGND VGND VPWR VPWR _36055_/CLK sky130_fd_sc_hd__clkbuf_16
X_26230_ _25115_/X _33526_/Q _26248_/S VGND VGND VPWR VPWR _26231_/A sky130_fd_sc_hd__mux2_1
X_23442_ _22901_/X _32277_/Q _23446_/S VGND VGND VPWR VPWR _23443_/A sky130_fd_sc_hd__mux2_1
X_35428_ _35555_/CLK _35428_/D VGND VGND VPWR VPWR _35428_/Q sky130_fd_sc_hd__dfxtp_1
X_20654_ _22458_/A VGND VGND VPWR VPWR _20654_/X sky130_fd_sc_hd__buf_4
XFILLER_23_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26161_ _26161_/A VGND VGND VPWR VPWR _33493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20585_ input73/X input74/X VGND VGND VPWR VPWR _22367_/A sky130_fd_sc_hd__nor2_4
X_23373_ _23421_/S VGND VGND VPWR VPWR _23392_/S sky130_fd_sc_hd__buf_4
X_35359_ _35937_/CLK _35359_/D VGND VGND VPWR VPWR _35359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25112_ input33/X VGND VGND VPWR VPWR _25112_/X sky130_fd_sc_hd__buf_2
XFILLER_99_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22324_ _22148_/X _22322_/X _22323_/X _22153_/X VGND VGND VPWR VPWR _22324_/X sky130_fd_sc_hd__a22o_1
X_26092_ _25112_/X _33461_/Q _26092_/S VGND VGND VPWR VPWR _26093_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_6_34__f_CLK clkbuf_5_17_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_34__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_152_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29920_ _35212_/Q _29243_/X _29922_/S VGND VGND VPWR VPWR _29921_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25043_ _25043_/A VGND VGND VPWR VPWR _32990_/D sky130_fd_sc_hd__clkbuf_1
X_22255_ _33531_/Q _33467_/Q _33403_/Q _33339_/Q _22076_/X _22077_/X VGND VGND VPWR
+ VPWR _22255_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21206_ _21202_/X _21205_/X _21030_/X _21031_/X VGND VGND VPWR VPWR _21223_/B sky130_fd_sc_hd__o211a_1
XFILLER_195_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22186_ _33785_/Q _33721_/Q _33657_/Q _33593_/Q _22149_/X _22150_/X VGND VGND VPWR
+ VPWR _22186_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29851_ _35179_/Q _29141_/X _29851_/S VGND VGND VPWR VPWR _29852_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28802_ _28802_/A VGND VGND VPWR VPWR _34712_/D sky130_fd_sc_hd__clkbuf_1
X_21137_ _32475_/Q _32347_/Q _32027_/Q _35995_/Q _20817_/X _20958_/X VGND VGND VPWR
+ VPWR _21137_/X sky130_fd_sc_hd__mux4_1
X_29782_ _29782_/A VGND VGND VPWR VPWR _35146_/D sky130_fd_sc_hd__clkbuf_1
X_26994_ _26993_/X _33861_/Q _27006_/S VGND VGND VPWR VPWR _26995_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21068_ _20949_/X _21066_/X _21067_/X _20955_/X VGND VGND VPWR VPWR _21068_/X sky130_fd_sc_hd__a22o_1
X_25945_ _25094_/X _33391_/Q _25957_/S VGND VGND VPWR VPWR _25946_/A sky130_fd_sc_hd__mux2_1
X_28733_ _26953_/X _34680_/Q _28747_/S VGND VGND VPWR VPWR _28734_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20019_ _20015_/X _20018_/X _19814_/X VGND VGND VPWR VPWR _20020_/D sky130_fd_sc_hd__o21ba_1
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28664_ _28664_/A VGND VGND VPWR VPWR _34647_/D sky130_fd_sc_hd__clkbuf_1
X_25876_ _24989_/X _33358_/Q _25894_/S VGND VGND VPWR VPWR _25877_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24827_ _24827_/A VGND VGND VPWR VPWR _32896_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27615_ _34150_/Q _24320_/X _27625_/S VGND VGND VPWR VPWR _27616_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28595_ _28595_/A VGND VGND VPWR VPWR _34614_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27546_ _27546_/A VGND VGND VPWR VPWR _34118_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24758_ _22935_/X _32864_/Q _24760_/S VGND VGND VPWR VPWR _24759_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23709_ _22889_/X _32401_/Q _23721_/S VGND VGND VPWR VPWR _23710_/A sky130_fd_sc_hd__mux2_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27477_ _27477_/A VGND VGND VPWR VPWR _34085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24689_ _23034_/X _32832_/Q _24707_/S VGND VGND VPWR VPWR _24690_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_59_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _34277_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_203_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17230_ _17224_/X _17229_/X _17161_/X VGND VGND VPWR VPWR _17231_/D sky130_fd_sc_hd__o21ba_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26428_ _25010_/X _33620_/Q _26434_/S VGND VGND VPWR VPWR _26429_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29216_ input49/X VGND VGND VPWR VPWR _29216_/X sky130_fd_sc_hd__buf_4
XFILLER_187_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29147_ _29147_/A VGND VGND VPWR VPWR _34860_/D sky130_fd_sc_hd__clkbuf_1
X_17161_ _17867_/A VGND VGND VPWR VPWR _17161_/X sky130_fd_sc_hd__clkbuf_4
X_26359_ _26359_/A VGND VGND VPWR VPWR _33587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16112_ _16106_/X _16111_/X _16011_/X VGND VGND VPWR VPWR _16134_/A sky130_fd_sc_hd__o21ba_1
XFILLER_31_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29078_ _29078_/A VGND VGND VPWR VPWR _34838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17092_ _16842_/X _17088_/X _17091_/X _16847_/X VGND VGND VPWR VPWR _17092_/X sky130_fd_sc_hd__a22o_1
XFILLER_196_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16043_ _16024_/X _16038_/X _16040_/X _16042_/X VGND VGND VPWR VPWR _16102_/B sky130_fd_sc_hd__o211a_1
XFILLER_129_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28029_ _28029_/A VGND VGND VPWR VPWR _34346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31040_ _35742_/Q _29101_/X _31046_/S VGND VGND VPWR VPWR _31041_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19802_ _20155_/A VGND VGND VPWR VPWR _19802_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17994_ _17994_/A VGND VGND VPWR VPWR _17994_/X sky130_fd_sc_hd__buf_6
XFILLER_96_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19733_ _35316_/Q _35252_/Q _35188_/Q _32308_/Q _19659_/X _19660_/X VGND VGND VPWR
+ VPWR _19733_/X sky130_fd_sc_hd__mux4_1
X_16945_ _16945_/A VGND VGND VPWR VPWR _31974_/D sky130_fd_sc_hd__clkbuf_1
X_32991_ _36062_/CLK _32991_/D VGND VGND VPWR VPWR _32991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34730_ _34794_/CLK _34730_/D VGND VGND VPWR VPWR _34730_/Q sky130_fd_sc_hd__dfxtp_1
X_31942_ _23336_/X _36170_/Q _31948_/S VGND VGND VPWR VPWR _31943_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19664_ _35058_/Q _34994_/Q _34930_/Q _34866_/Q _19456_/X _19457_/X VGND VGND VPWR
+ VPWR _19664_/X sky130_fd_sc_hd__mux4_1
X_16876_ _16801_/X _16874_/X _16875_/X _16806_/X VGND VGND VPWR VPWR _16876_/X sky130_fd_sc_hd__a22o_1
XFILLER_49_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18615_ _20147_/A VGND VGND VPWR VPWR _18615_/X sky130_fd_sc_hd__clkbuf_8
XTAP_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34661_ _36001_/CLK _34661_/D VGND VGND VPWR VPWR _34661_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19595_ _19454_/X _19593_/X _19594_/X _19459_/X VGND VGND VPWR VPWR _19595_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31873_ _23228_/X _36137_/Q _31877_/S VGND VGND VPWR VPWR _31874_/A sky130_fd_sc_hd__mux2_1
X_33612_ _34124_/CLK _33612_/D VGND VGND VPWR VPWR _33612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18546_ _18542_/X _18545_/X _18311_/X VGND VGND VPWR VPWR _18570_/A sky130_fd_sc_hd__o21ba_1
X_30824_ _30824_/A VGND VGND VPWR VPWR _35639_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34592_ _34782_/CLK _34592_/D VGND VGND VPWR VPWR _34592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33543_ _33544_/CLK _33543_/D VGND VGND VPWR VPWR _33543_/Q sky130_fd_sc_hd__dfxtp_1
X_18477_ _33489_/Q _33425_/Q _33361_/Q _33297_/Q _18298_/X _18299_/X VGND VGND VPWR
+ VPWR _18477_/X sky130_fd_sc_hd__mux4_1
X_30755_ _23114_/X _35607_/Q _30755_/S VGND VGND VPWR VPWR _30756_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_390 _36209_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17428_ _17932_/A VGND VGND VPWR VPWR _17428_/X sky130_fd_sc_hd__buf_4
X_33474_ _34050_/CLK _33474_/D VGND VGND VPWR VPWR _33474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30686_ _35574_/Q _29175_/X _30704_/S VGND VGND VPWR VPWR _30687_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35213_ _35277_/CLK _35213_/D VGND VGND VPWR VPWR _35213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32425_ _35050_/CLK _32425_/D VGND VGND VPWR VPWR _32425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36193_ _36200_/CLK _36193_/D VGND VGND VPWR VPWR _36193_/Q sky130_fd_sc_hd__dfxtp_1
X_17359_ _17712_/A VGND VGND VPWR VPWR _17359_/X sky130_fd_sc_hd__buf_6
XFILLER_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35144_ _35784_/CLK _35144_/D VGND VGND VPWR VPWR _35144_/Q sky130_fd_sc_hd__dfxtp_1
X_20370_ _20208_/X _20368_/X _20369_/X _20211_/X VGND VGND VPWR VPWR _20370_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32356_ _36004_/CLK _32356_/D VGND VGND VPWR VPWR _32356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19029_ _34528_/Q _32416_/Q _34400_/Q _34336_/Q _18819_/X _18820_/X VGND VGND VPWR
+ VPWR _19029_/X sky130_fd_sc_hd__mux4_1
X_31307_ _31307_/A VGND VGND VPWR VPWR _35868_/D sky130_fd_sc_hd__clkbuf_1
X_35075_ _35075_/CLK _35075_/D VGND VGND VPWR VPWR _35075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32287_ _34782_/CLK _32287_/D VGND VGND VPWR VPWR _32287_/Q sky130_fd_sc_hd__dfxtp_1
X_22040_ _22040_/A VGND VGND VPWR VPWR _36212_/D sky130_fd_sc_hd__buf_6
X_31238_ _35836_/Q input41/X _31244_/S VGND VGND VPWR VPWR _31239_/A sky130_fd_sc_hd__mux2_1
X_34026_ _34283_/CLK _34026_/D VGND VGND VPWR VPWR _34026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31169_ _35803_/Q input5/X _31181_/S VGND VGND VPWR VPWR _31170_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35977_ _35977_/CLK _35977_/D VGND VGND VPWR VPWR _35977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23991_ _22904_/X _32534_/Q _23993_/S VGND VGND VPWR VPWR _23992_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25730_ _25730_/A VGND VGND VPWR VPWR _33290_/D sky130_fd_sc_hd__clkbuf_1
X_34928_ _35954_/CLK _34928_/D VGND VGND VPWR VPWR _34928_/Q sky130_fd_sc_hd__dfxtp_1
X_22942_ _23075_/S VGND VGND VPWR VPWR _22970_/S sky130_fd_sc_hd__buf_4
XFILLER_28_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25661_ _25661_/A VGND VGND VPWR VPWR _33257_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22873_ _22873_/A _22873_/B _22873_/C _22873_/D VGND VGND VPWR VPWR _22874_/A sky130_fd_sc_hd__or4_4
XFILLER_216_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34859_ _34859_/CLK _34859_/D VGND VGND VPWR VPWR _34859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27400_ _34049_/Q _24404_/X _27416_/S VGND VGND VPWR VPWR _27401_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24612_ _24612_/A VGND VGND VPWR VPWR _32795_/D sky130_fd_sc_hd__clkbuf_1
X_28380_ _28380_/A VGND VGND VPWR VPWR _34512_/D sky130_fd_sc_hd__clkbuf_1
X_21824_ _21749_/X _21822_/X _21823_/X _21752_/X VGND VGND VPWR VPWR _21824_/X sky130_fd_sc_hd__a22o_1
X_25592_ _25592_/A VGND VGND VPWR VPWR _33226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27331_ _27331_/A VGND VGND VPWR VPWR _34016_/D sky130_fd_sc_hd__clkbuf_1
X_24543_ _24543_/A VGND VGND VPWR VPWR _32764_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21755_ _34540_/Q _32428_/Q _34412_/Q _34348_/Q _21472_/X _21473_/X VGND VGND VPWR
+ VPWR _21755_/X sky130_fd_sc_hd__mux4_1
XFILLER_240_952 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20706_ _20577_/X _20704_/X _20705_/X _20587_/X VGND VGND VPWR VPWR _20706_/X sky130_fd_sc_hd__a22o_1
X_27262_ _27289_/S VGND VGND VPWR VPWR _27281_/S sky130_fd_sc_hd__buf_4
X_24474_ _24474_/A VGND VGND VPWR VPWR _32731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21686_ _21686_/A _21686_/B _21686_/C _21686_/D VGND VGND VPWR VPWR _21687_/A sky130_fd_sc_hd__or4_4
XFILLER_180_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29001_ _34807_/Q _24373_/X _29017_/S VGND VGND VPWR VPWR _29002_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26213_ _25091_/X _33518_/Q _26227_/S VGND VGND VPWR VPWR _26214_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23425_ _26549_/C _31680_/A VGND VGND VPWR VPWR _30735_/B sky130_fd_sc_hd__nor2_8
X_20637_ _22511_/A VGND VGND VPWR VPWR _20637_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_123_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27193_ _26875_/X _33951_/Q _27197_/S VGND VGND VPWR VPWR _27194_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26144_ _28373_/B _26685_/B VGND VGND VPWR VPWR _26277_/S sky130_fd_sc_hd__nand2_8
XFILLER_165_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23356_ _23356_/A VGND VGND VPWR VPWR _32237_/D sky130_fd_sc_hd__clkbuf_1
X_20568_ _18344_/X _20566_/X _20567_/X _18354_/X VGND VGND VPWR VPWR _20568_/X sky130_fd_sc_hd__a22o_1
XFILLER_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_926 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22307_ _33212_/Q _32572_/Q _35964_/Q _35900_/Q _22027_/X _22028_/X VGND VGND VPWR
+ VPWR _22307_/X sky130_fd_sc_hd__mux4_1
X_26075_ _26075_/A VGND VGND VPWR VPWR _33452_/D sky130_fd_sc_hd__clkbuf_1
X_23287_ _32213_/Q _23286_/X _23301_/S VGND VGND VPWR VPWR _23288_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20499_ _35851_/Q _32231_/Q _35723_/Q _35659_/Q _18289_/X _18291_/X VGND VGND VPWR
+ VPWR _20499_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29903_ _29903_/A VGND VGND VPWR VPWR _35203_/D sky130_fd_sc_hd__clkbuf_1
X_25026_ input3/X VGND VGND VPWR VPWR _25026_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22238_ _33210_/Q _32570_/Q _35962_/Q _35898_/Q _22027_/X _22028_/X VGND VGND VPWR
+ VPWR _22238_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29834_ _29834_/A VGND VGND VPWR VPWR _35170_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22169_ _35768_/Q _35128_/Q _34488_/Q _33848_/Q _22093_/X _22094_/X VGND VGND VPWR
+ VPWR _22169_/X sky130_fd_sc_hd__mux4_1
XTAP_6955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29765_ _35138_/Q _29213_/X _29779_/S VGND VGND VPWR VPWR _29766_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26977_ input46/X VGND VGND VPWR VPWR _26977_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_121_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16730_ _35040_/Q _34976_/Q _34912_/Q _34848_/Q _16450_/X _16451_/X VGND VGND VPWR
+ VPWR _16730_/X sky130_fd_sc_hd__mux4_1
X_28716_ _26928_/X _34672_/Q _28726_/S VGND VGND VPWR VPWR _28717_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25928_ _25069_/X _33383_/Q _25936_/S VGND VGND VPWR VPWR _25929_/A sky130_fd_sc_hd__mux2_1
X_29696_ _29696_/A VGND VGND VPWR VPWR _35105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16661_ _16661_/A _16661_/B _16661_/C _16661_/D VGND VGND VPWR VPWR _16662_/A sky130_fd_sc_hd__or4_1
XFILLER_235_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25859_ _25859_/A VGND VGND VPWR VPWR _33350_/D sky130_fd_sc_hd__clkbuf_1
X_28647_ _26826_/X _34639_/Q _28663_/S VGND VGND VPWR VPWR _28648_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18400_ _20167_/A VGND VGND VPWR VPWR _18400_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_74_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16592_ _16592_/A VGND VGND VPWR VPWR _31964_/D sky130_fd_sc_hd__clkbuf_1
X_19380_ _35306_/Q _35242_/Q _35178_/Q _32298_/Q _19306_/X _19307_/X VGND VGND VPWR
+ VPWR _19380_/X sky130_fd_sc_hd__mux4_1
X_28578_ _28578_/A VGND VGND VPWR VPWR _34606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18331_ _32462_/Q _32334_/Q _32014_/Q _35982_/Q _18328_/X _20163_/A VGND VGND VPWR
+ VPWR _18331_/X sky130_fd_sc_hd__mux4_1
X_27529_ _27529_/A VGND VGND VPWR VPWR _34110_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18262_ _35597_/Q _35533_/Q _35469_/Q _35405_/Q _16005_/X _16007_/X VGND VGND VPWR
+ VPWR _18262_/X sky130_fd_sc_hd__mux4_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30540_ _23253_/X _35505_/Q _30548_/S VGND VGND VPWR VPWR _30541_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17213_ _17063_/X _17211_/X _17212_/X _17067_/X VGND VGND VPWR VPWR _17213_/X sky130_fd_sc_hd__a22o_1
XFILLER_202_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18193_ _33291_/Q _36171_/Q _33163_/Q _33099_/Q _16028_/X _17157_/A VGND VGND VPWR
+ VPWR _18193_/X sky130_fd_sc_hd__mux4_1
X_30471_ _23093_/X _35472_/Q _30485_/S VGND VGND VPWR VPWR _30472_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32210_ _35833_/CLK _32210_/D VGND VGND VPWR VPWR _32210_/Q sky130_fd_sc_hd__dfxtp_1
X_17144_ _35564_/Q _35500_/Q _35436_/Q _35372_/Q _16897_/X _16898_/X VGND VGND VPWR
+ VPWR _17144_/X sky130_fd_sc_hd__mux4_1
X_33190_ _35943_/CLK _33190_/D VGND VGND VPWR VPWR _33190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32141_ _35811_/CLK _32141_/D VGND VGND VPWR VPWR _32141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17075_ _17932_/A VGND VGND VPWR VPWR _17075_/X sky130_fd_sc_hd__buf_4
XFILLER_170_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16026_ _17908_/A VGND VGND VPWR VPWR _16026_/X sky130_fd_sc_hd__clkbuf_4
X_32072_ _36171_/CLK _32072_/D VGND VGND VPWR VPWR _32072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31023_ _35734_/Q _29076_/X _31025_/S VGND VGND VPWR VPWR _31024_/A sky130_fd_sc_hd__mux2_1
X_35900_ _36028_/CLK _35900_/D VGND VGND VPWR VPWR _35900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35831_ _35831_/CLK _35831_/D VGND VGND VPWR VPWR _35831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17977_ _17973_/X _17976_/X _17834_/X VGND VGND VPWR VPWR _18003_/A sky130_fd_sc_hd__o21ba_1
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19716_ _20208_/A VGND VGND VPWR VPWR _19716_/X sky130_fd_sc_hd__clkbuf_4
X_16928_ _35814_/Q _32190_/Q _35686_/Q _35622_/Q _16607_/X _16608_/X VGND VGND VPWR
+ VPWR _16928_/X sky130_fd_sc_hd__mux4_1
X_35762_ _35827_/CLK _35762_/D VGND VGND VPWR VPWR _35762_/Q sky130_fd_sc_hd__dfxtp_1
X_32974_ _36049_/CLK _32974_/D VGND VGND VPWR VPWR _32974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34713_ _36200_/CLK _34713_/D VGND VGND VPWR VPWR _34713_/Q sky130_fd_sc_hd__dfxtp_1
X_31925_ _31925_/A VGND VGND VPWR VPWR _36161_/D sky130_fd_sc_hd__clkbuf_1
X_19647_ _20155_/A VGND VGND VPWR VPWR _19647_/X sky130_fd_sc_hd__buf_4
XFILLER_226_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35693_ _35949_/CLK _35693_/D VGND VGND VPWR VPWR _35693_/Q sky130_fd_sc_hd__dfxtp_1
X_16859_ _32996_/Q _32932_/Q _32868_/Q _32804_/Q _16636_/X _16637_/X VGND VGND VPWR
+ VPWR _16859_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_1471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34644_ _34775_/CLK _34644_/D VGND VGND VPWR VPWR _34644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19578_ _33008_/Q _32944_/Q _32880_/Q _32816_/Q _19289_/X _19290_/X VGND VGND VPWR
+ VPWR _19578_/X sky130_fd_sc_hd__mux4_1
X_31856_ _23145_/X _36129_/Q _31856_/S VGND VGND VPWR VPWR _31857_/A sky130_fd_sc_hd__mux2_1
X_18529_ _20294_/A VGND VGND VPWR VPWR _18529_/X sky130_fd_sc_hd__buf_6
X_30807_ _30807_/A VGND VGND VPWR VPWR _35631_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34575_ _35215_/CLK _34575_/D VGND VGND VPWR VPWR _34575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31787_ _36096_/Q input46/X _31805_/S VGND VGND VPWR VPWR _31788_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21540_ _34534_/Q _32422_/Q _34406_/Q _34342_/Q _21472_/X _21473_/X VGND VGND VPWR
+ VPWR _21540_/X sky130_fd_sc_hd__mux4_1
X_33526_ _34039_/CLK _33526_/D VGND VGND VPWR VPWR _33526_/Q sky130_fd_sc_hd__dfxtp_1
X_30738_ _30738_/A VGND VGND VPWR VPWR _35598_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33457_ _34033_/CLK _33457_/D VGND VGND VPWR VPWR _33457_/Q sky130_fd_sc_hd__dfxtp_1
X_21471_ _21396_/X _21469_/X _21470_/X _21399_/X VGND VGND VPWR VPWR _21471_/X sky130_fd_sc_hd__a22o_1
X_30669_ _35566_/Q _29151_/X _30683_/S VGND VGND VPWR VPWR _30670_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1042 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23210_ _23210_/A VGND VGND VPWR VPWR _32186_/D sky130_fd_sc_hd__clkbuf_1
X_20422_ _20418_/X _20421_/X _20167_/X VGND VGND VPWR VPWR _20423_/D sky130_fd_sc_hd__o21ba_1
X_32408_ _35226_/CLK _32408_/D VGND VGND VPWR VPWR _32408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36176_ _36185_/CLK _36176_/D VGND VGND VPWR VPWR _36176_/Q sky130_fd_sc_hd__dfxtp_1
X_24190_ _22997_/X _32628_/Q _24192_/S VGND VGND VPWR VPWR _24191_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33388_ _34292_/CLK _33388_/D VGND VGND VPWR VPWR _33388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35127_ _35766_/CLK _35127_/D VGND VGND VPWR VPWR _35127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23141_ _23141_/A VGND VGND VPWR VPWR _32159_/D sky130_fd_sc_hd__clkbuf_1
X_20353_ _33222_/Q _32582_/Q _35974_/Q _35910_/Q _20080_/X _20081_/X VGND VGND VPWR
+ VPWR _20353_/X sky130_fd_sc_hd__mux4_1
X_32339_ _32978_/CLK _32339_/D VGND VGND VPWR VPWR _32339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23072_ _23071_/X _32076_/Q _23075_/S VGND VGND VPWR VPWR _23073_/A sky130_fd_sc_hd__mux2_1
X_20284_ _33028_/Q _32964_/Q _32900_/Q _32836_/Q _19995_/X _19996_/X VGND VGND VPWR
+ VPWR _20284_/X sky130_fd_sc_hd__mux4_1
X_35058_ _35826_/CLK _35058_/D VGND VGND VPWR VPWR _35058_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_11_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_11_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XTAP_6218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34009_ _35284_/CLK _34009_/D VGND VGND VPWR VPWR _34009_/Q sky130_fd_sc_hd__dfxtp_1
X_26900_ input18/X VGND VGND VPWR VPWR _26900_/X sky130_fd_sc_hd__clkbuf_4
X_22023_ _35828_/Q _32206_/Q _35700_/Q _35636_/Q _21913_/X _21914_/X VGND VGND VPWR
+ VPWR _22023_/X sky130_fd_sc_hd__mux4_1
XTAP_6229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27880_ _27880_/A VGND VGND VPWR VPWR _34275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26831_ _26831_/A VGND VGND VPWR VPWR _33808_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29550_ _35036_/Q _29095_/X _29560_/S VGND VGND VPWR VPWR _29551_/A sky130_fd_sc_hd__mux2_1
X_26762_ _26762_/A VGND VGND VPWR VPWR _33777_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_26_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_26_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XTAP_4849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23974_ _24106_/S VGND VGND VPWR VPWR _23993_/S sky130_fd_sc_hd__buf_4
XFILLER_25_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28501_ _28501_/A VGND VGND VPWR VPWR _34570_/D sky130_fd_sc_hd__clkbuf_1
X_25713_ _33282_/Q _24407_/X _25727_/S VGND VGND VPWR VPWR _25714_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22925_ _22925_/A VGND VGND VPWR VPWR _32028_/D sky130_fd_sc_hd__clkbuf_1
X_26693_ _26693_/A VGND VGND VPWR VPWR _33744_/D sky130_fd_sc_hd__clkbuf_1
X_29481_ _29481_/A VGND VGND VPWR VPWR _35003_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28432_ _28432_/A VGND VGND VPWR VPWR _34537_/D sky130_fd_sc_hd__clkbuf_1
X_25644_ _25644_/A VGND VGND VPWR VPWR _33249_/D sky130_fd_sc_hd__clkbuf_1
X_22856_ _33037_/Q _32973_/Q _32909_/Q _32845_/Q _20580_/X _20583_/X VGND VGND VPWR
+ VPWR _22856_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28363_ _34505_/Q _24428_/X _28363_/S VGND VGND VPWR VPWR _28364_/A sky130_fd_sc_hd__mux2_1
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21807_ _21801_/X _21806_/X _21728_/X VGND VGND VPWR VPWR _21831_/A sky130_fd_sc_hd__o21ba_1
X_25575_ _33218_/Q _24407_/X _25589_/S VGND VGND VPWR VPWR _25576_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22787_ _22501_/X _22785_/X _22786_/X _22506_/X VGND VGND VPWR VPWR _22787_/X sky130_fd_sc_hd__a22o_1
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27314_ _34008_/Q _24276_/X _27332_/S VGND VGND VPWR VPWR _27315_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24526_ _24526_/A VGND VGND VPWR VPWR _32756_/D sky130_fd_sc_hd__clkbuf_1
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28294_ _34472_/Q _24326_/X _28300_/S VGND VGND VPWR VPWR _28295_/A sky130_fd_sc_hd__mux2_1
X_21738_ _21732_/X _21735_/X _21736_/X _21737_/X VGND VGND VPWR VPWR _21763_/B sky130_fd_sc_hd__o211a_1
XFILLER_196_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27245_ _27245_/A VGND VGND VPWR VPWR _33975_/D sky130_fd_sc_hd__clkbuf_1
X_24457_ _24457_/A VGND VGND VPWR VPWR _32723_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21669_ _21662_/X _21668_/X _21383_/X _21384_/X VGND VGND VPWR VPWR _21686_/B sky130_fd_sc_hd__o211a_1
XFILLER_240_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23408_ _23408_/A VGND VGND VPWR VPWR _32262_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27176_ _26850_/X _33943_/Q _27176_/S VGND VGND VPWR VPWR _27177_/A sky130_fd_sc_hd__mux2_1
X_24388_ input41/X VGND VGND VPWR VPWR _24388_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26127_ _26127_/A VGND VGND VPWR VPWR _33477_/D sky130_fd_sc_hd__clkbuf_1
X_23339_ input58/X VGND VGND VPWR VPWR _23339_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_180_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26058_ _26058_/A VGND VGND VPWR VPWR _33444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17900_ _17900_/A VGND VGND VPWR VPWR _32001_/D sky130_fd_sc_hd__clkbuf_2
X_25009_ _25009_/A VGND VGND VPWR VPWR _32979_/D sky130_fd_sc_hd__clkbuf_1
X_18880_ _18593_/X _18878_/X _18879_/X _18596_/X VGND VGND VPWR VPWR _18880_/X sky130_fd_sc_hd__a22o_1
XFILLER_79_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17831_ _33536_/Q _33472_/Q _33408_/Q _33344_/Q _17829_/X _17830_/X VGND VGND VPWR
+ VPWR _17831_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29817_ _29817_/A VGND VGND VPWR VPWR _35162_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17762_ _17762_/A VGND VGND VPWR VPWR _17762_/X sky130_fd_sc_hd__clkbuf_4
X_29748_ _35130_/Q _29188_/X _29758_/S VGND VGND VPWR VPWR _29749_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19501_ _19495_/X _19498_/X _19499_/X _19500_/X VGND VGND VPWR VPWR _19501_/X sky130_fd_sc_hd__a22o_1
X_16713_ _32992_/Q _32928_/Q _32864_/Q _32800_/Q _16636_/X _16637_/X VGND VGND VPWR
+ VPWR _16713_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17693_ _17408_/X _17691_/X _17692_/X _17414_/X VGND VGND VPWR VPWR _17693_/X sky130_fd_sc_hd__a22o_1
X_29679_ _35097_/Q _29086_/X _29695_/S VGND VGND VPWR VPWR _29680_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_290_CLK clkbuf_6_57__f_CLK/X VGND VGND VPWR VPWR _32959_/CLK sky130_fd_sc_hd__clkbuf_16
X_31710_ _31710_/A VGND VGND VPWR VPWR _36059_/D sky130_fd_sc_hd__clkbuf_1
X_19432_ _19355_/X _19430_/X _19431_/X _19361_/X VGND VGND VPWR VPWR _19432_/X sky130_fd_sc_hd__a22o_1
X_16644_ _17858_/A VGND VGND VPWR VPWR _16644_/X sky130_fd_sc_hd__buf_4
XFILLER_207_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32690_ _34032_/CLK _32690_/D VGND VGND VPWR VPWR _32690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31641_ _36027_/Q input40/X _31649_/S VGND VGND VPWR VPWR _31642_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19363_ _20208_/A VGND VGND VPWR VPWR _19363_/X sky130_fd_sc_hd__buf_4
XFILLER_245_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16575_ _35804_/Q _32179_/Q _35676_/Q _35612_/Q _16254_/X _16255_/X VGND VGND VPWR
+ VPWR _16575_/X sky130_fd_sc_hd__mux4_1
XFILLER_188_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18314_ _20201_/A VGND VGND VPWR VPWR _18314_/X sky130_fd_sc_hd__buf_2
XFILLER_31_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34360_ _35577_/CLK _34360_/D VGND VGND VPWR VPWR _34360_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19294_ _20155_/A VGND VGND VPWR VPWR _19294_/X sky130_fd_sc_hd__buf_4
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31572_ _35994_/Q input4/X _31586_/S VGND VGND VPWR VPWR _31573_/A sky130_fd_sc_hd__mux2_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33311_ _33692_/CLK _33311_/D VGND VGND VPWR VPWR _33311_/Q sky130_fd_sc_hd__dfxtp_1
X_18245_ _33805_/Q _33741_/Q _33677_/Q _33613_/Q _16020_/X _16021_/X VGND VGND VPWR
+ VPWR _18245_/X sky130_fd_sc_hd__mux4_1
X_30523_ _23228_/X _35497_/Q _30527_/S VGND VGND VPWR VPWR _30524_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34291_ _34291_/CLK _34291_/D VGND VGND VPWR VPWR _34291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36030_ _36031_/CLK _36030_/D VGND VGND VPWR VPWR _36030_/Q sky130_fd_sc_hd__dfxtp_1
X_30454_ _30454_/A VGND VGND VPWR VPWR _35464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33242_ _33244_/CLK _33242_/D VGND VGND VPWR VPWR _33242_/Q sky130_fd_sc_hd__dfxtp_1
X_18176_ _34826_/Q _34762_/Q _34698_/Q _34634_/Q _17994_/X _17995_/X VGND VGND VPWR
+ VPWR _18176_/X sky130_fd_sc_hd__mux4_1
XFILLER_198_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17127_ _16849_/X _17125_/X _17126_/X _16852_/X VGND VGND VPWR VPWR _17127_/X sky130_fd_sc_hd__a22o_1
X_33173_ _36114_/CLK _33173_/D VGND VGND VPWR VPWR _33173_/Q sky130_fd_sc_hd__dfxtp_1
X_30385_ _30385_/A VGND VGND VPWR VPWR _35431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32124_ _35562_/CLK _32124_/D VGND VGND VPWR VPWR _32124_/Q sky130_fd_sc_hd__dfxtp_1
X_17058_ _17982_/A VGND VGND VPWR VPWR _17058_/X sky130_fd_sc_hd__buf_6
XFILLER_171_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16009_ _15997_/X _16000_/X _16003_/X _16008_/X VGND VGND VPWR VPWR _16009_/X sky130_fd_sc_hd__a22o_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32055_ _36023_/CLK _32055_/D VGND VGND VPWR VPWR _32055_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31006_ _31138_/S VGND VGND VPWR VPWR _31025_/S sky130_fd_sc_hd__buf_4
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35814_ _35814_/CLK _35814_/D VGND VGND VPWR VPWR _35814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35745_ _35745_/CLK _35745_/D VGND VGND VPWR VPWR _35745_/Q sky130_fd_sc_hd__dfxtp_1
X_32957_ _36095_/CLK _32957_/D VGND VGND VPWR VPWR _32957_/Q sky130_fd_sc_hd__dfxtp_1
X_20971_ _20893_/X _20967_/X _20970_/X _20896_/X VGND VGND VPWR VPWR _20971_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_281_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _36156_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_26_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22710_ _35784_/Q _35144_/Q _34504_/Q _33864_/Q _22446_/X _22447_/X VGND VGND VPWR
+ VPWR _22710_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31908_ _31908_/A VGND VGND VPWR VPWR _36153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23690_ _32394_/Q _23336_/X _23696_/S VGND VGND VPWR VPWR _23691_/A sky130_fd_sc_hd__mux2_1
X_35676_ _35803_/CLK _35676_/D VGND VGND VPWR VPWR _35676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32888_ _36024_/CLK _32888_/D VGND VGND VPWR VPWR _32888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34627_ _35331_/CLK _34627_/D VGND VGND VPWR VPWR _34627_/Q sky130_fd_sc_hd__dfxtp_1
X_22641_ _22637_/X _22640_/X _22434_/X VGND VGND VPWR VPWR _22663_/A sky130_fd_sc_hd__o21ba_2
XFILLER_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31839_ _31839_/A VGND VGND VPWR VPWR _36120_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25360_ _25041_/X _33118_/Q _25366_/S VGND VGND VPWR VPWR _25361_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22572_ _34308_/Q _34244_/Q _34180_/Q _34116_/Q _22395_/X _22396_/X VGND VGND VPWR
+ VPWR _22572_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34558_ _35581_/CLK _34558_/D VGND VGND VPWR VPWR _34558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24311_ input14/X VGND VGND VPWR VPWR _24311_/X sky130_fd_sc_hd__buf_4
XFILLER_221_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33509_ _35991_/CLK _33509_/D VGND VGND VPWR VPWR _33509_/Q sky130_fd_sc_hd__dfxtp_1
X_21523_ _22582_/A VGND VGND VPWR VPWR _21523_/X sky130_fd_sc_hd__buf_8
XFILLER_193_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25291_ _25140_/X _33086_/Q _25293_/S VGND VGND VPWR VPWR _25292_/A sky130_fd_sc_hd__mux2_1
X_34489_ _35766_/CLK _34489_/D VGND VGND VPWR VPWR _34489_/Q sky130_fd_sc_hd__dfxtp_1
X_27030_ _27030_/A VGND VGND VPWR VPWR _33873_/D sky130_fd_sc_hd__clkbuf_1
X_36228_ _36228_/CLK _36228_/D VGND VGND VPWR VPWR _36228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24242_ _23074_/X _32653_/Q _24242_/S VGND VGND VPWR VPWR _24243_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21454_ _21448_/X _21453_/X _21375_/X VGND VGND VPWR VPWR _21478_/A sky130_fd_sc_hd__o21ba_1
XFILLER_222_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20405_ _32520_/Q _32392_/Q _32072_/Q _36040_/Q _20282_/X _19307_/A VGND VGND VPWR
+ VPWR _20405_/X sky130_fd_sc_hd__mux4_1
XFILLER_193_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36159_ _36159_/CLK _36159_/D VGND VGND VPWR VPWR _36159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24173_ _24242_/S VGND VGND VPWR VPWR _24192_/S sky130_fd_sc_hd__buf_4
X_21385_ _21379_/X _21382_/X _21383_/X _21384_/X VGND VGND VPWR VPWR _21410_/B sky130_fd_sc_hd__o211a_1
XFILLER_208_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23124_ input4/X VGND VGND VPWR VPWR _23124_/X sky130_fd_sc_hd__buf_6
X_20336_ _34310_/Q _34246_/Q _34182_/Q _34118_/Q _20095_/X _20096_/X VGND VGND VPWR
+ VPWR _20336_/X sky130_fd_sc_hd__mux4_1
X_28981_ _28981_/A VGND VGND VPWR VPWR _34797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23055_ _23055_/A VGND VGND VPWR VPWR _32070_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27932_ _27932_/A VGND VGND VPWR VPWR _34300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20267_ _20160_/X _20265_/X _20266_/X _20165_/X VGND VGND VPWR VPWR _20267_/X sky130_fd_sc_hd__a22o_1
XTAP_6026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22006_ _21802_/X _22004_/X _22005_/X _21805_/X VGND VGND VPWR VPWR _22006_/X sky130_fd_sc_hd__a22o_1
XFILLER_248_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20198_ _20194_/X _20197_/X _20167_/X VGND VGND VPWR VPWR _20199_/D sky130_fd_sc_hd__o21ba_1
XTAP_5325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27863_ _27863_/A VGND VGND VPWR VPWR _34267_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29602_ _35061_/Q _29172_/X _29602_/S VGND VGND VPWR VPWR _29603_/A sky130_fd_sc_hd__mux2_1
X_26814_ _26814_/A VGND VGND VPWR VPWR _33802_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27794_ _34235_/Q _24385_/X _27802_/S VGND VGND VPWR VPWR _27795_/A sky130_fd_sc_hd__mux2_1
XTAP_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29533_ _35028_/Q _29070_/X _29539_/S VGND VGND VPWR VPWR _29534_/A sky130_fd_sc_hd__mux2_1
XTAP_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23957_ _23957_/A VGND VGND VPWR VPWR _32518_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26745_ _26745_/A VGND VGND VPWR VPWR _33769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_272_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _34302_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_901 _26142_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_912 _26829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22908_ _22907_/X _32023_/Q _22908_/S VGND VGND VPWR VPWR _22909_/A sky130_fd_sc_hd__mux2_1
XTAP_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26676_ _26676_/A VGND VGND VPWR VPWR _33737_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29464_ _29464_/A VGND VGND VPWR VPWR _34995_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_923 _27154_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23888_ _23888_/A VGND VGND VPWR VPWR _32485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_934 _29247_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_945 _29517_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_956 _29787_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28415_ _28415_/A VGND VGND VPWR VPWR _34529_/D sky130_fd_sc_hd__clkbuf_1
X_22839_ _34572_/Q _32460_/Q _34444_/Q _34380_/Q _20663_/X _20665_/X VGND VGND VPWR
+ VPWR _22839_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25627_ _33241_/Q _24280_/X _25643_/S VGND VGND VPWR VPWR _25628_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29395_ _29395_/A VGND VGND VPWR VPWR _34962_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_967 _31138_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_978 _17855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_989 _17860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16360_ _32982_/Q _32918_/Q _32854_/Q _32790_/Q _16283_/X _16284_/X VGND VGND VPWR
+ VPWR _16360_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28346_ _28346_/A VGND VGND VPWR VPWR _34496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25558_ _33210_/Q _24382_/X _25568_/S VGND VGND VPWR VPWR _25559_/A sky130_fd_sc_hd__mux2_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24509_ _22972_/X _32748_/Q _24527_/S VGND VGND VPWR VPWR _24510_/A sky130_fd_sc_hd__mux2_1
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28277_ _34464_/Q _24301_/X _28279_/S VGND VGND VPWR VPWR _28278_/A sky130_fd_sc_hd__mux2_1
X_16291_ _17858_/A VGND VGND VPWR VPWR _16291_/X sky130_fd_sc_hd__buf_4
X_25489_ _33177_/Q _24280_/X _25505_/S VGND VGND VPWR VPWR _25490_/A sky130_fd_sc_hd__mux2_1
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18030_ _35077_/Q _35013_/Q _34949_/Q _34885_/Q _17862_/X _17863_/X VGND VGND VPWR
+ VPWR _18030_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27228_ _27228_/A VGND VGND VPWR VPWR _33967_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27159_ _27159_/A VGND VGND VPWR VPWR _33934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30170_ _35330_/Q _29213_/X _30184_/S VGND VGND VPWR VPWR _30171_/A sky130_fd_sc_hd__mux2_1
X_19981_ _19977_/X _19980_/X _19814_/X VGND VGND VPWR VPWR _19982_/D sky130_fd_sc_hd__o21ba_1
XFILLER_207_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18932_ _32734_/Q _32670_/Q _32606_/Q _36062_/Q _18866_/X _18650_/X VGND VGND VPWR
+ VPWR _18932_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1300 _17867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1311 input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1322 _31993_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1333 _20232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18863_ _34012_/Q _33948_/Q _33884_/Q _32156_/Q _18614_/X _18615_/X VGND VGND VPWR
+ VPWR _18863_/X sky130_fd_sc_hd__mux4_1
XTAP_6560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1344 _22501_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1355 _22508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1366 _24354_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17814_ _33215_/Q _32575_/Q _35967_/Q _35903_/Q _17780_/X _17781_/X VGND VGND VPWR
+ VPWR _17814_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1377 _26869_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33860_ _35780_/CLK _33860_/D VGND VGND VPWR VPWR _33860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1388 _31408_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18794_ _20158_/A VGND VGND VPWR VPWR _18794_/X sky130_fd_sc_hd__buf_4
XTAP_5870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32811_ _36075_/CLK _32811_/D VGND VGND VPWR VPWR _32811_/Q sky130_fd_sc_hd__dfxtp_1
X_17745_ _34813_/Q _34749_/Q _34685_/Q _34621_/Q _17641_/X _17642_/X VGND VGND VPWR
+ VPWR _17745_/X sky130_fd_sc_hd__mux4_1
X_33791_ _34303_/CLK _33791_/D VGND VGND VPWR VPWR _33791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_263_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _36159_/CLK sky130_fd_sc_hd__clkbuf_16
X_35530_ _35978_/CLK _35530_/D VGND VGND VPWR VPWR _35530_/Q sky130_fd_sc_hd__dfxtp_1
X_32742_ _36135_/CLK _32742_/D VGND VGND VPWR VPWR _32742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17676_ _35323_/Q _35259_/Q _35195_/Q _32315_/Q _17359_/X _17360_/X VGND VGND VPWR
+ VPWR _17676_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19415_ _35051_/Q _34987_/Q _34923_/Q _34859_/Q _19103_/X _19104_/X VGND VGND VPWR
+ VPWR _19415_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35461_ _35909_/CLK _35461_/D VGND VGND VPWR VPWR _35461_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16627_ _16489_/X _16625_/X _16626_/X _16494_/X VGND VGND VPWR VPWR _16627_/X sky130_fd_sc_hd__a22o_1
X_32673_ _36065_/CLK _32673_/D VGND VGND VPWR VPWR _32673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34412_ _35304_/CLK _34412_/D VGND VGND VPWR VPWR _34412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19346_ _19346_/A _19346_/B _19346_/C _19346_/D VGND VGND VPWR VPWR _19347_/A sky130_fd_sc_hd__or4_4
X_31624_ _36019_/Q input31/X _31628_/S VGND VGND VPWR VPWR _31625_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35392_ _35909_/CLK _35392_/D VGND VGND VPWR VPWR _35392_/Q sky130_fd_sc_hd__dfxtp_1
X_16558_ _16558_/A VGND VGND VPWR VPWR _31963_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34343_ _35302_/CLK _34343_/D VGND VGND VPWR VPWR _34343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_1167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31555_ _35986_/Q input45/X _31565_/S VGND VGND VPWR VPWR _31556_/A sky130_fd_sc_hd__mux2_1
X_19277_ _19277_/A VGND VGND VPWR VPWR _32103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16489_ _17901_/A VGND VGND VPWR VPWR _16489_/X sky130_fd_sc_hd__buf_4
XFILLER_164_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18228_ _18224_/X _18227_/X _17842_/A _17843_/A VGND VGND VPWR VPWR _18243_/B sky130_fd_sc_hd__o211a_1
X_30506_ _23145_/X _35489_/Q _30506_/S VGND VGND VPWR VPWR _30507_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34274_ _35992_/CLK _34274_/D VGND VGND VPWR VPWR _34274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31486_ _31486_/A VGND VGND VPWR VPWR _35953_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36013_ _36013_/CLK _36013_/D VGND VGND VPWR VPWR _36013_/Q sky130_fd_sc_hd__dfxtp_1
X_33225_ _35975_/CLK _33225_/D VGND VGND VPWR VPWR _33225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18159_ _34058_/Q _33994_/Q _33930_/Q _32266_/Q _16058_/X _16060_/X VGND VGND VPWR
+ VPWR _18159_/X sky130_fd_sc_hd__mux4_1
X_30437_ _23303_/X _35456_/Q _30455_/S VGND VGND VPWR VPWR _30438_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33156_ _36166_/CLK _33156_/D VGND VGND VPWR VPWR _33156_/Q sky130_fd_sc_hd__dfxtp_1
X_21170_ _22582_/A VGND VGND VPWR VPWR _21170_/X sky130_fd_sc_hd__buf_6
XFILLER_117_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30368_ _30368_/A VGND VGND VPWR VPWR _35423_/D sky130_fd_sc_hd__clkbuf_1
X_20121_ _35071_/Q _35007_/Q _34943_/Q _34879_/Q _19809_/X _19810_/X VGND VGND VPWR
+ VPWR _20121_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32107_ _35552_/CLK _32107_/D VGND VGND VPWR VPWR _32107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30299_ _30299_/A VGND VGND VPWR VPWR _35391_/D sky130_fd_sc_hd__clkbuf_1
X_33087_ _36097_/CLK _33087_/D VGND VGND VPWR VPWR _33087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20052_ _20052_/A _20052_/B _20052_/C _20052_/D VGND VGND VPWR VPWR _20053_/A sky130_fd_sc_hd__or4_4
XFILLER_63_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32038_ _36005_/CLK _32038_/D VGND VGND VPWR VPWR _32038_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24860_ _22886_/X _32912_/Q _24874_/S VGND VGND VPWR VPWR _24861_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23811_ _23811_/A VGND VGND VPWR VPWR _32449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24791_ _24791_/A VGND VGND VPWR VPWR _32879_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33989_ _34057_/CLK _33989_/D VGND VGND VPWR VPWR _33989_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_254_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _36165_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26530_ _26530_/A VGND VGND VPWR VPWR _33668_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_208 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35728_ _35728_/CLK _35728_/D VGND VGND VPWR VPWR _35728_/Q sky130_fd_sc_hd__dfxtp_1
X_23742_ _22938_/X _32417_/Q _23742_/S VGND VGND VPWR VPWR _23743_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20954_ _33238_/Q _36118_/Q _33110_/Q _33046_/Q _20952_/X _20953_/X VGND VGND VPWR
+ VPWR _20954_/X sky130_fd_sc_hd__mux4_1
XANTENNA_219 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26461_ _26461_/A VGND VGND VPWR VPWR _33635_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35659_ _35787_/CLK _35659_/D VGND VGND VPWR VPWR _35659_/Q sky130_fd_sc_hd__dfxtp_1
X_23673_ _23673_/A VGND VGND VPWR VPWR _32385_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20885_ _32980_/Q _32916_/Q _32852_/Q _32788_/Q _20883_/X _20884_/X VGND VGND VPWR
+ VPWR _20885_/X sky130_fd_sc_hd__mux4_1
X_28200_ _28200_/A VGND VGND VPWR VPWR _34427_/D sky130_fd_sc_hd__clkbuf_1
X_25412_ _25412_/A VGND VGND VPWR VPWR _33142_/D sky130_fd_sc_hd__clkbuf_1
X_22624_ _22305_/X _22622_/X _22623_/X _22308_/X VGND VGND VPWR VPWR _22624_/X sky130_fd_sc_hd__a22o_1
X_29180_ _34871_/Q _29179_/X _29204_/S VGND VGND VPWR VPWR _29181_/A sky130_fd_sc_hd__mux2_1
X_26392_ _25156_/X _33603_/Q _26404_/S VGND VGND VPWR VPWR _26393_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28131_ _28131_/A VGND VGND VPWR VPWR _34394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25343_ _25016_/X _33110_/Q _25345_/S VGND VGND VPWR VPWR _25344_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22555_ _22300_/X _22553_/X _22554_/X _22303_/X VGND VGND VPWR VPWR _22555_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28062_ _26959_/X _34362_/Q _28072_/S VGND VGND VPWR VPWR _28063_/A sky130_fd_sc_hd__mux2_1
X_21506_ _34533_/Q _32421_/Q _34405_/Q _34341_/Q _21472_/X _21473_/X VGND VGND VPWR
+ VPWR _21506_/X sky130_fd_sc_hd__mux4_1
X_25274_ _25322_/S VGND VGND VPWR VPWR _25293_/S sky130_fd_sc_hd__buf_4
X_22486_ _35777_/Q _35137_/Q _34497_/Q _33857_/Q _22446_/X _22447_/X VGND VGND VPWR
+ VPWR _22486_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27013_ _27013_/A VGND VGND VPWR VPWR _33867_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24225_ _24225_/A VGND VGND VPWR VPWR _32644_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21437_ _35043_/Q _34979_/Q _34915_/Q _34851_/Q _21403_/X _21404_/X VGND VGND VPWR
+ VPWR _21437_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24156_ _24156_/A VGND VGND VPWR VPWR _32611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21368_ _34274_/Q _34210_/Q _34146_/Q _34082_/Q _21336_/X _21337_/X VGND VGND VPWR
+ VPWR _21368_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23107_ _23107_/A VGND VGND VPWR VPWR _32148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20319_ _35845_/Q _32224_/Q _35717_/Q _35653_/Q _18289_/X _18291_/X VGND VGND VPWR
+ VPWR _20319_/X sky130_fd_sc_hd__mux4_1
X_24087_ _24087_/A VGND VGND VPWR VPWR _32579_/D sky130_fd_sc_hd__clkbuf_1
X_28964_ _28964_/A VGND VGND VPWR VPWR _34789_/D sky130_fd_sc_hd__clkbuf_1
X_21299_ _34016_/Q _33952_/Q _33888_/Q _32160_/Q _21267_/X _21268_/X VGND VGND VPWR
+ VPWR _21299_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23038_ input47/X VGND VGND VPWR VPWR _23038_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27915_ _27915_/A VGND VGND VPWR VPWR _34292_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28895_ _26993_/X _34757_/Q _28903_/S VGND VGND VPWR VPWR _28896_/A sky130_fd_sc_hd__mux2_1
XTAP_5122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_493_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _35039_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27846_ _27846_/A VGND VGND VPWR VPWR _34259_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27777_ _34227_/Q _24360_/X _27781_/S VGND VGND VPWR VPWR _27778_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24989_ input1/X VGND VGND VPWR VPWR _24989_/X sky130_fd_sc_hd__buf_4
XTAP_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_245_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _34309_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29516_ _29516_/A VGND VGND VPWR VPWR _35020_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _17416_/X _17528_/X _17529_/X _17420_/X VGND VGND VPWR VPWR _17530_/X sky130_fd_sc_hd__a22o_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26728_ _26728_/A VGND VGND VPWR VPWR _33761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_720 _21754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_731 _20980_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_742 _21763_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29447_ _29447_/A VGND VGND VPWR VPWR _34987_/D sky130_fd_sc_hd__clkbuf_1
X_17461_ _33205_/Q _32565_/Q _35957_/Q _35893_/Q _17427_/X _17428_/X VGND VGND VPWR
+ VPWR _17461_/X sky130_fd_sc_hd__mux4_1
X_26659_ _25150_/X _33729_/Q _26675_/S VGND VGND VPWR VPWR _26660_/A sky130_fd_sc_hd__mux2_1
XANTENNA_753 _22443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_764 _22500_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_775 _22578_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19200_ _33189_/Q _32549_/Q _35941_/Q _35877_/Q _19021_/X _19022_/X VGND VGND VPWR
+ VPWR _19200_/X sky130_fd_sc_hd__mux4_1
XANTENNA_786 _22634_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16412_ _16412_/A _16412_/B _16412_/C _16412_/D VGND VGND VPWR VPWR _16413_/A sky130_fd_sc_hd__or4_4
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_797 _22874_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29378_ _23339_/X _34955_/Q _29382_/S VGND VGND VPWR VPWR _29379_/A sky130_fd_sc_hd__mux2_1
X_17392_ _34803_/Q _34739_/Q _34675_/Q _34611_/Q _17288_/X _17289_/X VGND VGND VPWR
+ VPWR _17392_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19131_ _18946_/X _19129_/X _19130_/X _18949_/X VGND VGND VPWR VPWR _19131_/X sky130_fd_sc_hd__a22o_1
X_16343_ _34262_/Q _34198_/Q _34134_/Q _34070_/Q _16005_/X _16007_/X VGND VGND VPWR
+ VPWR _16343_/X sky130_fd_sc_hd__mux4_1
XFILLER_207_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28329_ _28329_/A VGND VGND VPWR VPWR _34488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16274_ _16136_/X _16272_/X _16273_/X _16141_/X VGND VGND VPWR VPWR _16274_/X sky130_fd_sc_hd__a22o_1
XFILLER_121_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19062_ _35041_/Q _34977_/Q _34913_/Q _34849_/Q _18750_/X _18751_/X VGND VGND VPWR
+ VPWR _19062_/X sky130_fd_sc_hd__mux4_1
X_31340_ _35884_/Q input24/X _31358_/S VGND VGND VPWR VPWR _31341_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18013_ _33285_/Q _36165_/Q _33157_/Q _33093_/Q _17764_/X _17765_/X VGND VGND VPWR
+ VPWR _18013_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31271_ _35852_/Q input59/X _31273_/S VGND VGND VPWR VPWR _31272_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33010_ _35765_/CLK _33010_/D VGND VGND VPWR VPWR _33010_/Q sky130_fd_sc_hd__dfxtp_1
X_30222_ _30222_/A VGND VGND VPWR VPWR _35354_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_1417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1070 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30153_ _35322_/Q _29188_/X _30163_/S VGND VGND VPWR VPWR _30154_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19964_ _19716_/X _19962_/X _19963_/X _19720_/X VGND VGND VPWR VPWR _19964_/X sky130_fd_sc_hd__a22o_1
X_18915_ _18911_/X _18914_/X _18741_/X VGND VGND VPWR VPWR _18923_/C sky130_fd_sc_hd__o21ba_1
XFILLER_68_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34961_ _36204_/CLK _34961_/D VGND VGND VPWR VPWR _34961_/Q sky130_fd_sc_hd__dfxtp_1
X_30084_ _35289_/Q _29086_/X _30100_/S VGND VGND VPWR VPWR _30085_/A sky130_fd_sc_hd__mux2_1
XTAP_7091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1130 _17842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19895_ _19708_/X _19893_/X _19894_/X _19714_/X VGND VGND VPWR VPWR _19895_/X sky130_fd_sc_hd__a22o_1
XFILLER_110_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1141 _20201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_484_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _35743_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33912_ _36152_/CLK _33912_/D VGND VGND VPWR VPWR _33912_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1152 _22455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18846_ _35547_/Q _35483_/Q _35419_/Q _35355_/Q _18844_/X _18845_/X VGND VGND VPWR
+ VPWR _18846_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1163 _22462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_34892_ _35277_/CLK _34892_/D VGND VGND VPWR VPWR _34892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1174 _21607_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1185 _22217_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1196 _22935_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33843_ _35827_/CLK _33843_/D VGND VGND VPWR VPWR _33843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18777_ _33177_/Q _32537_/Q _35929_/Q _35865_/Q _18668_/X _18669_/X VGND VGND VPWR
+ VPWR _18777_/X sky130_fd_sc_hd__mux4_1
XFILLER_243_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15989_ _17795_/A VGND VGND VPWR VPWR _15989_/X sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_236_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _35328_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_236_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17728_ _34045_/Q _33981_/Q _33917_/Q _32253_/Q _17726_/X _17727_/X VGND VGND VPWR
+ VPWR _17728_/X sky130_fd_sc_hd__mux4_1
X_33774_ _34288_/CLK _33774_/D VGND VGND VPWR VPWR _33774_/Q sky130_fd_sc_hd__dfxtp_1
X_30986_ _30986_/A VGND VGND VPWR VPWR _35716_/D sky130_fd_sc_hd__clkbuf_1
X_35513_ _35578_/CLK _35513_/D VGND VGND VPWR VPWR _35513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32725_ _36116_/CLK _32725_/D VGND VGND VPWR VPWR _32725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17659_ _32763_/Q _32699_/Q _32635_/Q _36091_/Q _17625_/X _17409_/X VGND VGND VPWR
+ VPWR _17659_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35444_ _35956_/CLK _35444_/D VGND VGND VPWR VPWR _35444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20670_ input75/X input76/X VGND VGND VPWR VPWR _22453_/A sky130_fd_sc_hd__or2_4
X_32656_ _33234_/CLK _32656_/D VGND VGND VPWR VPWR _32656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31607_ _36011_/Q input22/X _31607_/S VGND VGND VPWR VPWR _31608_/A sky130_fd_sc_hd__mux2_1
X_19329_ _33001_/Q _32937_/Q _32873_/Q _32809_/Q _19289_/X _19290_/X VGND VGND VPWR
+ VPWR _19329_/X sky130_fd_sc_hd__mux4_1
X_35375_ _35822_/CLK _35375_/D VGND VGND VPWR VPWR _35375_/Q sky130_fd_sc_hd__dfxtp_1
X_32587_ _35979_/CLK _32587_/D VGND VGND VPWR VPWR _32587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34326_ _34706_/CLK _34326_/D VGND VGND VPWR VPWR _34326_/Q sky130_fd_sc_hd__dfxtp_1
X_22340_ _22300_/X _22338_/X _22339_/X _22303_/X VGND VGND VPWR VPWR _22340_/X sky130_fd_sc_hd__a22o_1
XFILLER_137_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31538_ _31538_/A VGND VGND VPWR VPWR _35978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34257_ _34259_/CLK _34257_/D VGND VGND VPWR VPWR _34257_/Q sky130_fd_sc_hd__dfxtp_1
X_22271_ _35579_/Q _35515_/Q _35451_/Q _35387_/Q _22203_/X _22204_/X VGND VGND VPWR
+ VPWR _22271_/X sky130_fd_sc_hd__mux4_1
X_31469_ _31469_/A VGND VGND VPWR VPWR _35945_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24010_ _22932_/X _32543_/Q _24014_/S VGND VGND VPWR VPWR _24011_/A sky130_fd_sc_hd__mux2_1
X_33208_ _36024_/CLK _33208_/D VGND VGND VPWR VPWR _33208_/Q sky130_fd_sc_hd__dfxtp_1
X_21222_ _21218_/X _21221_/X _21055_/X VGND VGND VPWR VPWR _21223_/D sky130_fd_sc_hd__o21ba_1
XFILLER_219_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34188_ _36048_/CLK _34188_/D VGND VGND VPWR VPWR _34188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21153_ _34523_/Q _32411_/Q _34395_/Q _34331_/Q _21119_/X _21120_/X VGND VGND VPWR
+ VPWR _21153_/X sky130_fd_sc_hd__mux4_1
X_33139_ _36147_/CLK _33139_/D VGND VGND VPWR VPWR _33139_/Q sky130_fd_sc_hd__dfxtp_1
X_20104_ _33279_/Q _36159_/Q _33151_/Q _33087_/Q _20064_/X _20065_/X VGND VGND VPWR
+ VPWR _20104_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25961_ _25961_/A VGND VGND VPWR VPWR _33398_/D sky130_fd_sc_hd__clkbuf_1
X_21084_ _35033_/Q _34969_/Q _34905_/Q _34841_/Q _21050_/X _21051_/X VGND VGND VPWR
+ VPWR _21084_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27700_ _34190_/Q _24244_/X _27718_/S VGND VGND VPWR VPWR _27701_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_475_CLK clkbuf_6_8__f_CLK/X VGND VGND VPWR VPWR _35876_/CLK sky130_fd_sc_hd__clkbuf_16
X_20035_ _33021_/Q _32957_/Q _32893_/Q _32829_/Q _19995_/X _19996_/X VGND VGND VPWR
+ VPWR _20035_/X sky130_fd_sc_hd__mux4_1
X_24912_ _22963_/X _32937_/Q _24916_/S VGND VGND VPWR VPWR _24913_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25892_ _25016_/X _33366_/Q _25894_/S VGND VGND VPWR VPWR _25893_/A sky130_fd_sc_hd__mux2_1
X_28680_ _26875_/X _34655_/Q _28684_/S VGND VGND VPWR VPWR _28681_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27631_ _27631_/A VGND VGND VPWR VPWR _34157_/D sky130_fd_sc_hd__clkbuf_1
X_24843_ _24843_/A VGND VGND VPWR VPWR _32904_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_838 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_227_CLK clkbuf_6_54__f_CLK/X VGND VGND VPWR VPWR _36038_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27562_ _27562_/A VGND VGND VPWR VPWR _30870_/B sky130_fd_sc_hd__buf_6
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24774_ _24774_/A VGND VGND VPWR VPWR _32871_/D sky130_fd_sc_hd__clkbuf_1
X_21986_ _35763_/Q _35123_/Q _34483_/Q _33843_/Q _21740_/X _21741_/X VGND VGND VPWR
+ VPWR _21986_/X sky130_fd_sc_hd__mux4_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_57__f_CLK clkbuf_5_28_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_57__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29301_ _23217_/X _34918_/Q _29311_/S VGND VGND VPWR VPWR _29302_/A sky130_fd_sc_hd__mux2_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26513_ _26513_/A VGND VGND VPWR VPWR _33660_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23725_ _23725_/A VGND VGND VPWR VPWR _32408_/D sky130_fd_sc_hd__clkbuf_1
X_20937_ _35029_/Q _34965_/Q _34901_/Q _34837_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _20937_/X sky130_fd_sc_hd__mux4_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27493_ _26919_/X _34093_/Q _27509_/S VGND VGND VPWR VPWR _27494_/A sky130_fd_sc_hd__mux2_1
XFILLER_226_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29232_ _34888_/Q _29231_/X _29235_/S VGND VGND VPWR VPWR _29233_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23656_ _23656_/A VGND VGND VPWR VPWR _32377_/D sky130_fd_sc_hd__clkbuf_1
X_26444_ _26444_/A VGND VGND VPWR VPWR _33627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20868_ _20687_/X _20866_/X _20867_/X _20697_/X VGND VGND VPWR VPWR _20868_/X sky130_fd_sc_hd__a22o_1
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22607_ _22501_/X _22605_/X _22606_/X _22506_/X VGND VGND VPWR VPWR _22607_/X sky130_fd_sc_hd__a22o_1
XFILLER_230_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26375_ _25131_/X _33595_/Q _26383_/S VGND VGND VPWR VPWR _26376_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29163_ input30/X VGND VGND VPWR VPWR _29163_/X sky130_fd_sc_hd__clkbuf_4
X_23587_ _23587_/A VGND VGND VPWR VPWR _32344_/D sky130_fd_sc_hd__clkbuf_1
X_20799_ _20674_/X _20797_/X _20798_/X _20684_/X VGND VGND VPWR VPWR _20799_/X sky130_fd_sc_hd__a22o_1
XFILLER_195_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28114_ _28114_/A VGND VGND VPWR VPWR _34386_/D sky130_fd_sc_hd__clkbuf_1
X_25326_ _25458_/S VGND VGND VPWR VPWR _25345_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_139_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22538_ _22538_/A VGND VGND VPWR VPWR _36226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29094_ _29094_/A VGND VGND VPWR VPWR _34843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25257_ _25257_/A VGND VGND VPWR VPWR _33069_/D sky130_fd_sc_hd__clkbuf_1
X_28045_ _26934_/X _34354_/Q _28051_/S VGND VGND VPWR VPWR _28046_/A sky130_fd_sc_hd__mux2_1
X_22469_ _22469_/A _22469_/B _22469_/C _22469_/D VGND VGND VPWR VPWR _22470_/A sky130_fd_sc_hd__or4_4
XFILLER_202_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24208_ _24208_/A VGND VGND VPWR VPWR _32636_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25188_ _25188_/A VGND VGND VPWR VPWR _33037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24139_ _24139_/A VGND VGND VPWR VPWR _32603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29996_ _29996_/A VGND VGND VPWR VPWR _35247_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16961_ _17796_/A VGND VGND VPWR VPWR _16961_/X sky130_fd_sc_hd__buf_4
X_28947_ _28947_/A VGND VGND VPWR VPWR _34781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18700_ _18588_/X _18698_/X _18699_/X _18591_/X VGND VGND VPWR VPWR _18700_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_466_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _35814_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_238_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19680_ _19355_/X _19678_/X _19679_/X _19361_/X VGND VGND VPWR VPWR _19680_/X sky130_fd_sc_hd__a22o_1
X_28878_ _26968_/X _34749_/Q _28882_/S VGND VGND VPWR VPWR _28879_/A sky130_fd_sc_hd__mux2_1
X_16892_ _16710_/X _16890_/X _16891_/X _16714_/X VGND VGND VPWR VPWR _16892_/X sky130_fd_sc_hd__a22o_1
XFILLER_204_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18631_ _18593_/X _18629_/X _18630_/X _18596_/X VGND VGND VPWR VPWR _18631_/X sky130_fd_sc_hd__a22o_1
XFILLER_237_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27829_ _34252_/Q _24437_/X _27831_/S VGND VGND VPWR VPWR _27830_/A sky130_fd_sc_hd__mux2_1
XTAP_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_218_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _35780_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_58_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30840_ _30840_/A VGND VGND VPWR VPWR _35647_/D sky130_fd_sc_hd__clkbuf_1
X_18562_ _18558_/X _18561_/X _18371_/X VGND VGND VPWR VPWR _18570_/C sky130_fd_sc_hd__o21ba_1
XTAP_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17513_ _17507_/X _17508_/X _17511_/X _17512_/X VGND VGND VPWR VPWR _17513_/X sky130_fd_sc_hd__a22o_1
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18493_ _35537_/Q _35473_/Q _35409_/Q _35345_/Q _18491_/X _18492_/X VGND VGND VPWR
+ VPWR _18493_/X sky130_fd_sc_hd__mux4_1
XTAP_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30771_ _30771_/A VGND VGND VPWR VPWR _35614_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_550 _20142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32510_ _36033_/CLK _32510_/D VGND VGND VPWR VPWR _32510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_561 _20146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_572 _20165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _34293_/Q _34229_/Q _34165_/Q _34101_/Q _17442_/X _17443_/X VGND VGND VPWR
+ VPWR _17444_/X sky130_fd_sc_hd__mux4_1
X_33490_ _33490_/CLK _33490_/D VGND VGND VPWR VPWR _33490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_583 _19449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_594 _19459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32441_ _35577_/CLK _32441_/D VGND VGND VPWR VPWR _32441_/Q sky130_fd_sc_hd__dfxtp_1
X_17375_ _34035_/Q _33971_/Q _33907_/Q _32243_/Q _17373_/X _17374_/X VGND VGND VPWR
+ VPWR _17375_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19114_ _18789_/X _19112_/X _19113_/X _18794_/X VGND VGND VPWR VPWR _19114_/X sky130_fd_sc_hd__a22o_1
XFILLER_203_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16326_ _35797_/Q _32172_/Q _35669_/Q _35605_/Q _16254_/X _16255_/X VGND VGND VPWR
+ VPWR _16326_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35160_ _35226_/CLK _35160_/D VGND VGND VPWR VPWR _35160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32372_ _34228_/CLK _32372_/D VGND VGND VPWR VPWR _32372_/Q sky130_fd_sc_hd__dfxtp_1
X_34111_ _36161_/CLK _34111_/D VGND VGND VPWR VPWR _34111_/Q sky130_fd_sc_hd__dfxtp_1
X_31323_ _35876_/Q input15/X _31337_/S VGND VGND VPWR VPWR _31324_/A sky130_fd_sc_hd__mux2_1
X_19045_ _33249_/Q _36129_/Q _33121_/Q _33057_/Q _19005_/X _19006_/X VGND VGND VPWR
+ VPWR _19045_/X sky130_fd_sc_hd__mux4_1
X_35091_ _35922_/CLK _35091_/D VGND VGND VPWR VPWR _35091_/Q sky130_fd_sc_hd__dfxtp_1
X_16257_ _35731_/Q _35091_/Q _34451_/Q _33811_/Q _16049_/X _16051_/X VGND VGND VPWR
+ VPWR _16257_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34042_ _36154_/CLK _34042_/D VGND VGND VPWR VPWR _34042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput204 _36229_/Q VGND VGND VPWR VPWR D2[55] sky130_fd_sc_hd__buf_2
X_31254_ _31254_/A VGND VGND VPWR VPWR _35843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16188_ _35793_/Q _32167_/Q _35665_/Q _35601_/Q _16045_/X _16046_/X VGND VGND VPWR
+ VPWR _16188_/X sky130_fd_sc_hd__mux4_1
Xoutput215 _36181_/Q VGND VGND VPWR VPWR D2[7] sky130_fd_sc_hd__buf_2
XFILLER_160_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput226 _32095_/Q VGND VGND VPWR VPWR D3[17] sky130_fd_sc_hd__buf_2
X_30205_ _30205_/A VGND VGND VPWR VPWR _35346_/D sky130_fd_sc_hd__clkbuf_1
Xoutput237 _32105_/Q VGND VGND VPWR VPWR D3[27] sky130_fd_sc_hd__buf_2
XFILLER_141_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput248 _32115_/Q VGND VGND VPWR VPWR D3[37] sky130_fd_sc_hd__buf_2
Xoutput259 _32125_/Q VGND VGND VPWR VPWR D3[47] sky130_fd_sc_hd__buf_2
X_31185_ _31185_/A VGND VGND VPWR VPWR _35810_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19947_ _35066_/Q _35002_/Q _34938_/Q _34874_/Q _19809_/X _19810_/X VGND VGND VPWR
+ VPWR _19947_/X sky130_fd_sc_hd__mux4_1
X_30136_ _35314_/Q _29163_/X _30142_/S VGND VGND VPWR VPWR _30137_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35993_ _35995_/CLK _35993_/D VGND VGND VPWR VPWR _35993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_457_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _34922_/CLK sky130_fd_sc_hd__clkbuf_16
X_34944_ _35075_/CLK _34944_/D VGND VGND VPWR VPWR _34944_/Q sky130_fd_sc_hd__dfxtp_1
X_30067_ _35281_/Q _29061_/X _30079_/S VGND VGND VPWR VPWR _30068_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19878_ _20231_/A VGND VGND VPWR VPWR _19878_/X sky130_fd_sc_hd__buf_6
XFILLER_110_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18829_ _18789_/X _18827_/X _18828_/X _18794_/X VGND VGND VPWR VPWR _18829_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34875_ _35386_/CLK _34875_/D VGND VGND VPWR VPWR _34875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_209_CLK clkbuf_6_52__f_CLK/X VGND VGND VPWR VPWR _35590_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21840_ _32751_/Q _32687_/Q _32623_/Q _36079_/Q _21519_/X _21656_/X VGND VGND VPWR
+ VPWR _21840_/X sky130_fd_sc_hd__mux4_1
X_33826_ _35876_/CLK _33826_/D VGND VGND VPWR VPWR _33826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33757_ _34080_/CLK _33757_/D VGND VGND VPWR VPWR _33757_/Q sky130_fd_sc_hd__dfxtp_1
X_21771_ _21767_/X _21770_/X _21728_/X VGND VGND VPWR VPWR _21793_/A sky130_fd_sc_hd__o21ba_1
X_30969_ _30969_/A VGND VGND VPWR VPWR _35708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23510_ _23510_/A VGND VGND VPWR VPWR _32309_/D sky130_fd_sc_hd__clkbuf_1
X_20722_ _20644_/X _20720_/X _20721_/X _20654_/X VGND VGND VPWR VPWR _20722_/X sky130_fd_sc_hd__a22o_1
X_32708_ _36100_/CLK _32708_/D VGND VGND VPWR VPWR _32708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24490_ _22945_/X _32739_/Q _24506_/S VGND VGND VPWR VPWR _24491_/A sky130_fd_sc_hd__mux2_1
X_33688_ _35671_/CLK _33688_/D VGND VGND VPWR VPWR _33688_/Q sky130_fd_sc_hd__dfxtp_1
X_23441_ _23441_/A VGND VGND VPWR VPWR _32276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35427_ _35940_/CLK _35427_/D VGND VGND VPWR VPWR _35427_/Q sky130_fd_sc_hd__dfxtp_1
X_20653_ _22367_/A VGND VGND VPWR VPWR _22458_/A sky130_fd_sc_hd__buf_12
X_32639_ _36097_/CLK _32639_/D VGND VGND VPWR VPWR _32639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26160_ _25013_/X _33493_/Q _26164_/S VGND VGND VPWR VPWR _26161_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35358_ _35744_/CLK _35358_/D VGND VGND VPWR VPWR _35358_/Q sky130_fd_sc_hd__dfxtp_1
X_23372_ _23372_/A VGND VGND VPWR VPWR _32245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1024 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20584_ _33742_/Q _33678_/Q _33614_/Q _33550_/Q _20580_/X _20583_/X VGND VGND VPWR
+ VPWR _20584_/X sky130_fd_sc_hd__mux4_1
X_25111_ _25111_/A VGND VGND VPWR VPWR _33012_/D sky130_fd_sc_hd__clkbuf_1
X_34309_ _34309_/CLK _34309_/D VGND VGND VPWR VPWR _34309_/Q sky130_fd_sc_hd__dfxtp_1
X_22323_ _34301_/Q _34237_/Q _34173_/Q _34109_/Q _22042_/X _22043_/X VGND VGND VPWR
+ VPWR _22323_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26091_ _26091_/A VGND VGND VPWR VPWR _33460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35289_ _36201_/CLK _35289_/D VGND VGND VPWR VPWR _35289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25042_ _25041_/X _32990_/Q _25051_/S VGND VGND VPWR VPWR _25043_/A sky130_fd_sc_hd__mux2_1
X_22254_ _22148_/X _22252_/X _22253_/X _22153_/X VGND VGND VPWR VPWR _22254_/X sky130_fd_sc_hd__a22o_1
XFILLER_152_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21205_ _20957_/X _21203_/X _21204_/X _20961_/X VGND VGND VPWR VPWR _21205_/X sky130_fd_sc_hd__a22o_1
X_29850_ _29850_/A VGND VGND VPWR VPWR _35178_/D sky130_fd_sc_hd__clkbuf_1
X_22185_ _22185_/A VGND VGND VPWR VPWR _36216_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28801_ _26853_/X _34712_/Q _28819_/S VGND VGND VPWR VPWR _28802_/A sky130_fd_sc_hd__mux2_1
X_21136_ _20949_/X _21134_/X _21135_/X _20955_/X VGND VGND VPWR VPWR _21136_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29781_ _35146_/Q _29237_/X _29787_/S VGND VGND VPWR VPWR _29782_/A sky130_fd_sc_hd__mux2_1
X_26993_ input51/X VGND VGND VPWR VPWR _26993_/X sky130_fd_sc_hd__buf_4
XFILLER_232_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_448_CLK clkbuf_6_9__f_CLK/X VGND VGND VPWR VPWR _36001_/CLK sky130_fd_sc_hd__clkbuf_16
X_28732_ _28732_/A VGND VGND VPWR VPWR _34679_/D sky130_fd_sc_hd__clkbuf_1
X_21067_ _33241_/Q _36121_/Q _33113_/Q _33049_/Q _20952_/X _20953_/X VGND VGND VPWR
+ VPWR _21067_/X sky130_fd_sc_hd__mux4_1
X_25944_ _25944_/A VGND VGND VPWR VPWR _33390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20018_ _19807_/X _20016_/X _20017_/X _19812_/X VGND VGND VPWR VPWR _20018_/X sky130_fd_sc_hd__a22o_1
XFILLER_247_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28663_ _26850_/X _34647_/Q _28663_/S VGND VGND VPWR VPWR _28664_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25875_ _26007_/S VGND VGND VPWR VPWR _25894_/S sky130_fd_sc_hd__buf_4
XFILLER_74_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27614_ _27614_/A VGND VGND VPWR VPWR _34149_/D sky130_fd_sc_hd__clkbuf_1
X_24826_ _23034_/X _32896_/Q _24844_/S VGND VGND VPWR VPWR _24827_/A sky130_fd_sc_hd__mux2_1
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28594_ _26946_/X _34614_/Q _28612_/S VGND VGND VPWR VPWR _28595_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27545_ _26996_/X _34118_/Q _27551_/S VGND VGND VPWR VPWR _27546_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21969_ _33779_/Q _33715_/Q _33651_/Q _33587_/Q _21796_/X _21797_/X VGND VGND VPWR
+ VPWR _21969_/X sky130_fd_sc_hd__mux4_1
X_24757_ _24757_/A VGND VGND VPWR VPWR _32863_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23708_ _23708_/A VGND VGND VPWR VPWR _32400_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24688_ _24715_/S VGND VGND VPWR VPWR _24707_/S sky130_fd_sc_hd__clkbuf_8
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27476_ _26894_/X _34085_/Q _27488_/S VGND VGND VPWR VPWR _27477_/A sky130_fd_sc_hd__mux2_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29215_ _29215_/A VGND VGND VPWR VPWR _34882_/D sky130_fd_sc_hd__clkbuf_1
X_26427_ _26427_/A VGND VGND VPWR VPWR _33619_/D sky130_fd_sc_hd__clkbuf_1
X_23639_ _23639_/A VGND VGND VPWR VPWR _32369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29146_ _34860_/Q _29144_/X _29173_/S VGND VGND VPWR VPWR _29147_/A sky130_fd_sc_hd__mux2_1
X_17160_ _17154_/X _17155_/X _17158_/X _17159_/X VGND VGND VPWR VPWR _17160_/X sky130_fd_sc_hd__a22o_1
XFILLER_70_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26358_ _25106_/X _33587_/Q _26362_/S VGND VGND VPWR VPWR _26359_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16111_ _15997_/X _16107_/X _16110_/X _16003_/X VGND VGND VPWR VPWR _16111_/X sky130_fd_sc_hd__a22o_1
XFILLER_196_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25309_ _25309_/A VGND VGND VPWR VPWR _33094_/D sky130_fd_sc_hd__clkbuf_1
X_26289_ _25004_/X _33554_/Q _26299_/S VGND VGND VPWR VPWR _26290_/A sky130_fd_sc_hd__mux2_1
X_29077_ _34838_/Q _29076_/X _29080_/S VGND VGND VPWR VPWR _29078_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17091_ _34283_/Q _34219_/Q _34155_/Q _34091_/Q _17089_/X _17090_/X VGND VGND VPWR
+ VPWR _17091_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16042_ _17843_/A VGND VGND VPWR VPWR _16042_/X sky130_fd_sc_hd__buf_2
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28028_ _26909_/X _34346_/Q _28030_/S VGND VGND VPWR VPWR _28029_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19801_ _19796_/X _19799_/X _19800_/X VGND VGND VPWR VPWR _19816_/C sky130_fd_sc_hd__o21ba_1
XFILLER_151_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17993_ _17989_/X _17992_/X _17853_/X VGND VGND VPWR VPWR _18003_/C sky130_fd_sc_hd__o21ba_1
X_29979_ _29979_/A VGND VGND VPWR VPWR _35239_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_439_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _36135_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_1103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19732_ _34804_/Q _34740_/Q _34676_/Q _34612_/Q _19588_/X _19589_/X VGND VGND VPWR
+ VPWR _19732_/X sky130_fd_sc_hd__mux4_1
X_16944_ _16944_/A _16944_/B _16944_/C _16944_/D VGND VGND VPWR VPWR _16945_/A sky130_fd_sc_hd__or4_4
XFILLER_96_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32990_ _35481_/CLK _32990_/D VGND VGND VPWR VPWR _32990_/Q sky130_fd_sc_hd__dfxtp_1
X_31941_ _31941_/A VGND VGND VPWR VPWR _36169_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19663_ _34546_/Q _32434_/Q _34418_/Q _34354_/Q _19525_/X _19526_/X VGND VGND VPWR
+ VPWR _19663_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16875_ _35044_/Q _34980_/Q _34916_/Q _34852_/Q _16803_/X _16804_/X VGND VGND VPWR
+ VPWR _16875_/X sky130_fd_sc_hd__mux4_1
XFILLER_231_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18614_ _20146_/A VGND VGND VPWR VPWR _18614_/X sky130_fd_sc_hd__buf_6
XTAP_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34660_ _35928_/CLK _34660_/D VGND VGND VPWR VPWR _34660_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19594_ _35056_/Q _34992_/Q _34928_/Q _34864_/Q _19456_/X _19457_/X VGND VGND VPWR
+ VPWR _19594_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31872_ _31872_/A VGND VGND VPWR VPWR _36136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33611_ _35977_/CLK _33611_/D VGND VGND VPWR VPWR _33611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18545_ _18443_/X _18543_/X _18544_/X _18446_/X VGND VGND VPWR VPWR _18545_/X sky130_fd_sc_hd__a22o_1
X_30823_ _23274_/X _35639_/Q _30839_/S VGND VGND VPWR VPWR _30824_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34591_ _35098_/CLK _34591_/D VGND VGND VPWR VPWR _34591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_40__f_CLK clkbuf_5_20_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_40__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_61_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33542_ _34053_/CLK _33542_/D VGND VGND VPWR VPWR _33542_/Q sky130_fd_sc_hd__dfxtp_1
X_18476_ _18436_/X _18474_/X _18475_/X _18441_/X VGND VGND VPWR VPWR _18476_/X sky130_fd_sc_hd__a22o_1
X_30754_ _30754_/A VGND VGND VPWR VPWR _35606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_380 _36208_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_391 _36209_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17427_ _17931_/A VGND VGND VPWR VPWR _17427_/X sky130_fd_sc_hd__buf_6
X_33473_ _34305_/CLK _33473_/D VGND VGND VPWR VPWR _33473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30685_ _30733_/S VGND VGND VPWR VPWR _30704_/S sky130_fd_sc_hd__buf_6
X_35212_ _35341_/CLK _35212_/D VGND VGND VPWR VPWR _35212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32424_ _34922_/CLK _32424_/D VGND VGND VPWR VPWR _32424_/Q sky130_fd_sc_hd__dfxtp_1
X_17358_ _34802_/Q _34738_/Q _34674_/Q _34610_/Q _17288_/X _17289_/X VGND VGND VPWR
+ VPWR _17358_/X sky130_fd_sc_hd__mux4_1
X_36192_ _36200_/CLK _36192_/D VGND VGND VPWR VPWR _36192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35143_ _35784_/CLK _35143_/D VGND VGND VPWR VPWR _35143_/Q sky130_fd_sc_hd__dfxtp_1
X_16309_ _16309_/A VGND VGND VPWR VPWR _31956_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32355_ _36003_/CLK _32355_/D VGND VGND VPWR VPWR _32355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17289_ _17995_/A VGND VGND VPWR VPWR _17289_/X sky130_fd_sc_hd__buf_4
XFILLER_105_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19028_ _18743_/X _19026_/X _19027_/X _18746_/X VGND VGND VPWR VPWR _19028_/X sky130_fd_sc_hd__a22o_1
X_31306_ _35868_/Q input6/X _31316_/S VGND VGND VPWR VPWR _31307_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35074_ _35075_/CLK _35074_/D VGND VGND VPWR VPWR _35074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32286_ _34781_/CLK _32286_/D VGND VGND VPWR VPWR _32286_/Q sky130_fd_sc_hd__dfxtp_1
X_34025_ _34282_/CLK _34025_/D VGND VGND VPWR VPWR _34025_/Q sky130_fd_sc_hd__dfxtp_1
X_31237_ _31237_/A VGND VGND VPWR VPWR _35835_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31168_ _31168_/A VGND VGND VPWR VPWR _35802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30119_ _35306_/Q _29138_/X _30121_/S VGND VGND VPWR VPWR _30120_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23990_ _23990_/A VGND VGND VPWR VPWR _32533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_1052 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35976_ _35977_/CLK _35976_/D VGND VGND VPWR VPWR _35976_/Q sky130_fd_sc_hd__dfxtp_1
X_31099_ _35770_/Q _29188_/X _31109_/S VGND VGND VPWR VPWR _31100_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22941_ input13/X VGND VGND VPWR VPWR _22941_/X sky130_fd_sc_hd__buf_2
XFILLER_214_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34927_ _35054_/CLK _34927_/D VGND VGND VPWR VPWR _34927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22872_ _22868_/X _22871_/X _22467_/A VGND VGND VPWR VPWR _22873_/D sky130_fd_sc_hd__o21ba_1
XFILLER_216_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25660_ _33257_/Q _24329_/X _25664_/S VGND VGND VPWR VPWR _25661_/A sky130_fd_sc_hd__mux2_1
X_34858_ _34922_/CLK _34858_/D VGND VGND VPWR VPWR _34858_/Q sky130_fd_sc_hd__dfxtp_1
X_24611_ _22920_/X _32795_/Q _24623_/S VGND VGND VPWR VPWR _24612_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21823_ _35310_/Q _35246_/Q _35182_/Q _32302_/Q _21606_/X _21607_/X VGND VGND VPWR
+ VPWR _21823_/X sky130_fd_sc_hd__mux4_1
X_25591_ _33226_/Q _24431_/X _25597_/S VGND VGND VPWR VPWR _25592_/A sky130_fd_sc_hd__mux2_1
X_33809_ _35729_/CLK _33809_/D VGND VGND VPWR VPWR _33809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34789_ _36003_/CLK _34789_/D VGND VGND VPWR VPWR _34789_/Q sky130_fd_sc_hd__dfxtp_1
X_24542_ _23022_/X _32764_/Q _24548_/S VGND VGND VPWR VPWR _24543_/A sky130_fd_sc_hd__mux2_1
X_27330_ _34016_/Q _24301_/X _27332_/S VGND VGND VPWR VPWR _27331_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21754_ _21754_/A VGND VGND VPWR VPWR _21754_/X sky130_fd_sc_hd__buf_4
XFILLER_227_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_964 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20705_ _34255_/Q _34191_/Q _34127_/Q _34063_/Q _20605_/X _20607_/X VGND VGND VPWR
+ VPWR _20705_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27261_ _27261_/A VGND VGND VPWR VPWR _33983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24473_ _22920_/X _32731_/Q _24485_/S VGND VGND VPWR VPWR _24474_/A sky130_fd_sc_hd__mux2_1
X_21685_ _21681_/X _21684_/X _21408_/X VGND VGND VPWR VPWR _21686_/D sky130_fd_sc_hd__o21ba_1
XFILLER_106_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29000_ _29000_/A VGND VGND VPWR VPWR _34806_/D sky130_fd_sc_hd__clkbuf_1
X_23424_ input85/X input84/X VGND VGND VPWR VPWR _31680_/A sky130_fd_sc_hd__nand2b_4
XFILLER_32_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26212_ _26212_/A VGND VGND VPWR VPWR _33517_/D sky130_fd_sc_hd__clkbuf_1
X_20636_ _32974_/Q _32910_/Q _32846_/Q _32782_/Q _20633_/X _20635_/X VGND VGND VPWR
+ VPWR _20636_/X sky130_fd_sc_hd__mux4_1
X_27192_ _27192_/A VGND VGND VPWR VPWR _33950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26143_ _26143_/A VGND VGND VPWR VPWR _33485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23355_ _32237_/Q _23241_/X _23371_/S VGND VGND VPWR VPWR _23356_/A sky130_fd_sc_hd__mux2_1
X_20567_ _35341_/Q _35277_/Q _35213_/Q _32333_/Q _18388_/X _18390_/X VGND VGND VPWR
+ VPWR _20567_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22306_ _35580_/Q _35516_/Q _35452_/Q _35388_/Q _22203_/X _22204_/X VGND VGND VPWR
+ VPWR _22306_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26074_ _25084_/X _33452_/Q _26092_/S VGND VGND VPWR VPWR _26075_/A sky130_fd_sc_hd__mux2_1
X_23286_ input40/X VGND VGND VPWR VPWR _23286_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_106_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20498_ _20494_/X _20497_/X _20142_/A _20143_/A VGND VGND VPWR VPWR _20513_/B sky130_fd_sc_hd__o211a_1
X_29902_ _35203_/Q _29216_/X _29914_/S VGND VGND VPWR VPWR _29903_/A sky130_fd_sc_hd__mux2_1
X_25025_ _25025_/A VGND VGND VPWR VPWR _32984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22237_ _35578_/Q _35514_/Q _35450_/Q _35386_/Q _22203_/X _22204_/X VGND VGND VPWR
+ VPWR _22237_/X sky130_fd_sc_hd__mux4_2
XFILLER_105_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29833_ _35170_/Q _29113_/X _29851_/S VGND VGND VPWR VPWR _29834_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_1147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22168_ _35832_/Q _32210_/Q _35704_/Q _35640_/Q _21913_/X _21914_/X VGND VGND VPWR
+ VPWR _22168_/X sky130_fd_sc_hd__mux4_1
XFILLER_26_1109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21119_ _22312_/A VGND VGND VPWR VPWR _21119_/X sky130_fd_sc_hd__buf_6
XFILLER_43_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29764_ _29764_/A VGND VGND VPWR VPWR _35137_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26976_ _26976_/A VGND VGND VPWR VPWR _33855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22099_ _21952_/X _22097_/X _22098_/X _21955_/X VGND VGND VPWR VPWR _22099_/X sky130_fd_sc_hd__a22o_1
XTAP_6989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28715_ _28715_/A VGND VGND VPWR VPWR _34671_/D sky130_fd_sc_hd__clkbuf_1
X_25927_ _25927_/A VGND VGND VPWR VPWR _33382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29695_ _35105_/Q _29110_/X _29695_/S VGND VGND VPWR VPWR _29696_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_1478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28646_ _28646_/A VGND VGND VPWR VPWR _34638_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16660_ _16656_/X _16659_/X _16455_/X VGND VGND VPWR VPWR _16661_/D sky130_fd_sc_hd__o21ba_1
XFILLER_75_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25858_ _25165_/X _33350_/Q _25864_/S VGND VGND VPWR VPWR _25859_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24809_ _23010_/X _32888_/Q _24823_/S VGND VGND VPWR VPWR _24810_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28577_ _26922_/X _34606_/Q _28591_/S VGND VGND VPWR VPWR _28578_/A sky130_fd_sc_hd__mux2_1
X_16591_ _16591_/A _16591_/B _16591_/C _16591_/D VGND VGND VPWR VPWR _16592_/A sky130_fd_sc_hd__or4_2
X_25789_ _25063_/X _33317_/Q _25801_/S VGND VGND VPWR VPWR _25790_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18330_ _20070_/A VGND VGND VPWR VPWR _20163_/A sky130_fd_sc_hd__buf_4
X_27528_ _26971_/X _34110_/Q _27530_/S VGND VGND VPWR VPWR _27529_/A sky130_fd_sc_hd__mux2_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ _15977_/X _18259_/X _18260_/X _15987_/X VGND VGND VPWR VPWR _18261_/X sky130_fd_sc_hd__a22o_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27459_ _26869_/X _34077_/Q _27467_/S VGND VGND VPWR VPWR _27460_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17212_ _33006_/Q _32942_/Q _32878_/Q _32814_/Q _16989_/X _16990_/X VGND VGND VPWR
+ VPWR _17212_/X sky130_fd_sc_hd__mux4_1
X_30470_ _30470_/A VGND VGND VPWR VPWR _35471_/D sky130_fd_sc_hd__clkbuf_1
X_18192_ _32779_/Q _32715_/Q _32651_/Q _36107_/Q _17978_/X _16873_/A VGND VGND VPWR
+ VPWR _18192_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17143_ _16994_/X _17139_/X _17142_/X _16997_/X VGND VGND VPWR VPWR _17143_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29129_ input18/X VGND VGND VPWR VPWR _29129_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_144_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32140_ _35815_/CLK _32140_/D VGND VGND VPWR VPWR _32140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17074_ _17931_/A VGND VGND VPWR VPWR _17074_/X sky130_fd_sc_hd__buf_6
XFILLER_7_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16025_ _17769_/A VGND VGND VPWR VPWR _17908_/A sky130_fd_sc_hd__buf_12
X_32071_ _32518_/CLK _32071_/D VGND VGND VPWR VPWR _32071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31022_ _31022_/A VGND VGND VPWR VPWR _35733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35830_ _35831_/CLK _35830_/D VGND VGND VPWR VPWR _35830_/Q sky130_fd_sc_hd__dfxtp_1
X_17976_ _17908_/X _17974_/X _17975_/X _17911_/X VGND VGND VPWR VPWR _17976_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_900 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19715_ _19708_/X _19710_/X _19713_/X _19714_/X VGND VGND VPWR VPWR _19715_/X sky130_fd_sc_hd__a22o_1
X_16927_ _16922_/X _16926_/X _16783_/X _16784_/X VGND VGND VPWR VPWR _16944_/B sky130_fd_sc_hd__o211a_1
X_32973_ _36045_/CLK _32973_/D VGND VGND VPWR VPWR _32973_/Q sky130_fd_sc_hd__dfxtp_1
X_35761_ _35953_/CLK _35761_/D VGND VGND VPWR VPWR _35761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1083 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31924_ _23307_/X _36161_/Q _31940_/S VGND VGND VPWR VPWR _31925_/A sky130_fd_sc_hd__mux2_1
X_19646_ _19640_/X _19645_/X _19436_/X _19437_/X VGND VGND VPWR VPWR _19667_/B sky130_fd_sc_hd__o211a_1
X_34712_ _34777_/CLK _34712_/D VGND VGND VPWR VPWR _34712_/Q sky130_fd_sc_hd__dfxtp_1
X_35692_ _35885_/CLK _35692_/D VGND VGND VPWR VPWR _35692_/Q sky130_fd_sc_hd__dfxtp_1
X_16858_ _32484_/Q _32356_/Q _32036_/Q _36004_/Q _16570_/X _16711_/X VGND VGND VPWR
+ VPWR _16858_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1029 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34643_ _36189_/CLK _34643_/D VGND VGND VPWR VPWR _34643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19577_ _32496_/Q _32368_/Q _32048_/Q _36016_/Q _19576_/X _19364_/X VGND VGND VPWR
+ VPWR _19577_/X sky130_fd_sc_hd__mux4_1
X_31855_ _31855_/A VGND VGND VPWR VPWR _36128_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16789_ _35746_/Q _35106_/Q _34466_/Q _33826_/Q _16787_/X _16788_/X VGND VGND VPWR
+ VPWR _16789_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18528_ _18524_/X _18527_/X _18371_/X VGND VGND VPWR VPWR _18538_/C sky130_fd_sc_hd__o21ba_1
X_30806_ _23247_/X _35631_/Q _30818_/S VGND VGND VPWR VPWR _30807_/A sky130_fd_sc_hd__mux2_1
X_34574_ _35280_/CLK _34574_/D VGND VGND VPWR VPWR _34574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31786_ _31813_/S VGND VGND VPWR VPWR _31805_/S sky130_fd_sc_hd__buf_6
XFILLER_222_964 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_896 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33525_ _34292_/CLK _33525_/D VGND VGND VPWR VPWR _33525_/Q sky130_fd_sc_hd__dfxtp_1
X_30737_ _23077_/X _35598_/Q _30755_/S VGND VGND VPWR VPWR _30738_/A sky130_fd_sc_hd__mux2_1
X_18459_ _35536_/Q _35472_/Q _35408_/Q _35344_/Q _18358_/X _18360_/X VGND VGND VPWR
+ VPWR _18459_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33456_ _33520_/CLK _33456_/D VGND VGND VPWR VPWR _33456_/Q sky130_fd_sc_hd__dfxtp_1
X_21470_ _35300_/Q _35236_/Q _35172_/Q _32292_/Q _21253_/X _21254_/X VGND VGND VPWR
+ VPWR _21470_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30668_ _30668_/A VGND VGND VPWR VPWR _35565_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20421_ _20160_/X _20419_/X _20420_/X _20165_/X VGND VGND VPWR VPWR _20421_/X sky130_fd_sc_hd__a22o_1
X_32407_ _36189_/CLK _32407_/D VGND VGND VPWR VPWR _32407_/Q sky130_fd_sc_hd__dfxtp_1
X_36175_ _36185_/CLK _36175_/D VGND VGND VPWR VPWR _36175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33387_ _33512_/CLK _33387_/D VGND VGND VPWR VPWR _33387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30599_ _30599_/A VGND VGND VPWR VPWR _35533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35126_ _35766_/CLK _35126_/D VGND VGND VPWR VPWR _35126_/Q sky130_fd_sc_hd__dfxtp_1
X_23140_ _32159_/Q _23139_/X _23146_/S VGND VGND VPWR VPWR _23141_/A sky130_fd_sc_hd__mux2_1
X_20352_ _35590_/Q _35526_/Q _35462_/Q _35398_/Q _20256_/X _20257_/X VGND VGND VPWR
+ VPWR _20352_/X sky130_fd_sc_hd__mux4_1
X_32338_ _36052_/CLK _32338_/D VGND VGND VPWR VPWR _32338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23071_ input59/X VGND VGND VPWR VPWR _23071_/X sky130_fd_sc_hd__clkbuf_4
X_35057_ _35954_/CLK _35057_/D VGND VGND VPWR VPWR _35057_/Q sky130_fd_sc_hd__dfxtp_1
X_20283_ _32516_/Q _32388_/Q _32068_/Q _36036_/Q _20282_/X _20070_/X VGND VGND VPWR
+ VPWR _20283_/X sky130_fd_sc_hd__mux4_1
X_32269_ _34316_/CLK _32269_/D VGND VGND VPWR VPWR _32269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34008_ _35284_/CLK _34008_/D VGND VGND VPWR VPWR _34008_/Q sky130_fd_sc_hd__dfxtp_1
X_22022_ _22015_/X _22021_/X _21736_/X _21737_/X VGND VGND VPWR VPWR _22039_/B sky130_fd_sc_hd__o211a_1
XTAP_6219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26830_ _26829_/X _33808_/Q _26851_/S VGND VGND VPWR VPWR _26831_/A sky130_fd_sc_hd__mux2_1
XTAP_5518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26761_ _33777_/Q _24354_/X _26769_/S VGND VGND VPWR VPWR _26762_/A sky130_fd_sc_hd__mux2_1
X_23973_ _30465_/B _31410_/A VGND VGND VPWR VPWR _24106_/S sky130_fd_sc_hd__nand2_8
XTAP_4839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35959_ _36023_/CLK _35959_/D VGND VGND VPWR VPWR _35959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28500_ _27008_/X _34570_/Q _28506_/S VGND VGND VPWR VPWR _28501_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25712_ _25712_/A VGND VGND VPWR VPWR _33281_/D sky130_fd_sc_hd__clkbuf_1
X_29480_ _23286_/X _35003_/Q _29488_/S VGND VGND VPWR VPWR _29481_/A sky130_fd_sc_hd__mux2_1
X_22924_ _22923_/X _32028_/Q _22939_/S VGND VGND VPWR VPWR _22925_/A sky130_fd_sc_hd__mux2_1
X_26692_ _33744_/Q _24252_/X _26706_/S VGND VGND VPWR VPWR _26693_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28431_ _26906_/X _34537_/Q _28435_/S VGND VGND VPWR VPWR _28432_/A sky130_fd_sc_hd__mux2_1
X_25643_ _33249_/Q _24304_/X _25643_/S VGND VGND VPWR VPWR _25644_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22855_ _32525_/Q _32397_/Q _32077_/Q _36045_/Q _22582_/X _21607_/A VGND VGND VPWR
+ VPWR _22855_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28362_ _28362_/A VGND VGND VPWR VPWR _34504_/D sky130_fd_sc_hd__clkbuf_1
X_21806_ _21802_/X _21803_/X _21804_/X _21805_/X VGND VGND VPWR VPWR _21806_/X sky130_fd_sc_hd__a22o_1
X_22786_ _34315_/Q _34251_/Q _34187_/Q _34123_/Q _20645_/X _20646_/X VGND VGND VPWR
+ VPWR _22786_/X sky130_fd_sc_hd__mux4_1
X_25574_ _25574_/A VGND VGND VPWR VPWR _33217_/D sky130_fd_sc_hd__clkbuf_1
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27313_ _27424_/S VGND VGND VPWR VPWR _27332_/S sky130_fd_sc_hd__clkbuf_8
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21737_ _22443_/A VGND VGND VPWR VPWR _21737_/X sky130_fd_sc_hd__clkbuf_4
X_24525_ _22997_/X _32756_/Q _24527_/S VGND VGND VPWR VPWR _24526_/A sky130_fd_sc_hd__mux2_1
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28293_ _28293_/A VGND VGND VPWR VPWR _34471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27244_ _26950_/X _33975_/Q _27260_/S VGND VGND VPWR VPWR _27245_/A sky130_fd_sc_hd__mux2_1
X_24456_ _22895_/X _32723_/Q _24464_/S VGND VGND VPWR VPWR _24457_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21668_ _21663_/X _21665_/X _21666_/X _21667_/X VGND VGND VPWR VPWR _21668_/X sky130_fd_sc_hd__a22o_1
XFILLER_229_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23407_ _32262_/Q _23322_/X _23413_/S VGND VGND VPWR VPWR _23408_/A sky130_fd_sc_hd__mux2_1
X_20619_ _32718_/Q _32654_/Q _32590_/Q _36046_/Q _22462_/A _22313_/A VGND VGND VPWR
+ VPWR _20619_/X sky130_fd_sc_hd__mux4_1
X_27175_ _27175_/A VGND VGND VPWR VPWR _33942_/D sky130_fd_sc_hd__clkbuf_1
X_24387_ _24387_/A VGND VGND VPWR VPWR _32699_/D sky130_fd_sc_hd__clkbuf_1
X_21599_ _22460_/A VGND VGND VPWR VPWR _21599_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23338_ _23338_/A VGND VGND VPWR VPWR _32230_/D sky130_fd_sc_hd__clkbuf_1
X_26126_ _25162_/X _33477_/Q _26134_/S VGND VGND VPWR VPWR _26127_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26057_ _25060_/X _33444_/Q _26071_/S VGND VGND VPWR VPWR _26058_/A sky130_fd_sc_hd__mux2_1
X_23269_ _23269_/A VGND VGND VPWR VPWR _32207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_4__f_CLK clkbuf_5_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_4__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_25008_ _25007_/X _32979_/Q _25020_/S VGND VGND VPWR VPWR _25009_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17830_ _17830_/A VGND VGND VPWR VPWR _17830_/X sky130_fd_sc_hd__clkbuf_4
X_29816_ _35162_/Q _29089_/X _29830_/S VGND VGND VPWR VPWR _29817_/A sky130_fd_sc_hd__mux2_1
XTAP_6753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17761_ _17761_/A VGND VGND VPWR VPWR _17761_/X sky130_fd_sc_hd__clkbuf_4
X_29747_ _29747_/A VGND VGND VPWR VPWR _35129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26959_ input39/X VGND VGND VPWR VPWR _26959_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_134_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19500_ _20206_/A VGND VGND VPWR VPWR _19500_/X sky130_fd_sc_hd__buf_2
X_16712_ _32480_/Q _32352_/Q _32032_/Q _36000_/Q _16570_/X _16711_/X VGND VGND VPWR
+ VPWR _16712_/X sky130_fd_sc_hd__mux4_1
XFILLER_247_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17692_ _33276_/Q _36156_/Q _33148_/Q _33084_/Q _17411_/X _17412_/X VGND VGND VPWR
+ VPWR _17692_/X sky130_fd_sc_hd__mux4_1
X_29678_ _29678_/A VGND VGND VPWR VPWR _35096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19431_ _33260_/Q _36140_/Q _33132_/Q _33068_/Q _19358_/X _19359_/X VGND VGND VPWR
+ VPWR _19431_/X sky130_fd_sc_hd__mux4_1
X_28629_ _26999_/X _34631_/Q _28633_/S VGND VGND VPWR VPWR _28630_/A sky130_fd_sc_hd__mux2_1
X_16643_ _35742_/Q _35102_/Q _34462_/Q _33822_/Q _16434_/X _16435_/X VGND VGND VPWR
+ VPWR _16643_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31640_ _31640_/A VGND VGND VPWR VPWR _36026_/D sky130_fd_sc_hd__clkbuf_1
X_19362_ _19355_/X _19357_/X _19360_/X _19361_/X VGND VGND VPWR VPWR _19362_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16574_ _16569_/X _16573_/X _16430_/X _16431_/X VGND VGND VPWR VPWR _16591_/B sky130_fd_sc_hd__o211a_2
XFILLER_203_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18313_ _20061_/A VGND VGND VPWR VPWR _20201_/A sky130_fd_sc_hd__buf_12
XFILLER_128_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1035 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31571_ _31571_/A VGND VGND VPWR VPWR _35993_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19293_ _19287_/X _19292_/X _19083_/X _19084_/X VGND VGND VPWR VPWR _19314_/B sky130_fd_sc_hd__o211a_1
XFILLER_188_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33310_ _33946_/CLK _33310_/D VGND VGND VPWR VPWR _33310_/Q sky130_fd_sc_hd__dfxtp_1
X_18244_ _18244_/A VGND VGND VPWR VPWR _32012_/D sky130_fd_sc_hd__clkbuf_1
X_30522_ _30522_/A VGND VGND VPWR VPWR _35496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34290_ _34291_/CLK _34290_/D VGND VGND VPWR VPWR _34290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33241_ _36059_/CLK _33241_/D VGND VGND VPWR VPWR _33241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18175_ _18171_/X _18174_/X _17853_/A VGND VGND VPWR VPWR _18183_/C sky130_fd_sc_hd__o21ba_1
X_30453_ _23330_/X _35464_/Q _30455_/S VGND VGND VPWR VPWR _30454_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17126_ _34028_/Q _33964_/Q _33900_/Q _32236_/Q _17020_/X _17021_/X VGND VGND VPWR
+ VPWR _17126_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33172_ _36115_/CLK _33172_/D VGND VGND VPWR VPWR _33172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30384_ _23220_/X _35431_/Q _30392_/S VGND VGND VPWR VPWR _30385_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32123_ _35562_/CLK _32123_/D VGND VGND VPWR VPWR _32123_/Q sky130_fd_sc_hd__dfxtp_1
X_17057_ _32746_/Q _32682_/Q _32618_/Q _36074_/Q _16919_/X _17056_/X VGND VGND VPWR
+ VPWR _17057_/X sky130_fd_sc_hd__mux4_1
XFILLER_217_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16008_ _33998_/Q _33934_/Q _33870_/Q _32142_/Q _16005_/X _16007_/X VGND VGND VPWR
+ VPWR _16008_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32054_ _36022_/CLK _32054_/D VGND VGND VPWR VPWR _32054_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31005_ _31275_/B _31140_/B VGND VGND VPWR VPWR _31138_/S sky130_fd_sc_hd__nor2_8
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35813_ _35814_/CLK _35813_/D VGND VGND VPWR VPWR _35813_/Q sky130_fd_sc_hd__dfxtp_1
X_17959_ _33219_/Q _32579_/Q _35971_/Q _35907_/Q _17780_/X _17781_/X VGND VGND VPWR
+ VPWR _17959_/X sky130_fd_sc_hd__mux4_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32956_ _36092_/CLK _32956_/D VGND VGND VPWR VPWR _32956_/Q sky130_fd_sc_hd__dfxtp_1
X_20970_ _33174_/Q _32534_/Q _35926_/Q _35862_/Q _20968_/X _20969_/X VGND VGND VPWR
+ VPWR _20970_/X sky130_fd_sc_hd__mux4_1
X_35744_ _35744_/CLK _35744_/D VGND VGND VPWR VPWR _35744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31907_ _23280_/X _36153_/Q _31919_/S VGND VGND VPWR VPWR _31908_/A sky130_fd_sc_hd__mux2_1
X_19629_ _19629_/A _19629_/B _19629_/C _19629_/D VGND VGND VPWR VPWR _19630_/A sky130_fd_sc_hd__or4_1
XFILLER_65_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32887_ _36024_/CLK _32887_/D VGND VGND VPWR VPWR _32887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35675_ _35675_/CLK _35675_/D VGND VGND VPWR VPWR _35675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22640_ _22508_/X _22638_/X _22639_/X _22511_/X VGND VGND VPWR VPWR _22640_/X sky130_fd_sc_hd__a22o_1
X_34626_ _35331_/CLK _34626_/D VGND VGND VPWR VPWR _34626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31838_ _23117_/X _36120_/Q _31856_/S VGND VGND VPWR VPWR _31839_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22571_ _33796_/Q _33732_/Q _33668_/Q _33604_/Q _22502_/X _22503_/X VGND VGND VPWR
+ VPWR _22571_/X sky130_fd_sc_hd__mux4_1
XFILLER_210_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34557_ _34620_/CLK _34557_/D VGND VGND VPWR VPWR _34557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31769_ _31769_/A VGND VGND VPWR VPWR _36087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21522_ _21302_/X _21520_/X _21521_/X _21308_/X VGND VGND VPWR VPWR _21522_/X sky130_fd_sc_hd__a22o_1
X_24310_ _24310_/A VGND VGND VPWR VPWR _32674_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25290_ _25290_/A VGND VGND VPWR VPWR _33085_/D sky130_fd_sc_hd__clkbuf_1
X_33508_ _33702_/CLK _33508_/D VGND VGND VPWR VPWR _33508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34488_ _35766_/CLK _34488_/D VGND VGND VPWR VPWR _34488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24241_ _24241_/A VGND VGND VPWR VPWR _32652_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36227_ _36228_/CLK _36227_/D VGND VGND VPWR VPWR _36227_/Q sky130_fd_sc_hd__dfxtp_1
X_21453_ _21449_/X _21450_/X _21451_/X _21452_/X VGND VGND VPWR VPWR _21453_/X sky130_fd_sc_hd__a22o_1
X_33439_ _33692_/CLK _33439_/D VGND VGND VPWR VPWR _33439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20404_ _19449_/A _20402_/X _20403_/X _19452_/A VGND VGND VPWR VPWR _20404_/X sky130_fd_sc_hd__a22o_1
XFILLER_181_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36158_ _36161_/CLK _36158_/D VGND VGND VPWR VPWR _36158_/Q sky130_fd_sc_hd__dfxtp_1
X_24172_ _24172_/A VGND VGND VPWR VPWR _32619_/D sky130_fd_sc_hd__clkbuf_1
X_21384_ _22443_/A VGND VGND VPWR VPWR _21384_/X sky130_fd_sc_hd__clkbuf_4
X_23123_ _23123_/A VGND VGND VPWR VPWR _32153_/D sky130_fd_sc_hd__clkbuf_1
X_20335_ _33798_/Q _33734_/Q _33670_/Q _33606_/Q _20202_/X _20203_/X VGND VGND VPWR
+ VPWR _20335_/X sky130_fd_sc_hd__mux4_1
X_35109_ _35749_/CLK _35109_/D VGND VGND VPWR VPWR _35109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36089_ _36089_/CLK _36089_/D VGND VGND VPWR VPWR _36089_/Q sky130_fd_sc_hd__dfxtp_1
X_28980_ _34797_/Q _24342_/X _28996_/S VGND VGND VPWR VPWR _28981_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23054_ _23053_/X _32070_/Q _23063_/S VGND VGND VPWR VPWR _23055_/A sky130_fd_sc_hd__mux2_1
XTAP_6005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27931_ _34300_/Q _24388_/X _27937_/S VGND VGND VPWR VPWR _27932_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20266_ _35075_/Q _35011_/Q _34947_/Q _34883_/Q _20162_/X _20163_/X VGND VGND VPWR
+ VPWR _20266_/X sky130_fd_sc_hd__mux4_1
XFILLER_227_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22005_ _34036_/Q _33972_/Q _33908_/Q _32244_/Q _21973_/X _21974_/X VGND VGND VPWR
+ VPWR _22005_/X sky130_fd_sc_hd__mux4_1
XTAP_6049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27862_ _34267_/Q _24286_/X _27874_/S VGND VGND VPWR VPWR _27863_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20197_ _20160_/X _20195_/X _20196_/X _20165_/X VGND VGND VPWR VPWR _20197_/X sky130_fd_sc_hd__a22o_1
XTAP_5326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29601_ _29601_/A VGND VGND VPWR VPWR _35060_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26813_ _33802_/Q _24431_/X _26819_/S VGND VGND VPWR VPWR _26814_/A sky130_fd_sc_hd__mux2_1
XTAP_5348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27793_ _27793_/A VGND VGND VPWR VPWR _34234_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29532_ _29532_/A VGND VGND VPWR VPWR _35027_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26744_ _33769_/Q _24329_/X _26748_/S VGND VGND VPWR VPWR _26745_/A sky130_fd_sc_hd__mux2_1
X_23956_ _23053_/X _32518_/Q _23962_/S VGND VGND VPWR VPWR _23957_/A sky130_fd_sc_hd__mux2_1
XTAP_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22907_ input64/X VGND VGND VPWR VPWR _22907_/X sky130_fd_sc_hd__buf_4
XANTENNA_902 _26277_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29463_ _23261_/X _34995_/Q _29467_/S VGND VGND VPWR VPWR _29464_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26675_ _25174_/X _33737_/Q _26675_/S VGND VGND VPWR VPWR _26676_/A sky130_fd_sc_hd__mux2_1
XTAP_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_913 _26919_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_924 _27424_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23887_ _22951_/X _32485_/Q _23899_/S VGND VGND VPWR VPWR _23888_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_935 _29061_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28414_ _26881_/X _34529_/Q _28414_/S VGND VGND VPWR VPWR _28415_/A sky130_fd_sc_hd__mux2_1
X_25626_ _25626_/A VGND VGND VPWR VPWR _33240_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_946 _29517_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22838_ _20644_/X _22836_/X _22837_/X _20654_/X VGND VGND VPWR VPWR _22838_/X sky130_fd_sc_hd__a22o_1
X_29394_ _23099_/X _34962_/Q _29404_/S VGND VGND VPWR VPWR _29395_/A sky130_fd_sc_hd__mux2_1
XANTENNA_957 _29922_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_968 _31273_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_979 _17855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28345_ _34496_/Q _24400_/X _28363_/S VGND VGND VPWR VPWR _28346_/A sky130_fd_sc_hd__mux2_1
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25557_ _25557_/A VGND VGND VPWR VPWR _33209_/D sky130_fd_sc_hd__clkbuf_1
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22769_ _35850_/Q _32230_/Q _35722_/Q _35658_/Q _20589_/X _20591_/X VGND VGND VPWR
+ VPWR _22769_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24508_ _24577_/S VGND VGND VPWR VPWR _24527_/S sky130_fd_sc_hd__buf_6
X_16290_ _35732_/Q _35092_/Q _34452_/Q _33812_/Q _16049_/X _16051_/X VGND VGND VPWR
+ VPWR _16290_/X sky130_fd_sc_hd__mux4_1
X_28276_ _28276_/A VGND VGND VPWR VPWR _34463_/D sky130_fd_sc_hd__clkbuf_1
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25488_ _25488_/A VGND VGND VPWR VPWR _33176_/D sky130_fd_sc_hd__clkbuf_1
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27227_ _26925_/X _33967_/Q _27239_/S VGND VGND VPWR VPWR _27228_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24439_ _24439_/A VGND VGND VPWR VPWR _32716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27158_ _26821_/X _33934_/Q _27176_/S VGND VGND VPWR VPWR _27159_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26109_ _25137_/X _33469_/Q _26113_/S VGND VGND VPWR VPWR _26110_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19980_ _19807_/X _19978_/X _19979_/X _19812_/X VGND VGND VPWR VPWR _19980_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27089_ _27089_/A VGND VGND VPWR VPWR _33901_/D sky130_fd_sc_hd__clkbuf_1
X_18931_ _18927_/X _18930_/X _18722_/X VGND VGND VPWR VPWR _18961_/A sky130_fd_sc_hd__o21ba_1
XFILLER_98_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1301 _16496_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1312 input11/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1323 _31993_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18862_ _33500_/Q _33436_/Q _33372_/Q _33308_/Q _18717_/X _18718_/X VGND VGND VPWR
+ VPWR _18862_/X sky130_fd_sc_hd__mux4_1
XTAP_6550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1334 _20165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1345 _22462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1356 _22511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17813_ _35583_/Q _35519_/Q _35455_/Q _35391_/Q _17603_/X _17604_/X VGND VGND VPWR
+ VPWR _17813_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1367 _24354_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1378 _26872_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18793_ _34266_/Q _34202_/Q _34138_/Q _34074_/Q _18683_/X _18684_/X VGND VGND VPWR
+ VPWR _18793_/X sky130_fd_sc_hd__mux4_1
XTAP_5860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1389 _17830_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32810_ _36075_/CLK _32810_/D VGND VGND VPWR VPWR _32810_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17744_ _17740_/X _17743_/X _17500_/X VGND VGND VPWR VPWR _17752_/C sky130_fd_sc_hd__o21ba_1
XFILLER_208_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33790_ _34303_/CLK _33790_/D VGND VGND VPWR VPWR _33790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32741_ _36070_/CLK _32741_/D VGND VGND VPWR VPWR _32741_/Q sky130_fd_sc_hd__dfxtp_1
X_17675_ _34811_/Q _34747_/Q _34683_/Q _34619_/Q _17641_/X _17642_/X VGND VGND VPWR
+ VPWR _17675_/X sky130_fd_sc_hd__mux4_1
XFILLER_247_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19414_ _34539_/Q _32427_/Q _34411_/Q _34347_/Q _19172_/X _19173_/X VGND VGND VPWR
+ VPWR _19414_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35460_ _35973_/CLK _35460_/D VGND VGND VPWR VPWR _35460_/Q sky130_fd_sc_hd__dfxtp_1
X_16626_ _34270_/Q _34206_/Q _34142_/Q _34078_/Q _16383_/X _16384_/X VGND VGND VPWR
+ VPWR _16626_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_917 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32672_ _36128_/CLK _32672_/D VGND VGND VPWR VPWR _32672_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34411_ _35050_/CLK _34411_/D VGND VGND VPWR VPWR _34411_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_10_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_10_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_19345_ _19341_/X _19344_/X _19108_/X VGND VGND VPWR VPWR _19346_/D sky130_fd_sc_hd__o21ba_1
X_31623_ _31623_/A VGND VGND VPWR VPWR _36018_/D sky130_fd_sc_hd__clkbuf_1
X_35391_ _36105_/CLK _35391_/D VGND VGND VPWR VPWR _35391_/Q sky130_fd_sc_hd__dfxtp_1
X_16557_ _16557_/A _16557_/B _16557_/C _16557_/D VGND VGND VPWR VPWR _16558_/A sky130_fd_sc_hd__or4_2
XFILLER_188_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34342_ _35942_/CLK _34342_/D VGND VGND VPWR VPWR _34342_/Q sky130_fd_sc_hd__dfxtp_1
X_31554_ _31554_/A VGND VGND VPWR VPWR _35985_/D sky130_fd_sc_hd__clkbuf_1
X_19276_ _19276_/A _19276_/B _19276_/C _19276_/D VGND VGND VPWR VPWR _19277_/A sky130_fd_sc_hd__or4_4
XFILLER_203_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16488_ _16488_/A VGND VGND VPWR VPWR _31961_/D sky130_fd_sc_hd__clkbuf_1
X_18227_ _17154_/A _18225_/X _18226_/X _17159_/A VGND VGND VPWR VPWR _18227_/X sky130_fd_sc_hd__a22o_1
X_30505_ _30505_/A VGND VGND VPWR VPWR _35488_/D sky130_fd_sc_hd__clkbuf_1
X_34273_ _36123_/CLK _34273_/D VGND VGND VPWR VPWR _34273_/Q sky130_fd_sc_hd__dfxtp_1
X_31485_ _23253_/X _35953_/Q _31493_/S VGND VGND VPWR VPWR _31486_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_5_25_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_25_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_117_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36012_ _36013_/CLK _36012_/D VGND VGND VPWR VPWR _36012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33224_ _35977_/CLK _33224_/D VGND VGND VPWR VPWR _33224_/Q sky130_fd_sc_hd__dfxtp_1
X_30436_ _30463_/S VGND VGND VPWR VPWR _30455_/S sky130_fd_sc_hd__buf_4
X_18158_ _33546_/Q _33482_/Q _33418_/Q _33354_/Q _16033_/X _16035_/X VGND VGND VPWR
+ VPWR _18158_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17109_ _16999_/X _17107_/X _17108_/X _17002_/X VGND VGND VPWR VPWR _17109_/X sky130_fd_sc_hd__a22o_1
X_33155_ _36100_/CLK _33155_/D VGND VGND VPWR VPWR _33155_/Q sky130_fd_sc_hd__dfxtp_1
X_18089_ _34567_/Q _32455_/Q _34439_/Q _34375_/Q _17931_/X _17932_/X VGND VGND VPWR
+ VPWR _18089_/X sky130_fd_sc_hd__mux4_1
X_30367_ _23139_/X _35423_/Q _30371_/S VGND VGND VPWR VPWR _30368_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20120_ _34559_/Q _32447_/Q _34431_/Q _34367_/Q _19878_/X _19879_/X VGND VGND VPWR
+ VPWR _20120_/X sky130_fd_sc_hd__mux4_1
X_32106_ _35552_/CLK _32106_/D VGND VGND VPWR VPWR _32106_/Q sky130_fd_sc_hd__dfxtp_1
X_33086_ _34046_/CLK _33086_/D VGND VGND VPWR VPWR _33086_/Q sky130_fd_sc_hd__dfxtp_1
X_30298_ _35391_/Q _29203_/X _30298_/S VGND VGND VPWR VPWR _30299_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20051_ _20047_/X _20050_/X _19814_/X VGND VGND VPWR VPWR _20052_/D sky130_fd_sc_hd__o21ba_1
X_32037_ _36069_/CLK _32037_/D VGND VGND VPWR VPWR _32037_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23810_ _23038_/X _32449_/Q _23826_/S VGND VGND VPWR VPWR _23811_/A sky130_fd_sc_hd__mux2_1
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24790_ _22982_/X _32879_/Q _24802_/S VGND VGND VPWR VPWR _24791_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33988_ _34306_/CLK _33988_/D VGND VGND VPWR VPWR _33988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35727_ _35727_/CLK _35727_/D VGND VGND VPWR VPWR _35727_/Q sky130_fd_sc_hd__dfxtp_1
X_20953_ _22503_/A VGND VGND VPWR VPWR _20953_/X sky130_fd_sc_hd__clkbuf_4
X_23741_ _23741_/A VGND VGND VPWR VPWR _32416_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32939_ _36075_/CLK _32939_/D VGND VGND VPWR VPWR _32939_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26460_ _25057_/X _33635_/Q _26476_/S VGND VGND VPWR VPWR _26461_/A sky130_fd_sc_hd__mux2_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35658_ _35852_/CLK _35658_/D VGND VGND VPWR VPWR _35658_/Q sky130_fd_sc_hd__dfxtp_1
X_23672_ _32385_/Q _23307_/X _23688_/S VGND VGND VPWR VPWR _23673_/A sky130_fd_sc_hd__mux2_1
X_20884_ _22430_/A VGND VGND VPWR VPWR _20884_/X sky130_fd_sc_hd__buf_4
XFILLER_14_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25411_ _25115_/X _33142_/Q _25429_/S VGND VGND VPWR VPWR _25412_/A sky130_fd_sc_hd__mux2_1
X_22623_ _33221_/Q _32581_/Q _35973_/Q _35909_/Q _22380_/X _22381_/X VGND VGND VPWR
+ VPWR _22623_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34609_ _34932_/CLK _34609_/D VGND VGND VPWR VPWR _34609_/Q sky130_fd_sc_hd__dfxtp_1
X_26391_ _26391_/A VGND VGND VPWR VPWR _33602_/D sky130_fd_sc_hd__clkbuf_1
X_35589_ _35973_/CLK _35589_/D VGND VGND VPWR VPWR _35589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28130_ _26860_/X _34394_/Q _28144_/S VGND VGND VPWR VPWR _28131_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22554_ _35779_/Q _35139_/Q _34499_/Q _33859_/Q _22446_/X _22447_/X VGND VGND VPWR
+ VPWR _22554_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25342_ _25342_/A VGND VGND VPWR VPWR _33109_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21505_ _21396_/X _21503_/X _21504_/X _21399_/X VGND VGND VPWR VPWR _21505_/X sky130_fd_sc_hd__a22o_1
X_28061_ _28061_/A VGND VGND VPWR VPWR _34361_/D sky130_fd_sc_hd__clkbuf_1
X_22485_ _35841_/Q _32220_/Q _35713_/Q _35649_/Q _22266_/X _22267_/X VGND VGND VPWR
+ VPWR _22485_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25273_ _25273_/A VGND VGND VPWR VPWR _33077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27012_ _27011_/X _33867_/Q _27018_/S VGND VGND VPWR VPWR _27013_/A sky130_fd_sc_hd__mux2_1
X_24224_ _23047_/X _32644_/Q _24234_/S VGND VGND VPWR VPWR _24225_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21436_ _34531_/Q _32419_/Q _34403_/Q _34339_/Q _21119_/X _21120_/X VGND VGND VPWR
+ VPWR _21436_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_17__f_CLK clkbuf_5_8_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_99_CLK/A sky130_fd_sc_hd__clkbuf_16
X_24155_ _22945_/X _32611_/Q _24171_/S VGND VGND VPWR VPWR _24156_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_190_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _35581_/CLK sky130_fd_sc_hd__clkbuf_16
X_21367_ _33762_/Q _33698_/Q _33634_/Q _33570_/Q _21090_/X _21091_/X VGND VGND VPWR
+ VPWR _21367_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23106_ _32148_/Q _23105_/X _23115_/S VGND VGND VPWR VPWR _23107_/A sky130_fd_sc_hd__mux2_1
X_20318_ _20314_/X _20317_/X _20142_/X _20143_/X VGND VGND VPWR VPWR _20333_/B sky130_fd_sc_hd__o211a_1
X_24086_ _23044_/X _32579_/Q _24098_/S VGND VGND VPWR VPWR _24087_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28963_ _34789_/Q _24317_/X _28975_/S VGND VGND VPWR VPWR _28964_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21298_ _33504_/Q _33440_/Q _33376_/Q _33312_/Q _21017_/X _21018_/X VGND VGND VPWR
+ VPWR _21298_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23037_ _23037_/A VGND VGND VPWR VPWR _32064_/D sky130_fd_sc_hd__clkbuf_1
X_27914_ _34292_/Q _24363_/X _27916_/S VGND VGND VPWR VPWR _27915_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_952 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20249_ _32515_/Q _32387_/Q _32067_/Q _36035_/Q _19929_/X _20070_/X VGND VGND VPWR
+ VPWR _20249_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28894_ _28894_/A VGND VGND VPWR VPWR _34756_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27845_ _34259_/Q _24261_/X _27853_/S VGND VGND VPWR VPWR _27846_/A sky130_fd_sc_hd__mux2_1
XTAP_5145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27776_ _27776_/A VGND VGND VPWR VPWR _34226_/D sky130_fd_sc_hd__clkbuf_1
X_24988_ _24988_/A VGND VGND VPWR VPWR _32973_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_839 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29515_ _23342_/X _35020_/Q _29517_/S VGND VGND VPWR VPWR _29516_/A sky130_fd_sc_hd__mux2_1
XTAP_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26727_ _33761_/Q _24304_/X _26727_/S VGND VGND VPWR VPWR _26728_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23939_ _23028_/X _32510_/Q _23941_/S VGND VGND VPWR VPWR _23940_/A sky130_fd_sc_hd__mux2_1
XTAP_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_710 _22465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_721 _21754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_732 _21157_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29446_ _23234_/X _34987_/Q _29446_/S VGND VGND VPWR VPWR _29447_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17460_ _35573_/Q _35509_/Q _35445_/Q _35381_/Q _17250_/X _17251_/X VGND VGND VPWR
+ VPWR _17460_/X sky130_fd_sc_hd__mux4_1
X_26658_ _26658_/A VGND VGND VPWR VPWR _33728_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_743 _21897_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_754 _22470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_765 _22500_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16411_ _16407_/X _16410_/X _16100_/X VGND VGND VPWR VPWR _16412_/D sky130_fd_sc_hd__o21ba_1
XFILLER_60_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_776 _22603_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25609_ _25609_/A VGND VGND VPWR VPWR _33232_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_787 _22634_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29377_ _29377_/A VGND VGND VPWR VPWR _34954_/D sky130_fd_sc_hd__clkbuf_1
X_17391_ _17387_/X _17390_/X _17147_/X VGND VGND VPWR VPWR _17399_/C sky130_fd_sc_hd__o21ba_1
XANTENNA_798 _22874_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26589_ _25047_/X _33696_/Q _26591_/S VGND VGND VPWR VPWR _26590_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19130_ _33187_/Q _32547_/Q _35939_/Q _35875_/Q _19021_/X _19022_/X VGND VGND VPWR
+ VPWR _19130_/X sky130_fd_sc_hd__mux4_1
X_16342_ _33750_/Q _33686_/Q _33622_/Q _33558_/Q _16137_/X _16138_/X VGND VGND VPWR
+ VPWR _16342_/X sky130_fd_sc_hd__mux4_1
X_28328_ _34488_/Q _24376_/X _28342_/S VGND VGND VPWR VPWR _28329_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19061_ _34529_/Q _32417_/Q _34401_/Q _34337_/Q _18819_/X _18820_/X VGND VGND VPWR
+ VPWR _19061_/X sky130_fd_sc_hd__mux4_1
X_16273_ _34260_/Q _34196_/Q _34132_/Q _34068_/Q _16005_/X _16007_/X VGND VGND VPWR
+ VPWR _16273_/X sky130_fd_sc_hd__mux4_1
X_28259_ _28259_/A VGND VGND VPWR VPWR _34455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18012_ _32773_/Q _32709_/Q _32645_/Q _36101_/Q _17978_/X _17762_/X VGND VGND VPWR
+ VPWR _18012_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31270_ _31270_/A VGND VGND VPWR VPWR _35851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30221_ _35354_/Q _29089_/X _30235_/S VGND VGND VPWR VPWR _30222_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_181_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _35985_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30152_ _30152_/A VGND VGND VPWR VPWR _35321_/D sky130_fd_sc_hd__clkbuf_1
X_19963_ _33019_/Q _32955_/Q _32891_/Q _32827_/Q _19642_/X _19643_/X VGND VGND VPWR
+ VPWR _19963_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18914_ _18593_/X _18912_/X _18913_/X _18596_/X VGND VGND VPWR VPWR _18914_/X sky130_fd_sc_hd__a22o_1
XTAP_7070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1120 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_34960_ _35026_/CLK _34960_/D VGND VGND VPWR VPWR _34960_/Q sky130_fd_sc_hd__dfxtp_1
X_30083_ _30083_/A VGND VGND VPWR VPWR _35288_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19894_ _33273_/Q _36153_/Q _33145_/Q _33081_/Q _19711_/X _19712_/X VGND VGND VPWR
+ VPWR _19894_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1131 _17908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1142 _20158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1153 _22455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33911_ _36152_/CLK _33911_/D VGND VGND VPWR VPWR _33911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18845_ _20257_/A VGND VGND VPWR VPWR _18845_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_41_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1164 _22508_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_34891_ _35788_/CLK _34891_/D VGND VGND VPWR VPWR _34891_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1175 _21757_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1186 _22217_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1197 _22938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33842_ _34997_/CLK _33842_/D VGND VGND VPWR VPWR _33842_/Q sky130_fd_sc_hd__dfxtp_1
X_18776_ _35545_/Q _35481_/Q _35417_/Q _35353_/Q _18491_/X _18492_/X VGND VGND VPWR
+ VPWR _18776_/X sky130_fd_sc_hd__mux4_1
X_15988_ _16057_/A VGND VGND VPWR VPWR _17795_/A sky130_fd_sc_hd__buf_12
XTAP_5690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17727_ _17847_/A VGND VGND VPWR VPWR _17727_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_82_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33773_ _34745_/CLK _33773_/D VGND VGND VPWR VPWR _33773_/Q sky130_fd_sc_hd__dfxtp_1
X_30985_ _35716_/Q _29219_/X _30995_/S VGND VGND VPWR VPWR _30986_/A sky130_fd_sc_hd__mux2_1
XFILLER_209_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35512_ _35638_/CLK _35512_/D VGND VGND VPWR VPWR _35512_/Q sky130_fd_sc_hd__dfxtp_1
X_32724_ _36052_/CLK _32724_/D VGND VGND VPWR VPWR _32724_/Q sky130_fd_sc_hd__dfxtp_1
X_17658_ _17654_/X _17657_/X _17481_/X VGND VGND VPWR VPWR _17682_/A sky130_fd_sc_hd__o21ba_1
XFILLER_23_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16609_ _35805_/Q _32180_/Q _35677_/Q _35613_/Q _16607_/X _16608_/X VGND VGND VPWR
+ VPWR _16609_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32655_ _36048_/CLK _32655_/D VGND VGND VPWR VPWR _32655_/Q sky130_fd_sc_hd__dfxtp_1
X_35443_ _36019_/CLK _35443_/D VGND VGND VPWR VPWR _35443_/Q sky130_fd_sc_hd__dfxtp_1
X_17589_ _33529_/Q _33465_/Q _33401_/Q _33337_/Q _17476_/X _17477_/X VGND VGND VPWR
+ VPWR _17589_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19328_ _32489_/Q _32361_/Q _32041_/Q _36009_/Q _19223_/X _19011_/X VGND VGND VPWR
+ VPWR _19328_/X sky130_fd_sc_hd__mux4_1
X_31606_ _31606_/A VGND VGND VPWR VPWR _36010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32586_ _35978_/CLK _32586_/D VGND VGND VPWR VPWR _32586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35374_ _35562_/CLK _35374_/D VGND VGND VPWR VPWR _35374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31537_ _23336_/X _35978_/Q _31543_/S VGND VGND VPWR VPWR _31538_/A sky130_fd_sc_hd__mux2_1
X_34325_ _36196_/CLK _34325_/D VGND VGND VPWR VPWR _34325_/Q sky130_fd_sc_hd__dfxtp_1
X_19259_ _19255_/X _19258_/X _19083_/X _19084_/X VGND VGND VPWR VPWR _19276_/B sky130_fd_sc_hd__o211a_1
XFILLER_176_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34256_ _34256_/CLK _34256_/D VGND VGND VPWR VPWR _34256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22270_ _21947_/X _22268_/X _22269_/X _21950_/X VGND VGND VPWR VPWR _22270_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_958 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31468_ _23228_/X _35945_/Q _31472_/S VGND VGND VPWR VPWR _31469_/A sky130_fd_sc_hd__mux2_1
X_21221_ _21048_/X _21219_/X _21220_/X _21053_/X VGND VGND VPWR VPWR _21221_/X sky130_fd_sc_hd__a22o_1
X_33207_ _36023_/CLK _33207_/D VGND VGND VPWR VPWR _33207_/Q sky130_fd_sc_hd__dfxtp_1
X_30419_ _30419_/A VGND VGND VPWR VPWR _35447_/D sky130_fd_sc_hd__clkbuf_1
X_34187_ _35851_/CLK _34187_/D VGND VGND VPWR VPWR _34187_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_172_CLK clkbuf_leaf_76_CLK/A VGND VGND VPWR VPWR _34316_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31399_ _31399_/A VGND VGND VPWR VPWR _35912_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33138_ _36146_/CLK _33138_/D VGND VGND VPWR VPWR _33138_/Q sky130_fd_sc_hd__dfxtp_1
X_21152_ _21043_/X _21150_/X _21151_/X _21046_/X VGND VGND VPWR VPWR _21152_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20103_ _32767_/Q _32703_/Q _32639_/Q _36095_/Q _19925_/X _20062_/X VGND VGND VPWR
+ VPWR _20103_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25960_ _25115_/X _33398_/Q _25978_/S VGND VGND VPWR VPWR _25961_/A sky130_fd_sc_hd__mux2_1
X_33069_ _35889_/CLK _33069_/D VGND VGND VPWR VPWR _33069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21083_ _34521_/Q _32409_/Q _34393_/Q _34329_/Q _20766_/X _20767_/X VGND VGND VPWR
+ VPWR _21083_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_972 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20034_ _32509_/Q _32381_/Q _32061_/Q _36029_/Q _19929_/X _19717_/X VGND VGND VPWR
+ VPWR _20034_/X sky130_fd_sc_hd__mux4_1
X_24911_ _24911_/A VGND VGND VPWR VPWR _32936_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25891_ _25891_/A VGND VGND VPWR VPWR _33365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27630_ _34157_/Q _24342_/X _27646_/S VGND VGND VPWR VPWR _27631_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24842_ _23059_/X _32904_/Q _24844_/S VGND VGND VPWR VPWR _24843_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27561_ _31680_/A _27561_/B VGND VGND VPWR VPWR _27562_/A sky130_fd_sc_hd__or2_1
XFILLER_6_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24773_ _22957_/X _32871_/Q _24781_/S VGND VGND VPWR VPWR _24774_/A sky130_fd_sc_hd__mux2_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21985_ _35827_/Q _32205_/Q _35699_/Q _35635_/Q _21913_/X _21914_/X VGND VGND VPWR
+ VPWR _21985_/X sky130_fd_sc_hd__mux4_1
XFILLER_227_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29300_ _29300_/A VGND VGND VPWR VPWR _34917_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26512_ _25134_/X _33660_/Q _26518_/S VGND VGND VPWR VPWR _26513_/A sky130_fd_sc_hd__mux2_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23724_ _22910_/X _32408_/Q _23742_/S VGND VGND VPWR VPWR _23725_/A sky130_fd_sc_hd__mux2_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ _34517_/Q _32405_/Q _34389_/Q _34325_/Q _20766_/X _20767_/X VGND VGND VPWR
+ VPWR _20936_/X sky130_fd_sc_hd__mux4_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27492_ _27492_/A VGND VGND VPWR VPWR _34092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29231_ input54/X VGND VGND VPWR VPWR _29231_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26443_ _25032_/X _33627_/Q _26455_/S VGND VGND VPWR VPWR _26444_/A sky130_fd_sc_hd__mux2_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20867_ _35027_/Q _34963_/Q _34899_/Q _34835_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _20867_/X sky130_fd_sc_hd__mux4_1
X_23655_ _32377_/Q _23280_/X _23667_/S VGND VGND VPWR VPWR _23656_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1019 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22606_ _34309_/Q _34245_/Q _34181_/Q _34117_/Q _22395_/X _22396_/X VGND VGND VPWR
+ VPWR _22606_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29162_ _29162_/A VGND VGND VPWR VPWR _34865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26374_ _26374_/A VGND VGND VPWR VPWR _33594_/D sky130_fd_sc_hd__clkbuf_1
X_20798_ _35281_/Q _35217_/Q _35153_/Q _32273_/Q _20679_/X _20681_/X VGND VGND VPWR
+ VPWR _20798_/X sky130_fd_sc_hd__mux4_1
X_23586_ _32344_/Q _23117_/X _23604_/S VGND VGND VPWR VPWR _23587_/A sky130_fd_sc_hd__mux2_1
X_28113_ _26835_/X _34386_/Q _28123_/S VGND VGND VPWR VPWR _28114_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25325_ _31815_/B _28643_/B VGND VGND VPWR VPWR _25458_/S sky130_fd_sc_hd__nand2_8
XFILLER_128_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22537_ _22537_/A _22537_/B _22537_/C _22537_/D VGND VGND VPWR VPWR _22538_/A sky130_fd_sc_hd__or4_4
XFILLER_224_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29093_ _34843_/Q _29092_/X _29111_/S VGND VGND VPWR VPWR _29094_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28044_ _28044_/A VGND VGND VPWR VPWR _34353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25256_ _25088_/X _33069_/Q _25272_/S VGND VGND VPWR VPWR _25257_/A sky130_fd_sc_hd__mux2_1
X_22468_ _22459_/X _22466_/X _22467_/X VGND VGND VPWR VPWR _22469_/D sky130_fd_sc_hd__o21ba_1
XFILLER_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24207_ _23022_/X _32636_/Q _24213_/S VGND VGND VPWR VPWR _24208_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_163_CLK clkbuf_6_30__f_CLK/X VGND VGND VPWR VPWR _36172_/CLK sky130_fd_sc_hd__clkbuf_16
X_21419_ _32739_/Q _32675_/Q _32611_/Q _36067_/Q _21166_/X _21303_/X VGND VGND VPWR
+ VPWR _21419_/X sky130_fd_sc_hd__mux4_1
X_25187_ _25186_/X _33037_/Q _25187_/S VGND VGND VPWR VPWR _25188_/A sky130_fd_sc_hd__mux2_1
X_22399_ _33535_/Q _33471_/Q _33407_/Q _33343_/Q _22076_/X _22077_/X VGND VGND VPWR
+ VPWR _22399_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24138_ _22920_/X _32603_/Q _24150_/S VGND VGND VPWR VPWR _24139_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29995_ _35247_/Q _29154_/X _30007_/S VGND VGND VPWR VPWR _29996_/A sky130_fd_sc_hd__mux2_1
X_16960_ _17795_/A VGND VGND VPWR VPWR _16960_/X sky130_fd_sc_hd__buf_4
XFILLER_151_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24069_ _23019_/X _32571_/Q _24077_/S VGND VGND VPWR VPWR _24070_/A sky130_fd_sc_hd__mux2_1
X_28946_ _34781_/Q _24292_/X _28954_/S VGND VGND VPWR VPWR _28947_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28877_ _28877_/A VGND VGND VPWR VPWR _34748_/D sky130_fd_sc_hd__clkbuf_1
X_16891_ _32997_/Q _32933_/Q _32869_/Q _32805_/Q _16636_/X _16637_/X VGND VGND VPWR
+ VPWR _16891_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18630_ _33173_/Q _32533_/Q _35925_/Q _35861_/Q _18363_/X _18365_/X VGND VGND VPWR
+ VPWR _18630_/X sky130_fd_sc_hd__mux4_1
X_27828_ _27828_/A VGND VGND VPWR VPWR _34251_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18561_ _18356_/X _18559_/X _18560_/X _18368_/X VGND VGND VPWR VPWR _18561_/X sky130_fd_sc_hd__a22o_1
XTAP_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27759_ _27759_/A VGND VGND VPWR VPWR _34218_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ _17865_/A VGND VGND VPWR VPWR _17512_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18492_ _20147_/A VGND VGND VPWR VPWR _18492_/X sky130_fd_sc_hd__buf_4
XTAP_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30770_ _23136_/X _35614_/Q _30776_/S VGND VGND VPWR VPWR _30771_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_540 _20256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_551 _20142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17443_ _17957_/A VGND VGND VPWR VPWR _17443_/X sky130_fd_sc_hd__buf_4
X_29429_ _29429_/A VGND VGND VPWR VPWR _34978_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_562 _20146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_573 _20165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_584 _19307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_595 _19459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32440_ _35320_/CLK _32440_/D VGND VGND VPWR VPWR _32440_/Q sky130_fd_sc_hd__dfxtp_1
X_17374_ _17847_/A VGND VGND VPWR VPWR _17374_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19113_ _34275_/Q _34211_/Q _34147_/Q _34083_/Q _19036_/X _19037_/X VGND VGND VPWR
+ VPWR _19113_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16325_ _16321_/X _16324_/X _16040_/X _16042_/X VGND VGND VPWR VPWR _16340_/B sky130_fd_sc_hd__o211a_1
XFILLER_41_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32371_ _34222_/CLK _32371_/D VGND VGND VPWR VPWR _32371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34110_ _36157_/CLK _34110_/D VGND VGND VPWR VPWR _34110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31322_ _31322_/A VGND VGND VPWR VPWR _35875_/D sky130_fd_sc_hd__clkbuf_1
X_19044_ _32737_/Q _32673_/Q _32609_/Q _36065_/Q _18866_/X _19003_/X VGND VGND VPWR
+ VPWR _19044_/X sky130_fd_sc_hd__mux4_1
X_35090_ _35729_/CLK _35090_/D VGND VGND VPWR VPWR _35090_/Q sky130_fd_sc_hd__dfxtp_1
X_16256_ _35795_/Q _32169_/Q _35667_/Q _35603_/Q _16254_/X _16255_/X VGND VGND VPWR
+ VPWR _16256_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34041_ _36154_/CLK _34041_/D VGND VGND VPWR VPWR _34041_/Q sky130_fd_sc_hd__dfxtp_1
X_31253_ _35843_/Q input49/X _31265_/S VGND VGND VPWR VPWR _31254_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_154_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _34822_/CLK sky130_fd_sc_hd__clkbuf_16
X_16187_ _16183_/X _16186_/X _16040_/X _16042_/X VGND VGND VPWR VPWR _16204_/B sky130_fd_sc_hd__o211a_1
Xoutput205 _36230_/Q VGND VGND VPWR VPWR D2[56] sky130_fd_sc_hd__buf_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput216 _36182_/Q VGND VGND VPWR VPWR D2[8] sky130_fd_sc_hd__buf_2
X_30204_ _35346_/Q _29064_/X _30214_/S VGND VGND VPWR VPWR _30205_/A sky130_fd_sc_hd__mux2_1
Xoutput227 _32096_/Q VGND VGND VPWR VPWR D3[18] sky130_fd_sc_hd__buf_2
XFILLER_99_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_833 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput238 _32106_/Q VGND VGND VPWR VPWR D3[28] sky130_fd_sc_hd__buf_2
X_31184_ _35810_/Q input13/X _31202_/S VGND VGND VPWR VPWR _31185_/A sky130_fd_sc_hd__mux2_1
Xoutput249 _32116_/Q VGND VGND VPWR VPWR D3[38] sky130_fd_sc_hd__buf_2
XFILLER_88_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_63__f_CLK clkbuf_5_31_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_63__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_142_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30135_ _30135_/A VGND VGND VPWR VPWR _35313_/D sky130_fd_sc_hd__clkbuf_1
X_19946_ _34554_/Q _32442_/Q _34426_/Q _34362_/Q _19878_/X _19879_/X VGND VGND VPWR
+ VPWR _19946_/X sky130_fd_sc_hd__mux4_1
X_35992_ _35992_/CLK _35992_/D VGND VGND VPWR VPWR _35992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30066_ _30066_/A VGND VGND VPWR VPWR _35280_/D sky130_fd_sc_hd__clkbuf_1
X_34943_ _35989_/CLK _34943_/D VGND VGND VPWR VPWR _34943_/Q sky130_fd_sc_hd__dfxtp_1
X_19877_ _19802_/X _19875_/X _19876_/X _19805_/X VGND VGND VPWR VPWR _19877_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18828_ _34267_/Q _34203_/Q _34139_/Q _34075_/Q _18683_/X _18684_/X VGND VGND VPWR
+ VPWR _18828_/X sky130_fd_sc_hd__mux4_1
X_34874_ _35002_/CLK _34874_/D VGND VGND VPWR VPWR _34874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33825_ _35745_/CLK _33825_/D VGND VGND VPWR VPWR _33825_/Q sky130_fd_sc_hd__dfxtp_1
X_18759_ _33753_/Q _33689_/Q _33625_/Q _33561_/Q _18437_/X _18438_/X VGND VGND VPWR
+ VPWR _18759_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21770_ _21449_/X _21768_/X _21769_/X _21452_/X VGND VGND VPWR VPWR _21770_/X sky130_fd_sc_hd__a22o_1
X_30968_ _35708_/Q _29194_/X _30974_/S VGND VGND VPWR VPWR _30969_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33756_ _34017_/CLK _33756_/D VGND VGND VPWR VPWR _33756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20721_ _35727_/Q _35087_/Q _34447_/Q _33807_/Q _20649_/X _20651_/X VGND VGND VPWR
+ VPWR _20721_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32707_ _36100_/CLK _32707_/D VGND VGND VPWR VPWR _32707_/Q sky130_fd_sc_hd__dfxtp_1
X_33687_ _35664_/CLK _33687_/D VGND VGND VPWR VPWR _33687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30899_ _35675_/Q _29092_/X _30911_/S VGND VGND VPWR VPWR _30900_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20652_ _35726_/Q _35086_/Q _34446_/Q _33806_/Q _20649_/X _20651_/X VGND VGND VPWR
+ VPWR _20652_/X sky130_fd_sc_hd__mux4_1
X_23440_ _22898_/X _32276_/Q _23446_/S VGND VGND VPWR VPWR _23441_/A sky130_fd_sc_hd__mux2_1
X_35426_ _35940_/CLK _35426_/D VGND VGND VPWR VPWR _35426_/Q sky130_fd_sc_hd__dfxtp_1
X_32638_ _32959_/CLK _32638_/D VGND VGND VPWR VPWR _32638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23371_ _32245_/Q _23267_/X _23371_/S VGND VGND VPWR VPWR _23372_/A sky130_fd_sc_hd__mux2_1
X_20583_ _22503_/A VGND VGND VPWR VPWR _20583_/X sky130_fd_sc_hd__buf_6
X_32569_ _36025_/CLK _32569_/D VGND VGND VPWR VPWR _32569_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_393_CLK clkbuf_6_34__f_CLK/X VGND VGND VPWR VPWR _35758_/CLK sky130_fd_sc_hd__clkbuf_16
X_35357_ _35935_/CLK _35357_/D VGND VGND VPWR VPWR _35357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25110_ _25109_/X _33012_/Q _25113_/S VGND VGND VPWR VPWR _25111_/A sky130_fd_sc_hd__mux2_1
X_34308_ _34308_/CLK _34308_/D VGND VGND VPWR VPWR _34308_/Q sky130_fd_sc_hd__dfxtp_1
X_22322_ _33789_/Q _33725_/Q _33661_/Q _33597_/Q _22149_/X _22150_/X VGND VGND VPWR
+ VPWR _22322_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26090_ _25109_/X _33460_/Q _26092_/S VGND VGND VPWR VPWR _26091_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35288_ _35675_/CLK _35288_/D VGND VGND VPWR VPWR _35288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22253_ _34299_/Q _34235_/Q _34171_/Q _34107_/Q _22042_/X _22043_/X VGND VGND VPWR
+ VPWR _22253_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25041_ input8/X VGND VGND VPWR VPWR _25041_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_145_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _35277_/CLK sky130_fd_sc_hd__clkbuf_16
X_34239_ _36161_/CLK _34239_/D VGND VGND VPWR VPWR _34239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21204_ _32989_/Q _32925_/Q _32861_/Q _32797_/Q _20883_/X _20884_/X VGND VGND VPWR
+ VPWR _21204_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22184_ _22184_/A _22184_/B _22184_/C _22184_/D VGND VGND VPWR VPWR _22185_/A sky130_fd_sc_hd__or4_4
XFILLER_69_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21135_ _33243_/Q _36123_/Q _33115_/Q _33051_/Q _20952_/X _20953_/X VGND VGND VPWR
+ VPWR _21135_/X sky130_fd_sc_hd__mux4_1
X_28800_ _28911_/S VGND VGND VPWR VPWR _28819_/S sky130_fd_sc_hd__buf_4
X_29780_ _29780_/A VGND VGND VPWR VPWR _35145_/D sky130_fd_sc_hd__clkbuf_1
X_26992_ _26992_/A VGND VGND VPWR VPWR _33860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28731_ _26950_/X _34679_/Q _28747_/S VGND VGND VPWR VPWR _28732_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21066_ _32729_/Q _32665_/Q _32601_/Q _36057_/Q _20813_/X _20950_/X VGND VGND VPWR
+ VPWR _21066_/X sky130_fd_sc_hd__mux4_1
X_25943_ _25091_/X _33390_/Q _25957_/S VGND VGND VPWR VPWR _25944_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20017_ _35068_/Q _35004_/Q _34940_/Q _34876_/Q _19809_/X _19810_/X VGND VGND VPWR
+ VPWR _20017_/X sky130_fd_sc_hd__mux4_1
XFILLER_24_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28662_ _28662_/A VGND VGND VPWR VPWR _34646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25874_ _31410_/B _26685_/B VGND VGND VPWR VPWR _26007_/S sky130_fd_sc_hd__nand2_8
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1029 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27613_ _34149_/Q _24317_/X _27625_/S VGND VGND VPWR VPWR _27614_/A sky130_fd_sc_hd__mux2_1
X_24825_ _24852_/S VGND VGND VPWR VPWR _24844_/S sky130_fd_sc_hd__buf_6
XFILLER_228_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28593_ _28641_/S VGND VGND VPWR VPWR _28612_/S sky130_fd_sc_hd__clkbuf_8
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27544_ _27544_/A VGND VGND VPWR VPWR _34117_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24756_ _22932_/X _32863_/Q _24760_/S VGND VGND VPWR VPWR _24757_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21968_ _21968_/A VGND VGND VPWR VPWR _36210_/D sky130_fd_sc_hd__buf_6
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23707_ _22886_/X _32400_/Q _23721_/S VGND VGND VPWR VPWR _23708_/A sky130_fd_sc_hd__mux2_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20919_ _32725_/Q _32661_/Q _32597_/Q _36053_/Q _20813_/X _22313_/A VGND VGND VPWR
+ VPWR _20919_/X sky130_fd_sc_hd__mux4_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27475_ _27475_/A VGND VGND VPWR VPWR _34084_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_226_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24687_ _24687_/A VGND VGND VPWR VPWR _32831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21899_ _33777_/Q _33713_/Q _33649_/Q _33585_/Q _21796_/X _21797_/X VGND VGND VPWR
+ VPWR _21899_/X sky130_fd_sc_hd__mux4_1
X_29214_ _34882_/Q _29213_/X _29235_/S VGND VGND VPWR VPWR _29215_/A sky130_fd_sc_hd__mux2_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26426_ _25007_/X _33619_/Q _26434_/S VGND VGND VPWR VPWR _26427_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23638_ _32369_/Q _23253_/X _23646_/S VGND VGND VPWR VPWR _23639_/A sky130_fd_sc_hd__mux2_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29145_ _29247_/S VGND VGND VPWR VPWR _29173_/S sky130_fd_sc_hd__buf_4
XFILLER_70_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26357_ _26357_/A VGND VGND VPWR VPWR _33586_/D sky130_fd_sc_hd__clkbuf_1
X_23569_ _32336_/Q _23093_/X _23583_/S VGND VGND VPWR VPWR _23570_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_384_CLK clkbuf_6_41__f_CLK/X VGND VGND VPWR VPWR _35955_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_167_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16110_ _33999_/Q _33935_/Q _33871_/Q _32143_/Q _16108_/X _16109_/X VGND VGND VPWR
+ VPWR _16110_/X sky130_fd_sc_hd__mux4_1
XFILLER_183_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25308_ _25165_/X _33094_/Q _25314_/S VGND VGND VPWR VPWR _25309_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_947 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29076_ input63/X VGND VGND VPWR VPWR _29076_/X sky130_fd_sc_hd__clkbuf_4
X_17090_ _17957_/A VGND VGND VPWR VPWR _17090_/X sky130_fd_sc_hd__buf_4
X_26288_ _26288_/A VGND VGND VPWR VPWR _33553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16041_ input70/X VGND VGND VPWR VPWR _17843_/A sky130_fd_sc_hd__buf_12
X_28027_ _28027_/A VGND VGND VPWR VPWR _34345_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_136_CLK clkbuf_6_22__f_CLK/X VGND VGND VPWR VPWR _35597_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_183_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25239_ _25063_/X _33061_/Q _25251_/S VGND VGND VPWR VPWR _25240_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19800_ _20153_/A VGND VGND VPWR VPWR _19800_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_237_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17992_ _17705_/X _17990_/X _17991_/X _17708_/X VGND VGND VPWR VPWR _17992_/X sky130_fd_sc_hd__a22o_1
XFILLER_46_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29978_ _35239_/Q _29129_/X _29986_/S VGND VGND VPWR VPWR _29979_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16943_ _16939_/X _16942_/X _16808_/X VGND VGND VPWR VPWR _16944_/D sky130_fd_sc_hd__o21ba_1
X_19731_ _19725_/X _19730_/X _19447_/X VGND VGND VPWR VPWR _19739_/C sky130_fd_sc_hd__o21ba_1
XFILLER_172_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28929_ _34773_/Q _24267_/X _28933_/S VGND VGND VPWR VPWR _28930_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31940_ _23333_/X _36169_/Q _31940_/S VGND VGND VPWR VPWR _31941_/A sky130_fd_sc_hd__mux2_1
X_16874_ _34532_/Q _32420_/Q _34404_/Q _34340_/Q _16872_/X _16873_/X VGND VGND VPWR
+ VPWR _16874_/X sky130_fd_sc_hd__mux4_1
X_19662_ _19449_/X _19658_/X _19661_/X _19452_/X VGND VGND VPWR VPWR _19662_/X sky130_fd_sc_hd__a22o_1
XFILLER_37_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18613_ _33493_/Q _33429_/Q _33365_/Q _33301_/Q _18298_/X _18299_/X VGND VGND VPWR
+ VPWR _18613_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19593_ _34544_/Q _32432_/Q _34416_/Q _34352_/Q _19525_/X _19526_/X VGND VGND VPWR
+ VPWR _19593_/X sky130_fd_sc_hd__mux4_1
X_31871_ _23223_/X _36136_/Q _31877_/S VGND VGND VPWR VPWR _31872_/A sky130_fd_sc_hd__mux2_1
XTAP_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33610_ _35977_/CLK _33610_/D VGND VGND VPWR VPWR _33610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30822_ _30822_/A VGND VGND VPWR VPWR _35638_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18544_ _34003_/Q _33939_/Q _33875_/Q _32147_/Q _18408_/X _18409_/X VGND VGND VPWR
+ VPWR _18544_/X sky130_fd_sc_hd__mux4_1
XTAP_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34590_ _34781_/CLK _34590_/D VGND VGND VPWR VPWR _34590_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18475_ _34257_/Q _34193_/Q _34129_/Q _34065_/Q _18305_/X _18307_/X VGND VGND VPWR
+ VPWR _18475_/X sky130_fd_sc_hd__mux4_1
X_33541_ _33545_/CLK _33541_/D VGND VGND VPWR VPWR _33541_/Q sky130_fd_sc_hd__dfxtp_1
X_30753_ _23111_/X _35606_/Q _30755_/S VGND VGND VPWR VPWR _30754_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_370 _36208_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_381 _36208_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_392 _36209_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17426_ _35572_/Q _35508_/Q _35444_/Q _35380_/Q _17250_/X _17251_/X VGND VGND VPWR
+ VPWR _17426_/X sky130_fd_sc_hd__mux4_1
X_33472_ _34305_/CLK _33472_/D VGND VGND VPWR VPWR _33472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30684_ _30684_/A VGND VGND VPWR VPWR _35573_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35211_ _35338_/CLK _35211_/D VGND VGND VPWR VPWR _35211_/Q sky130_fd_sc_hd__dfxtp_1
X_32423_ _35302_/CLK _32423_/D VGND VGND VPWR VPWR _32423_/Q sky130_fd_sc_hd__dfxtp_1
X_17357_ _17351_/X _17356_/X _17147_/X VGND VGND VPWR VPWR _17367_/C sky130_fd_sc_hd__o21ba_1
X_36191_ _36191_/CLK _36191_/D VGND VGND VPWR VPWR _36191_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_375_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _36076_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_159_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16308_ _16308_/A _16308_/B _16308_/C _16308_/D VGND VGND VPWR VPWR _16309_/A sky130_fd_sc_hd__or4_4
XFILLER_105_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35142_ _35845_/CLK _35142_/D VGND VGND VPWR VPWR _35142_/Q sky130_fd_sc_hd__dfxtp_1
X_32354_ _36004_/CLK _32354_/D VGND VGND VPWR VPWR _32354_/Q sky130_fd_sc_hd__dfxtp_1
X_17288_ _17994_/A VGND VGND VPWR VPWR _17288_/X sky130_fd_sc_hd__buf_6
XFILLER_105_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19027_ _35296_/Q _35232_/Q _35168_/Q _32288_/Q _18953_/X _18954_/X VGND VGND VPWR
+ VPWR _19027_/X sky130_fd_sc_hd__mux4_1
X_31305_ _31305_/A VGND VGND VPWR VPWR _35867_/D sky130_fd_sc_hd__clkbuf_1
X_35073_ _35075_/CLK _35073_/D VGND VGND VPWR VPWR _35073_/Q sky130_fd_sc_hd__dfxtp_1
X_16239_ _16239_/A VGND VGND VPWR VPWR _31954_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_127_CLK clkbuf_6_23__f_CLK/X VGND VGND VPWR VPWR _34260_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_173_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32285_ _35293_/CLK _32285_/D VGND VGND VPWR VPWR _32285_/Q sky130_fd_sc_hd__dfxtp_1
X_34024_ _34153_/CLK _34024_/D VGND VGND VPWR VPWR _34024_/Q sky130_fd_sc_hd__dfxtp_1
X_31236_ _35835_/Q input40/X _31244_/S VGND VGND VPWR VPWR _31237_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31167_ _35802_/Q input4/X _31181_/S VGND VGND VPWR VPWR _31168_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30118_ _30118_/A VGND VGND VPWR VPWR _35305_/D sky130_fd_sc_hd__clkbuf_1
X_19929_ _20282_/A VGND VGND VPWR VPWR _19929_/X sky130_fd_sc_hd__buf_6
X_35975_ _35975_/CLK _35975_/D VGND VGND VPWR VPWR _35975_/Q sky130_fd_sc_hd__dfxtp_1
X_31098_ _31098_/A VGND VGND VPWR VPWR _35769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30049_ _35273_/Q _29234_/X _30049_/S VGND VGND VPWR VPWR _30050_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34926_ _35054_/CLK _34926_/D VGND VGND VPWR VPWR _34926_/Q sky130_fd_sc_hd__dfxtp_1
X_22940_ _22940_/A VGND VGND VPWR VPWR _32033_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22871_ _20656_/X _22869_/X _22870_/X _20668_/X VGND VGND VPWR VPWR _22871_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34857_ _35943_/CLK _34857_/D VGND VGND VPWR VPWR _34857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24610_ _24610_/A VGND VGND VPWR VPWR _32794_/D sky130_fd_sc_hd__clkbuf_1
X_33808_ _35728_/CLK _33808_/D VGND VGND VPWR VPWR _33808_/Q sky130_fd_sc_hd__dfxtp_1
X_21822_ _34798_/Q _34734_/Q _34670_/Q _34606_/Q _21535_/X _21536_/X VGND VGND VPWR
+ VPWR _21822_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25590_ _25590_/A VGND VGND VPWR VPWR _33225_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34788_ _36003_/CLK _34788_/D VGND VGND VPWR VPWR _34788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24541_ _24541_/A VGND VGND VPWR VPWR _32763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33739_ _35977_/CLK _33739_/D VGND VGND VPWR VPWR _33739_/Q sky130_fd_sc_hd__dfxtp_1
X_21753_ _21749_/X _21750_/X _21751_/X _21752_/X VGND VGND VPWR VPWR _21753_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20704_ _33743_/Q _33679_/Q _33615_/Q _33551_/Q _20580_/X _20583_/X VGND VGND VPWR
+ VPWR _20704_/X sky130_fd_sc_hd__mux4_1
X_27260_ _26974_/X _33983_/Q _27260_/S VGND VGND VPWR VPWR _27261_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24472_ _24472_/A VGND VGND VPWR VPWR _32730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21684_ _21401_/X _21682_/X _21683_/X _21406_/X VGND VGND VPWR VPWR _21684_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26211_ _25088_/X _33517_/Q _26227_/S VGND VGND VPWR VPWR _26212_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23423_ _30329_/A _29049_/B _30329_/B VGND VGND VPWR VPWR _29384_/A sky130_fd_sc_hd__nor3b_4
X_35409_ _35922_/CLK _35409_/D VGND VGND VPWR VPWR _35409_/Q sky130_fd_sc_hd__dfxtp_1
X_20635_ _22430_/A VGND VGND VPWR VPWR _20635_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_366_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _36147_/CLK sky130_fd_sc_hd__clkbuf_16
X_27191_ _26872_/X _33950_/Q _27197_/S VGND VGND VPWR VPWR _27192_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26142_ _25186_/X _33485_/Q _26142_/S VGND VGND VPWR VPWR _26143_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20566_ _34829_/Q _34765_/Q _34701_/Q _34637_/Q _20294_/X _20295_/X VGND VGND VPWR
+ VPWR _20566_/X sky130_fd_sc_hd__mux4_1
X_23354_ _23354_/A VGND VGND VPWR VPWR _32236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22305_ _22460_/A VGND VGND VPWR VPWR _22305_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_118_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _34006_/CLK sky130_fd_sc_hd__clkbuf_16
X_26073_ _26142_/S VGND VGND VPWR VPWR _26092_/S sky130_fd_sc_hd__buf_4
X_20497_ _19454_/A _20495_/X _20496_/X _19459_/A VGND VGND VPWR VPWR _20497_/X sky130_fd_sc_hd__a22o_1
X_23285_ _23285_/A VGND VGND VPWR VPWR _32212_/D sky130_fd_sc_hd__clkbuf_1
X_29901_ _29901_/A VGND VGND VPWR VPWR _35202_/D sky130_fd_sc_hd__clkbuf_1
X_25024_ _25022_/X _32984_/Q _25051_/S VGND VGND VPWR VPWR _25025_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22236_ _21947_/X _22234_/X _22235_/X _21950_/X VGND VGND VPWR VPWR _22236_/X sky130_fd_sc_hd__a22o_1
XFILLER_195_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22167_ _22163_/X _22166_/X _22089_/X _22090_/X VGND VGND VPWR VPWR _22184_/B sky130_fd_sc_hd__o211a_1
X_29832_ _29922_/S VGND VGND VPWR VPWR _29851_/S sky130_fd_sc_hd__buf_4
XTAP_6924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21118_ _21043_/X _21116_/X _21117_/X _21046_/X VGND VGND VPWR VPWR _21118_/X sky130_fd_sc_hd__a22o_1
XTAP_6957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29763_ _35137_/Q _29210_/X _29779_/S VGND VGND VPWR VPWR _29764_/A sky130_fd_sc_hd__mux2_1
X_26975_ _26974_/X _33855_/Q _26975_/S VGND VGND VPWR VPWR _26976_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22098_ _33206_/Q _32566_/Q _35958_/Q _35894_/Q _22027_/X _22028_/X VGND VGND VPWR
+ VPWR _22098_/X sky130_fd_sc_hd__mux4_1
XTAP_6979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25926_ _25066_/X _33382_/Q _25936_/S VGND VGND VPWR VPWR _25927_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28714_ _26925_/X _34671_/Q _28726_/S VGND VGND VPWR VPWR _28715_/A sky130_fd_sc_hd__mux2_1
X_21049_ _34520_/Q _32408_/Q _34392_/Q _34328_/Q _20766_/X _20767_/X VGND VGND VPWR
+ VPWR _21049_/X sky130_fd_sc_hd__mux4_1
X_29694_ _29694_/A VGND VGND VPWR VPWR _35104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1041 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28645_ _26821_/X _34638_/Q _28663_/S VGND VGND VPWR VPWR _28646_/A sky130_fd_sc_hd__mux2_1
X_25857_ _25857_/A VGND VGND VPWR VPWR _33349_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24808_ _24808_/A VGND VGND VPWR VPWR _32887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28576_ _28576_/A VGND VGND VPWR VPWR _34605_/D sky130_fd_sc_hd__clkbuf_1
X_16590_ _16586_/X _16589_/X _16455_/X VGND VGND VPWR VPWR _16591_/D sky130_fd_sc_hd__o21ba_1
XFILLER_90_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25788_ _25788_/A VGND VGND VPWR VPWR _33316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27527_ _27527_/A VGND VGND VPWR VPWR _34109_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24739_ _22907_/X _32855_/Q _24739_/S VGND VGND VPWR VPWR _24740_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _35789_/Q _35149_/Q _34509_/Q _33869_/Q _16108_/X _16109_/X VGND VGND VPWR
+ VPWR _18260_/X sky130_fd_sc_hd__mux4_1
XFILLER_202_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27458_ _27458_/A VGND VGND VPWR VPWR _34076_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _32494_/Q _32366_/Q _32046_/Q _36014_/Q _16923_/X _17064_/X VGND VGND VPWR
+ VPWR _17211_/X sky130_fd_sc_hd__mux4_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26409_ _26409_/A VGND VGND VPWR VPWR _33611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18191_ _18187_/X _18190_/X _17834_/A VGND VGND VPWR VPWR _18213_/A sky130_fd_sc_hd__o21ba_1
XFILLER_204_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27389_ _34044_/Q _24388_/X _27395_/S VGND VGND VPWR VPWR _27390_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_1406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_357_CLK clkbuf_6_41__f_CLK/X VGND VGND VPWR VPWR _36019_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17142_ _35756_/Q _35116_/Q _34476_/Q _33836_/Q _17140_/X _17141_/X VGND VGND VPWR
+ VPWR _17142_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29128_ _29128_/A VGND VGND VPWR VPWR _34854_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_109_CLK clkbuf_6_22__f_CLK/X VGND VGND VPWR VPWR _35279_/CLK sky130_fd_sc_hd__clkbuf_16
X_29059_ _34832_/Q _29058_/X _29080_/S VGND VGND VPWR VPWR _29060_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17073_ _35562_/Q _35498_/Q _35434_/Q _35370_/Q _16897_/X _16898_/X VGND VGND VPWR
+ VPWR _17073_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16024_ _16014_/X _16019_/X _16022_/X _16023_/X VGND VGND VPWR VPWR _16024_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32070_ _32518_/CLK _32070_/D VGND VGND VPWR VPWR _32070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31021_ _35733_/Q _29073_/X _31025_/S VGND VGND VPWR VPWR _31022_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17975_ _34052_/Q _33988_/Q _33924_/Q _32260_/Q _17726_/X _17727_/X VGND VGND VPWR
+ VPWR _17975_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19714_ _20206_/A VGND VGND VPWR VPWR _19714_/X sky130_fd_sc_hd__clkbuf_4
X_35760_ _35760_/CLK _35760_/D VGND VGND VPWR VPWR _35760_/Q sky130_fd_sc_hd__dfxtp_1
X_16926_ _16710_/X _16924_/X _16925_/X _16714_/X VGND VGND VPWR VPWR _16926_/X sky130_fd_sc_hd__a22o_1
XFILLER_215_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32972_ _35917_/CLK _32972_/D VGND VGND VPWR VPWR _32972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34711_ _36202_/CLK _34711_/D VGND VGND VPWR VPWR _34711_/Q sky130_fd_sc_hd__dfxtp_1
X_31923_ _31923_/A VGND VGND VPWR VPWR _36160_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19645_ _19363_/X _19641_/X _19644_/X _19367_/X VGND VGND VPWR VPWR _19645_/X sky130_fd_sc_hd__a22o_1
X_35691_ _35818_/CLK _35691_/D VGND VGND VPWR VPWR _35691_/Q sky130_fd_sc_hd__dfxtp_1
X_16857_ _16702_/X _16855_/X _16856_/X _16708_/X VGND VGND VPWR VPWR _16857_/X sky130_fd_sc_hd__a22o_1
XFILLER_226_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_915 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34642_ _34775_/CLK _34642_/D VGND VGND VPWR VPWR _34642_/Q sky130_fd_sc_hd__dfxtp_1
X_16788_ _17995_/A VGND VGND VPWR VPWR _16788_/X sky130_fd_sc_hd__buf_4
X_31854_ _23142_/X _36128_/Q _31856_/S VGND VGND VPWR VPWR _31855_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19576_ _20282_/A VGND VGND VPWR VPWR _19576_/X sky130_fd_sc_hd__buf_6
XFILLER_244_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18527_ _18356_/X _18525_/X _18526_/X _18368_/X VGND VGND VPWR VPWR _18527_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30805_ _30805_/A VGND VGND VPWR VPWR _35630_/D sky130_fd_sc_hd__clkbuf_1
X_34573_ _35981_/CLK _34573_/D VGND VGND VPWR VPWR _34573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31785_ _31785_/A VGND VGND VPWR VPWR _36095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33524_ _33779_/CLK _33524_/D VGND VGND VPWR VPWR _33524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18458_ _18344_/X _18456_/X _18457_/X _18354_/X VGND VGND VPWR VPWR _18458_/X sky130_fd_sc_hd__a22o_1
X_30736_ _30868_/S VGND VGND VPWR VPWR _30755_/S sky130_fd_sc_hd__buf_4
XFILLER_107_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17409_ _17762_/A VGND VGND VPWR VPWR _17409_/X sky130_fd_sc_hd__clkbuf_4
X_18389_ _20062_/A VGND VGND VPWR VPWR _19173_/A sky130_fd_sc_hd__buf_12
XFILLER_21_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30667_ _35565_/Q _29148_/X _30683_/S VGND VGND VPWR VPWR _30668_/A sky130_fd_sc_hd__mux2_1
X_33455_ _33520_/CLK _33455_/D VGND VGND VPWR VPWR _33455_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_348_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _34289_/CLK sky130_fd_sc_hd__clkbuf_16
X_20420_ _35080_/Q _35016_/Q _34952_/Q _34888_/Q _20162_/X _20163_/X VGND VGND VPWR
+ VPWR _20420_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32406_ _35669_/CLK _32406_/D VGND VGND VPWR VPWR _32406_/Q sky130_fd_sc_hd__dfxtp_1
X_36174_ _36185_/CLK _36174_/D VGND VGND VPWR VPWR _36174_/Q sky130_fd_sc_hd__dfxtp_1
X_30598_ _23345_/X _35533_/Q _30598_/S VGND VGND VPWR VPWR _30599_/A sky130_fd_sc_hd__mux2_1
X_33386_ _33512_/CLK _33386_/D VGND VGND VPWR VPWR _33386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20351_ _18277_/X _20349_/X _20350_/X _18287_/X VGND VGND VPWR VPWR _20351_/X sky130_fd_sc_hd__a22o_1
XFILLER_140_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35125_ _35829_/CLK _35125_/D VGND VGND VPWR VPWR _35125_/Q sky130_fd_sc_hd__dfxtp_1
X_32337_ _36049_/CLK _32337_/D VGND VGND VPWR VPWR _32337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23070_ _23070_/A VGND VGND VPWR VPWR _32075_/D sky130_fd_sc_hd__clkbuf_1
X_32268_ _34316_/CLK _32268_/D VGND VGND VPWR VPWR _32268_/Q sky130_fd_sc_hd__dfxtp_1
X_20282_ _20282_/A VGND VGND VPWR VPWR _20282_/X sky130_fd_sc_hd__buf_6
X_35056_ _35760_/CLK _35056_/D VGND VGND VPWR VPWR _35056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22021_ _22016_/X _22018_/X _22019_/X _22020_/X VGND VGND VPWR VPWR _22021_/X sky130_fd_sc_hd__a22o_1
XTAP_6209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34007_ _35280_/CLK _34007_/D VGND VGND VPWR VPWR _34007_/Q sky130_fd_sc_hd__dfxtp_1
X_31219_ _35827_/Q input31/X _31223_/S VGND VGND VPWR VPWR _31220_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32199_ _35822_/CLK _32199_/D VGND VGND VPWR VPWR _32199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26760_ _26760_/A VGND VGND VPWR VPWR _33776_/D sky130_fd_sc_hd__clkbuf_1
X_23972_ _30329_/A _30329_/B _29049_/B VGND VGND VPWR VPWR _31410_/A sky130_fd_sc_hd__nor3_4
XTAP_4829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35958_ _35958_/CLK _35958_/D VGND VGND VPWR VPWR _35958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25711_ _33281_/Q _24404_/X _25727_/S VGND VGND VPWR VPWR _25712_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34909_ _35036_/CLK _34909_/D VGND VGND VPWR VPWR _34909_/Q sky130_fd_sc_hd__dfxtp_1
X_22923_ input6/X VGND VGND VPWR VPWR _22923_/X sky130_fd_sc_hd__buf_4
X_26691_ _26691_/A VGND VGND VPWR VPWR _33743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1029 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35889_ _35889_/CLK _35889_/D VGND VGND VPWR VPWR _35889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28430_ _28430_/A VGND VGND VPWR VPWR _34536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25642_ _25642_/A VGND VGND VPWR VPWR _33248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22854_ _21749_/A _22852_/X _22853_/X _21752_/A VGND VGND VPWR VPWR _22854_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28361_ _34504_/Q _24425_/X _28363_/S VGND VGND VPWR VPWR _28362_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21805_ _22511_/A VGND VGND VPWR VPWR _21805_/X sky130_fd_sc_hd__clkbuf_4
X_25573_ _33217_/Q _24404_/X _25589_/S VGND VGND VPWR VPWR _25574_/A sky130_fd_sc_hd__mux2_1
XFILLER_227_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22785_ _33803_/Q _33739_/Q _33675_/Q _33611_/Q _22502_/X _22503_/X VGND VGND VPWR
+ VPWR _22785_/X sky130_fd_sc_hd__mux4_1
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27312_ _27312_/A VGND VGND VPWR VPWR _34007_/D sky130_fd_sc_hd__clkbuf_1
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24524_ _24524_/A VGND VGND VPWR VPWR _32755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28292_ _34471_/Q _24323_/X _28300_/S VGND VGND VPWR VPWR _28293_/A sky130_fd_sc_hd__mux2_1
X_21736_ _22442_/A VGND VGND VPWR VPWR _21736_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_197_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27243_ _27243_/A VGND VGND VPWR VPWR _33974_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24455_ _24455_/A VGND VGND VPWR VPWR _32722_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_339_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _34296_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21667_ _22511_/A VGND VGND VPWR VPWR _21667_/X sky130_fd_sc_hd__buf_4
XFILLER_61_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23406_ _23406_/A VGND VGND VPWR VPWR _32261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27174_ _26847_/X _33942_/Q _27176_/S VGND VGND VPWR VPWR _27175_/A sky130_fd_sc_hd__mux2_1
X_20618_ _22362_/A VGND VGND VPWR VPWR _22313_/A sky130_fd_sc_hd__buf_4
XFILLER_240_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24386_ _32699_/Q _24385_/X _24398_/S VGND VGND VPWR VPWR _24387_/A sky130_fd_sc_hd__mux2_1
X_21598_ _21594_/X _21595_/X _21596_/X _21597_/X VGND VGND VPWR VPWR _21598_/X sky130_fd_sc_hd__a22o_1
X_26125_ _26125_/A VGND VGND VPWR VPWR _33476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23337_ _32230_/Q _23336_/X _23346_/S VGND VGND VPWR VPWR _23338_/A sky130_fd_sc_hd__mux2_1
X_20549_ _34061_/Q _33997_/Q _33933_/Q _32269_/Q _18358_/X _18360_/X VGND VGND VPWR
+ VPWR _20549_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26056_ _26056_/A VGND VGND VPWR VPWR _33443_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23268_ _32207_/Q _23267_/X _23268_/S VGND VGND VPWR VPWR _23269_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25007_ input56/X VGND VGND VPWR VPWR _25007_/X sky130_fd_sc_hd__buf_4
XFILLER_69_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22219_ _34298_/Q _34234_/Q _34170_/Q _34106_/Q _22042_/X _22043_/X VGND VGND VPWR
+ VPWR _22219_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23199_ input16/X VGND VGND VPWR VPWR _23199_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29815_ _29815_/A VGND VGND VPWR VPWR _35161_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17760_ _17756_/X _17759_/X _17481_/X VGND VGND VPWR VPWR _17792_/A sky130_fd_sc_hd__o21ba_1
X_29746_ _35129_/Q _29185_/X _29758_/S VGND VGND VPWR VPWR _29747_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26958_ _26958_/A VGND VGND VPWR VPWR _33849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16711_ _17770_/A VGND VGND VPWR VPWR _16711_/X sky130_fd_sc_hd__clkbuf_4
X_17691_ _32764_/Q _32700_/Q _32636_/Q _36092_/Q _17625_/X _17409_/X VGND VGND VPWR
+ VPWR _17691_/X sky130_fd_sc_hd__mux4_1
X_25909_ _25041_/X _33374_/Q _25915_/S VGND VGND VPWR VPWR _25910_/A sky130_fd_sc_hd__mux2_1
X_26889_ _26888_/X _33827_/Q _26913_/S VGND VGND VPWR VPWR _26890_/A sky130_fd_sc_hd__mux2_1
X_29677_ _35096_/Q _29082_/X _29695_/S VGND VGND VPWR VPWR _29678_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19430_ _32748_/Q _32684_/Q _32620_/Q _36076_/Q _19219_/X _19356_/X VGND VGND VPWR
+ VPWR _19430_/X sky130_fd_sc_hd__mux4_1
X_16642_ _35806_/Q _32181_/Q _35678_/Q _35614_/Q _16607_/X _16608_/X VGND VGND VPWR
+ VPWR _16642_/X sky130_fd_sc_hd__mux4_1
X_28628_ _28628_/A VGND VGND VPWR VPWR _34630_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19361_ _20206_/A VGND VGND VPWR VPWR _19361_/X sky130_fd_sc_hd__clkbuf_8
X_16573_ _16357_/X _16571_/X _16572_/X _16361_/X VGND VGND VPWR VPWR _16573_/X sky130_fd_sc_hd__a22o_1
X_28559_ _28559_/A VGND VGND VPWR VPWR _34597_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18312_ _18293_/X _18309_/X _18311_/X VGND VGND VPWR VPWR _18402_/A sky130_fd_sc_hd__o21ba_1
XFILLER_231_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31570_ _35993_/Q input3/X _31586_/S VGND VGND VPWR VPWR _31571_/A sky130_fd_sc_hd__mux2_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19292_ _19010_/X _19288_/X _19291_/X _19014_/X VGND VGND VPWR VPWR _19292_/X sky130_fd_sc_hd__a22o_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _18243_/A _18243_/B _18243_/C _18243_/D VGND VGND VPWR VPWR _18244_/A sky130_fd_sc_hd__or4_4
XFILLER_128_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30521_ _23223_/X _35496_/Q _30527_/S VGND VGND VPWR VPWR _30522_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18174_ _15997_/X _18172_/X _18173_/X _16003_/X VGND VGND VPWR VPWR _18174_/X sky130_fd_sc_hd__a22o_1
X_30452_ _30452_/A VGND VGND VPWR VPWR _35463_/D sky130_fd_sc_hd__clkbuf_1
X_33240_ _36121_/CLK _33240_/D VGND VGND VPWR VPWR _33240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17125_ _33516_/Q _33452_/Q _33388_/Q _33324_/Q _17123_/X _17124_/X VGND VGND VPWR
+ VPWR _17125_/X sky130_fd_sc_hd__mux4_2
X_33171_ _36114_/CLK _33171_/D VGND VGND VPWR VPWR _33171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30383_ _30383_/A VGND VGND VPWR VPWR _35430_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32122_ _35562_/CLK _32122_/D VGND VGND VPWR VPWR _32122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17056_ _17762_/A VGND VGND VPWR VPWR _17056_/X sky130_fd_sc_hd__buf_6
XFILLER_239_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16007_ _17957_/A VGND VGND VPWR VPWR _16007_/X sky130_fd_sc_hd__buf_4
X_32053_ _36021_/CLK _32053_/D VGND VGND VPWR VPWR _32053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31004_ _31004_/A VGND VGND VPWR VPWR _35725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35812_ _35814_/CLK _35812_/D VGND VGND VPWR VPWR _35812_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _35587_/Q _35523_/Q _35459_/Q _35395_/Q _17956_/X _17957_/X VGND VGND VPWR
+ VPWR _17958_/X sky130_fd_sc_hd__mux4_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35743_ _35743_/CLK _35743_/D VGND VGND VPWR VPWR _35743_/Q sky130_fd_sc_hd__dfxtp_1
X_16909_ _16905_/X _16908_/X _16808_/X VGND VGND VPWR VPWR _16910_/D sky130_fd_sc_hd__o21ba_1
X_32955_ _36090_/CLK _32955_/D VGND VGND VPWR VPWR _32955_/Q sky130_fd_sc_hd__dfxtp_1
X_17889_ _33217_/Q _32577_/Q _35969_/Q _35905_/Q _17780_/X _17781_/X VGND VGND VPWR
+ VPWR _17889_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31906_ _31906_/A VGND VGND VPWR VPWR _36152_/D sky130_fd_sc_hd__clkbuf_1
X_19628_ _19624_/X _19627_/X _19461_/X VGND VGND VPWR VPWR _19629_/D sky130_fd_sc_hd__o21ba_1
XFILLER_53_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35674_ _35675_/CLK _35674_/D VGND VGND VPWR VPWR _35674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32886_ _36022_/CLK _32886_/D VGND VGND VPWR VPWR _32886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34625_ _35330_/CLK _34625_/D VGND VGND VPWR VPWR _34625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31837_ _31948_/S VGND VGND VPWR VPWR _31856_/S sky130_fd_sc_hd__buf_4
X_19559_ _34543_/Q _32431_/Q _34415_/Q _34351_/Q _19525_/X _19526_/X VGND VGND VPWR
+ VPWR _19559_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22570_ _22570_/A VGND VGND VPWR VPWR _36227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34556_ _34620_/CLK _34556_/D VGND VGND VPWR VPWR _34556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31768_ _36087_/Q input36/X _31784_/S VGND VGND VPWR VPWR _31769_/A sky130_fd_sc_hd__mux2_1
X_33507_ _33507_/CLK _33507_/D VGND VGND VPWR VPWR _33507_/Q sky130_fd_sc_hd__dfxtp_1
X_21521_ _33254_/Q _36134_/Q _33126_/Q _33062_/Q _21305_/X _21306_/X VGND VGND VPWR
+ VPWR _21521_/X sky130_fd_sc_hd__mux4_1
X_30719_ _35590_/Q _29225_/X _30725_/S VGND VGND VPWR VPWR _30720_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34487_ _35831_/CLK _34487_/D VGND VGND VPWR VPWR _34487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31699_ _31699_/A VGND VGND VPWR VPWR _36054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36226_ _36228_/CLK _36226_/D VGND VGND VPWR VPWR _36226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24240_ _23071_/X _32652_/Q _24242_/S VGND VGND VPWR VPWR _24241_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21452_ _22511_/A VGND VGND VPWR VPWR _21452_/X sky130_fd_sc_hd__clkbuf_4
X_33438_ _33946_/CLK _33438_/D VGND VGND VPWR VPWR _33438_/Q sky130_fd_sc_hd__dfxtp_1
X_20403_ _33288_/Q _36168_/Q _33160_/Q _33096_/Q _18328_/X _19457_/A VGND VGND VPWR
+ VPWR _20403_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_928 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36157_ _36157_/CLK _36157_/D VGND VGND VPWR VPWR _36157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24171_ _22969_/X _32619_/Q _24171_/S VGND VGND VPWR VPWR _24172_/A sky130_fd_sc_hd__mux2_1
X_21383_ _22442_/A VGND VGND VPWR VPWR _21383_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_147_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33369_ _35284_/CLK _33369_/D VGND VGND VPWR VPWR _33369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23122_ _32153_/Q _23121_/X _23146_/S VGND VGND VPWR VPWR _23123_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35108_ _35748_/CLK _35108_/D VGND VGND VPWR VPWR _35108_/Q sky130_fd_sc_hd__dfxtp_1
X_20334_ _20334_/A VGND VGND VPWR VPWR _32133_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_123_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36088_ _36088_/CLK _36088_/D VGND VGND VPWR VPWR _36088_/Q sky130_fd_sc_hd__dfxtp_1
X_20265_ _34563_/Q _32451_/Q _34435_/Q _34371_/Q _20231_/X _20232_/X VGND VGND VPWR
+ VPWR _20265_/X sky130_fd_sc_hd__mux4_1
X_23053_ input52/X VGND VGND VPWR VPWR _23053_/X sky130_fd_sc_hd__buf_4
X_27930_ _27930_/A VGND VGND VPWR VPWR _34299_/D sky130_fd_sc_hd__clkbuf_1
X_35039_ _35039_/CLK _35039_/D VGND VGND VPWR VPWR _35039_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22004_ _33524_/Q _33460_/Q _33396_/Q _33332_/Q _21723_/X _21724_/X VGND VGND VPWR
+ VPWR _22004_/X sky130_fd_sc_hd__mux4_1
XTAP_6039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27861_ _27861_/A VGND VGND VPWR VPWR _34266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20196_ _35073_/Q _35009_/Q _34945_/Q _34881_/Q _20162_/X _20163_/X VGND VGND VPWR
+ VPWR _20196_/X sky130_fd_sc_hd__mux4_1
XTAP_5305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29600_ _35060_/Q _29169_/X _29602_/S VGND VGND VPWR VPWR _29601_/A sky130_fd_sc_hd__mux2_1
X_26812_ _26812_/A VGND VGND VPWR VPWR _33801_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27792_ _34234_/Q _24382_/X _27802_/S VGND VGND VPWR VPWR _27793_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29531_ _35027_/Q _29067_/X _29539_/S VGND VGND VPWR VPWR _29532_/A sky130_fd_sc_hd__mux2_1
XTAP_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26743_ _26743_/A VGND VGND VPWR VPWR _33768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23955_ _23955_/A VGND VGND VPWR VPWR _32517_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22906_ _22906_/A VGND VGND VPWR VPWR _32022_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29462_ _29462_/A VGND VGND VPWR VPWR _34994_/D sky130_fd_sc_hd__clkbuf_1
X_26674_ _26674_/A VGND VGND VPWR VPWR _33736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_903 _26277_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23886_ _23886_/A VGND VGND VPWR VPWR _32484_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_914 _26956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_925 _27509_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_936 _29067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25625_ _33240_/Q _24276_/X _25643_/S VGND VGND VPWR VPWR _25626_/A sky130_fd_sc_hd__mux2_1
X_28413_ _28413_/A VGND VGND VPWR VPWR _34528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22837_ _35340_/Q _35276_/Q _35212_/Q _32332_/Q _20688_/X _20690_/X VGND VGND VPWR
+ VPWR _22837_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29393_ _29393_/A VGND VGND VPWR VPWR _34961_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_947 _29517_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_958 _29922_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_969 _31273_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28344_ _28371_/S VGND VGND VPWR VPWR _28363_/S sky130_fd_sc_hd__buf_4
XFILLER_169_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25556_ _33209_/Q _24379_/X _25568_/S VGND VGND VPWR VPWR _25557_/A sky130_fd_sc_hd__mux2_1
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22768_ _22764_/X _22767_/X _22442_/A _22443_/A VGND VGND VPWR VPWR _22783_/B sky130_fd_sc_hd__o211a_1
XFILLER_38_1356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24507_ _24507_/A VGND VGND VPWR VPWR _32747_/D sky130_fd_sc_hd__clkbuf_1
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21719_ _21719_/A VGND VGND VPWR VPWR _36203_/D sky130_fd_sc_hd__clkbuf_1
X_28275_ _34463_/Q _24298_/X _28279_/S VGND VGND VPWR VPWR _28276_/A sky130_fd_sc_hd__mux2_1
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25487_ _33176_/Q _24276_/X _25505_/S VGND VGND VPWR VPWR _25488_/A sky130_fd_sc_hd__mux2_1
X_22699_ _34056_/Q _33992_/Q _33928_/Q _32264_/Q _20658_/X _20660_/X VGND VGND VPWR
+ VPWR _22699_/X sky130_fd_sc_hd__mux4_1
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27226_ _27226_/A VGND VGND VPWR VPWR _33966_/D sky130_fd_sc_hd__clkbuf_1
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24438_ _32716_/Q _24437_/X _24441_/S VGND VGND VPWR VPWR _24439_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27157_ _27289_/S VGND VGND VPWR VPWR _27176_/S sky130_fd_sc_hd__buf_4
X_24369_ input35/X VGND VGND VPWR VPWR _24369_/X sky130_fd_sc_hd__buf_4
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26108_ _26108_/A VGND VGND VPWR VPWR _33468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27088_ _26919_/X _33901_/Q _27104_/S VGND VGND VPWR VPWR _27089_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26039_ _26039_/A VGND VGND VPWR VPWR _33435_/D sky130_fd_sc_hd__clkbuf_1
X_18930_ _18796_/X _18928_/X _18929_/X _18799_/X VGND VGND VPWR VPWR _18930_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_40_CLK clkbuf_6_7__f_CLK/X VGND VGND VPWR VPWR _33244_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_1302 _16525_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1313 input11/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18861_ _18789_/X _18859_/X _18860_/X _18794_/X VGND VGND VPWR VPWR _18861_/X sky130_fd_sc_hd__a22o_1
XTAP_6540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1324 _18124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1335 _19452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1346 _22443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17812_ _17700_/X _17810_/X _17811_/X _17703_/X VGND VGND VPWR VPWR _17812_/X sky130_fd_sc_hd__a22o_1
XANTENNA_1357 _22892_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1368 _24394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18792_ _33754_/Q _33690_/Q _33626_/Q _33562_/Q _18790_/X _18791_/X VGND VGND VPWR
+ VPWR _18792_/X sky130_fd_sc_hd__mux4_1
XTAP_6595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1379 _26928_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17743_ _17705_/X _17741_/X _17742_/X _17708_/X VGND VGND VPWR VPWR _17743_/X sky130_fd_sc_hd__a22o_1
X_29729_ _35121_/Q _29160_/X _29737_/S VGND VGND VPWR VPWR _29730_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32740_ _36069_/CLK _32740_/D VGND VGND VPWR VPWR _32740_/Q sky130_fd_sc_hd__dfxtp_1
X_17674_ _17670_/X _17673_/X _17500_/X VGND VGND VPWR VPWR _17682_/C sky130_fd_sc_hd__o21ba_1
XFILLER_36_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19413_ _19096_/X _19411_/X _19412_/X _19099_/X VGND VGND VPWR VPWR _19413_/X sky130_fd_sc_hd__a22o_1
XFILLER_35_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16625_ _33758_/Q _33694_/Q _33630_/Q _33566_/Q _16490_/X _16491_/X VGND VGND VPWR
+ VPWR _16625_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32671_ _34271_/CLK _32671_/D VGND VGND VPWR VPWR _32671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_929 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34410_ _35050_/CLK _34410_/D VGND VGND VPWR VPWR _34410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19344_ _19101_/X _19342_/X _19343_/X _19106_/X VGND VGND VPWR VPWR _19344_/X sky130_fd_sc_hd__a22o_1
X_31622_ _36018_/Q input30/X _31628_/S VGND VGND VPWR VPWR _31623_/A sky130_fd_sc_hd__mux2_1
X_16556_ _16552_/X _16555_/X _16455_/X VGND VGND VPWR VPWR _16557_/D sky130_fd_sc_hd__o21ba_1
X_35390_ _35966_/CLK _35390_/D VGND VGND VPWR VPWR _35390_/Q sky130_fd_sc_hd__dfxtp_1
X_34341_ _35941_/CLK _34341_/D VGND VGND VPWR VPWR _34341_/Q sky130_fd_sc_hd__dfxtp_1
X_31553_ _35985_/Q input34/X _31565_/S VGND VGND VPWR VPWR _31554_/A sky130_fd_sc_hd__mux2_1
X_19275_ _19271_/X _19274_/X _19108_/X VGND VGND VPWR VPWR _19276_/D sky130_fd_sc_hd__o21ba_1
X_16487_ _16487_/A _16487_/B _16487_/C _16487_/D VGND VGND VPWR VPWR _16488_/A sky130_fd_sc_hd__or4_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18226_ _33036_/Q _32972_/Q _32908_/Q _32844_/Q _15980_/X _15983_/X VGND VGND VPWR
+ VPWR _18226_/X sky130_fd_sc_hd__mux4_1
X_30504_ _23142_/X _35488_/Q _30506_/S VGND VGND VPWR VPWR _30505_/A sky130_fd_sc_hd__mux2_1
X_31484_ _31484_/A VGND VGND VPWR VPWR _35952_/D sky130_fd_sc_hd__clkbuf_1
X_34272_ _35675_/CLK _34272_/D VGND VGND VPWR VPWR _34272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36011_ _36011_/CLK _36011_/D VGND VGND VPWR VPWR _36011_/Q sky130_fd_sc_hd__dfxtp_1
X_33223_ _36168_/CLK _33223_/D VGND VGND VPWR VPWR _33223_/Q sky130_fd_sc_hd__dfxtp_1
X_30435_ _30435_/A VGND VGND VPWR VPWR _35455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18157_ _17901_/X _18155_/X _18156_/X _17906_/X VGND VGND VPWR VPWR _18157_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17108_ _33195_/Q _32555_/Q _35947_/Q _35883_/Q _17074_/X _17075_/X VGND VGND VPWR
+ VPWR _17108_/X sky130_fd_sc_hd__mux4_1
X_18088_ _17855_/X _18086_/X _18087_/X _17858_/X VGND VGND VPWR VPWR _18088_/X sky130_fd_sc_hd__a22o_1
X_33154_ _36159_/CLK _33154_/D VGND VGND VPWR VPWR _33154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30366_ _30366_/A VGND VGND VPWR VPWR _35422_/D sky130_fd_sc_hd__clkbuf_1
X_32105_ _35808_/CLK _32105_/D VGND VGND VPWR VPWR _32105_/Q sky130_fd_sc_hd__dfxtp_1
X_17039_ _34793_/Q _34729_/Q _34665_/Q _34601_/Q _16935_/X _16936_/X VGND VGND VPWR
+ VPWR _17039_/X sky130_fd_sc_hd__mux4_1
XFILLER_171_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33085_ _36095_/CLK _33085_/D VGND VGND VPWR VPWR _33085_/Q sky130_fd_sc_hd__dfxtp_1
X_30297_ _30297_/A VGND VGND VPWR VPWR _35390_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_31_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _34267_/CLK sky130_fd_sc_hd__clkbuf_16
X_20050_ _19807_/X _20048_/X _20049_/X _19812_/X VGND VGND VPWR VPWR _20050_/X sky130_fd_sc_hd__a22o_1
X_32036_ _36004_/CLK _32036_/D VGND VGND VPWR VPWR _32036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33987_ _34057_/CLK _33987_/D VGND VGND VPWR VPWR _33987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35726_ _35727_/CLK _35726_/D VGND VGND VPWR VPWR _35726_/Q sky130_fd_sc_hd__dfxtp_1
X_23740_ _22935_/X _32416_/Q _23742_/S VGND VGND VPWR VPWR _23741_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20952_ _22502_/A VGND VGND VPWR VPWR _20952_/X sky130_fd_sc_hd__buf_4
XFILLER_66_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32938_ _36075_/CLK _32938_/D VGND VGND VPWR VPWR _32938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35657_ _35848_/CLK _35657_/D VGND VGND VPWR VPWR _35657_/Q sky130_fd_sc_hd__dfxtp_1
X_23671_ _23671_/A VGND VGND VPWR VPWR _32384_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_98_CLK clkbuf_leaf_99_CLK/A VGND VGND VPWR VPWR _36196_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20883_ _22429_/A VGND VGND VPWR VPWR _20883_/X sky130_fd_sc_hd__buf_4
X_32869_ _36069_/CLK _32869_/D VGND VGND VPWR VPWR _32869_/Q sky130_fd_sc_hd__dfxtp_1
X_25410_ _25458_/S VGND VGND VPWR VPWR _25429_/S sky130_fd_sc_hd__buf_4
XFILLER_198_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22622_ _35589_/Q _35525_/Q _35461_/Q _35397_/Q _22556_/X _22557_/X VGND VGND VPWR
+ VPWR _22622_/X sky130_fd_sc_hd__mux4_1
X_34608_ _34797_/CLK _34608_/D VGND VGND VPWR VPWR _34608_/Q sky130_fd_sc_hd__dfxtp_1
X_26390_ _25153_/X _33602_/Q _26404_/S VGND VGND VPWR VPWR _26391_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35588_ _35715_/CLK _35588_/D VGND VGND VPWR VPWR _35588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25341_ _25013_/X _33109_/Q _25345_/S VGND VGND VPWR VPWR _25342_/A sky130_fd_sc_hd__mux2_1
X_22553_ _35843_/Q _32222_/Q _35715_/Q _35651_/Q _22266_/X _22267_/X VGND VGND VPWR
+ VPWR _22553_/X sky130_fd_sc_hd__mux4_1
X_34539_ _35944_/CLK _34539_/D VGND VGND VPWR VPWR _34539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28060_ _26956_/X _34361_/Q _28072_/S VGND VGND VPWR VPWR _28061_/A sky130_fd_sc_hd__mux2_1
X_21504_ _35301_/Q _35237_/Q _35173_/Q _32293_/Q _21253_/X _21254_/X VGND VGND VPWR
+ VPWR _21504_/X sky130_fd_sc_hd__mux4_1
X_25272_ _25112_/X _33077_/Q _25272_/S VGND VGND VPWR VPWR _25273_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_978 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22484_ _22480_/X _22483_/X _22442_/X _22443_/X VGND VGND VPWR VPWR _22499_/B sky130_fd_sc_hd__o211a_1
X_27011_ input58/X VGND VGND VPWR VPWR _27011_/X sky130_fd_sc_hd__buf_2
XFILLER_120_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36209_ _36211_/CLK _36209_/D VGND VGND VPWR VPWR _36209_/Q sky130_fd_sc_hd__dfxtp_1
X_24223_ _24223_/A VGND VGND VPWR VPWR _32643_/D sky130_fd_sc_hd__clkbuf_1
X_21435_ _21396_/X _21433_/X _21434_/X _21399_/X VGND VGND VPWR VPWR _21435_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24154_ _24154_/A VGND VGND VPWR VPWR _32610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21366_ _21366_/A VGND VGND VPWR VPWR _36193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23105_ input61/X VGND VGND VPWR VPWR _23105_/X sky130_fd_sc_hd__buf_6
X_20317_ _20069_/X _20315_/X _20316_/X _20073_/X VGND VGND VPWR VPWR _20317_/X sky130_fd_sc_hd__a22o_1
XFILLER_235_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24085_ _24085_/A VGND VGND VPWR VPWR _32578_/D sky130_fd_sc_hd__clkbuf_1
X_28962_ _28962_/A VGND VGND VPWR VPWR _34788_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_22_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _36201_/CLK sky130_fd_sc_hd__clkbuf_16
X_21297_ _21089_/X _21295_/X _21296_/X _21094_/X VGND VGND VPWR VPWR _21297_/X sky130_fd_sc_hd__a22o_1
XFILLER_235_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23036_ _23034_/X _32064_/Q _23063_/S VGND VGND VPWR VPWR _23037_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27913_ _27913_/A VGND VGND VPWR VPWR _34291_/D sky130_fd_sc_hd__clkbuf_1
X_20248_ _20061_/X _20246_/X _20247_/X _20067_/X VGND VGND VPWR VPWR _20248_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28893_ _26990_/X _34756_/Q _28903_/S VGND VGND VPWR VPWR _28894_/A sky130_fd_sc_hd__mux2_1
XTAP_5102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27844_ _27844_/A VGND VGND VPWR VPWR _34258_/D sky130_fd_sc_hd__clkbuf_1
X_20179_ _33281_/Q _36161_/Q _33153_/Q _33089_/Q _20064_/X _20065_/X VGND VGND VPWR
+ VPWR _20179_/X sky130_fd_sc_hd__mux4_1
XTAP_5135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24987_ _23074_/X _32973_/Q _24987_/S VGND VGND VPWR VPWR _24988_/A sky130_fd_sc_hd__mux2_1
XTAP_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27775_ _34226_/Q _24357_/X _27781_/S VGND VGND VPWR VPWR _27776_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29514_ _29514_/A VGND VGND VPWR VPWR _35019_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23938_ _23938_/A VGND VGND VPWR VPWR _32509_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26726_ _26726_/A VGND VGND VPWR VPWR _33760_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_700 _22458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_711 _22465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_722 _21473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26657_ _25146_/X _33728_/Q _26675_/S VGND VGND VPWR VPWR _26658_/A sky130_fd_sc_hd__mux2_1
XTAP_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29445_ _29445_/A VGND VGND VPWR VPWR _34986_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_733 _21191_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23869_ _23869_/A VGND VGND VPWR VPWR _32476_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_744 _22072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _35286_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_755 _22470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16410_ _16087_/X _16408_/X _16409_/X _16097_/X VGND VGND VPWR VPWR _16410_/X sky130_fd_sc_hd__a22o_1
XFILLER_72_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_766 _22511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25608_ _33232_/Q _24252_/X _25622_/S VGND VGND VPWR VPWR _25609_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17390_ _17352_/X _17388_/X _17389_/X _17355_/X VGND VGND VPWR VPWR _17390_/X sky130_fd_sc_hd__a22o_1
XANTENNA_777 _22604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29376_ _23336_/X _34954_/Q _29382_/S VGND VGND VPWR VPWR _29377_/A sky130_fd_sc_hd__mux2_1
X_26588_ _26588_/A VGND VGND VPWR VPWR _33695_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_788 _22663_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_799 _23075_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16341_ _16341_/A VGND VGND VPWR VPWR _31957_/D sky130_fd_sc_hd__clkbuf_1
X_28327_ _28327_/A VGND VGND VPWR VPWR _34487_/D sky130_fd_sc_hd__clkbuf_1
X_25539_ _33201_/Q _24354_/X _25547_/S VGND VGND VPWR VPWR _25540_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19060_ _18743_/X _19058_/X _19059_/X _18746_/X VGND VGND VPWR VPWR _19060_/X sky130_fd_sc_hd__a22o_1
X_16272_ _33748_/Q _33684_/Q _33620_/Q _33556_/Q _16137_/X _16138_/X VGND VGND VPWR
+ VPWR _16272_/X sky130_fd_sc_hd__mux4_1
X_28258_ _34455_/Q _24273_/X _28258_/S VGND VGND VPWR VPWR _28259_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18011_ _18007_/X _18010_/X _17834_/X VGND VGND VPWR VPWR _18033_/A sky130_fd_sc_hd__o21ba_2
X_27209_ _27209_/A VGND VGND VPWR VPWR _33958_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28189_ _26946_/X _34422_/Q _28207_/S VGND VGND VPWR VPWR _28190_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30220_ _30220_/A VGND VGND VPWR VPWR _35353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30151_ _35321_/Q _29185_/X _30163_/S VGND VGND VPWR VPWR _30152_/A sky130_fd_sc_hd__mux2_1
X_19962_ _32507_/Q _32379_/Q _32059_/Q _36027_/Q _19929_/X _19717_/X VGND VGND VPWR
+ VPWR _19962_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_13_CLK clkbuf_6_3__f_CLK/X VGND VGND VPWR VPWR _35929_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18913_ _33181_/Q _32541_/Q _35933_/Q _35869_/Q _18668_/X _18669_/X VGND VGND VPWR
+ VPWR _18913_/X sky130_fd_sc_hd__mux4_1
XTAP_7060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30082_ _35288_/Q _29082_/X _30100_/S VGND VGND VPWR VPWR _30083_/A sky130_fd_sc_hd__mux2_1
XTAP_7071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19893_ _32761_/Q _32697_/Q _32633_/Q _36089_/Q _19572_/X _19709_/X VGND VGND VPWR
+ VPWR _19893_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1110 _32122_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1121 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1132 _17908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33910_ _36150_/CLK _33910_/D VGND VGND VPWR VPWR _33910_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1143 _20232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18844_ _20256_/A VGND VGND VPWR VPWR _18844_/X sky130_fd_sc_hd__buf_4
X_34890_ _35340_/CLK _34890_/D VGND VGND VPWR VPWR _34890_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1154 _22455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1165 _22370_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1176 _22467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1187 _22503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33841_ _35760_/CLK _33841_/D VGND VGND VPWR VPWR _33841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1198 _22988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18775_ _18588_/X _18773_/X _18774_/X _18591_/X VGND VGND VPWR VPWR _18775_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15987_ _17906_/A VGND VGND VPWR VPWR _15987_/X sky130_fd_sc_hd__buf_4
XTAP_5680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17726_ _17846_/A VGND VGND VPWR VPWR _17726_/X sky130_fd_sc_hd__buf_4
X_33772_ _35315_/CLK _33772_/D VGND VGND VPWR VPWR _33772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30984_ _30984_/A VGND VGND VPWR VPWR _35715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35511_ _35638_/CLK _35511_/D VGND VGND VPWR VPWR _35511_/Q sky130_fd_sc_hd__dfxtp_1
X_32723_ _36052_/CLK _32723_/D VGND VGND VPWR VPWR _32723_/Q sky130_fd_sc_hd__dfxtp_1
X_17657_ _17555_/X _17655_/X _17656_/X _17558_/X VGND VGND VPWR VPWR _17657_/X sky130_fd_sc_hd__a22o_1
XFILLER_169_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16608_ _17796_/A VGND VGND VPWR VPWR _16608_/X sky130_fd_sc_hd__clkbuf_4
X_35442_ _36018_/CLK _35442_/D VGND VGND VPWR VPWR _35442_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_23__f_CLK clkbuf_5_11_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_23__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_32654_ _33234_/CLK _32654_/D VGND VGND VPWR VPWR _32654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17588_ _17548_/X _17586_/X _17587_/X _17553_/X VGND VGND VPWR VPWR _17588_/X sky130_fd_sc_hd__a22o_1
XFILLER_16_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31605_ _36010_/Q input21/X _31607_/S VGND VGND VPWR VPWR _31606_/A sky130_fd_sc_hd__mux2_1
X_19327_ _19002_/X _19325_/X _19326_/X _19008_/X VGND VGND VPWR VPWR _19327_/X sky130_fd_sc_hd__a22o_1
X_16539_ _16357_/X _16537_/X _16538_/X _16361_/X VGND VGND VPWR VPWR _16539_/X sky130_fd_sc_hd__a22o_1
X_35373_ _35946_/CLK _35373_/D VGND VGND VPWR VPWR _35373_/Q sky130_fd_sc_hd__dfxtp_1
X_32585_ _35977_/CLK _32585_/D VGND VGND VPWR VPWR _32585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34324_ _35031_/CLK _34324_/D VGND VGND VPWR VPWR _34324_/Q sky130_fd_sc_hd__dfxtp_1
X_31536_ _31536_/A VGND VGND VPWR VPWR _35977_/D sky130_fd_sc_hd__clkbuf_1
X_19258_ _19010_/X _19256_/X _19257_/X _19014_/X VGND VGND VPWR VPWR _19258_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18209_ _34571_/Q _32459_/Q _34443_/Q _34379_/Q _17931_/X _17932_/X VGND VGND VPWR
+ VPWR _18209_/X sky130_fd_sc_hd__mux4_1
X_34255_ _34256_/CLK _34255_/D VGND VGND VPWR VPWR _34255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31467_ _31467_/A VGND VGND VPWR VPWR _35944_/D sky130_fd_sc_hd__clkbuf_1
X_19189_ _19002_/X _19187_/X _19188_/X _19008_/X VGND VGND VPWR VPWR _19189_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21220_ _35037_/Q _34973_/Q _34909_/Q _34845_/Q _21050_/X _21051_/X VGND VGND VPWR
+ VPWR _21220_/X sky130_fd_sc_hd__mux4_1
X_33206_ _36022_/CLK _33206_/D VGND VGND VPWR VPWR _33206_/Q sky130_fd_sc_hd__dfxtp_1
X_30418_ _23274_/X _35447_/Q _30434_/S VGND VGND VPWR VPWR _30419_/A sky130_fd_sc_hd__mux2_1
X_34186_ _35851_/CLK _34186_/D VGND VGND VPWR VPWR _34186_/Q sky130_fd_sc_hd__dfxtp_1
X_31398_ _35912_/Q input54/X _31400_/S VGND VGND VPWR VPWR _31399_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33137_ _33520_/CLK _33137_/D VGND VGND VPWR VPWR _33137_/Q sky130_fd_sc_hd__dfxtp_1
X_21151_ _35291_/Q _35227_/Q _35163_/Q _32283_/Q _20900_/X _20901_/X VGND VGND VPWR
+ VPWR _21151_/X sky130_fd_sc_hd__mux4_1
X_30349_ _30349_/A VGND VGND VPWR VPWR _35414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20102_ _20098_/X _20101_/X _19781_/X VGND VGND VPWR VPWR _20124_/A sky130_fd_sc_hd__o21ba_1
XFILLER_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21082_ _21043_/X _21080_/X _21081_/X _21046_/X VGND VGND VPWR VPWR _21082_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33068_ _36076_/CLK _33068_/D VGND VGND VPWR VPWR _33068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20033_ _19708_/X _20031_/X _20032_/X _19714_/X VGND VGND VPWR VPWR _20033_/X sky130_fd_sc_hd__a22o_1
X_24910_ _22960_/X _32936_/Q _24916_/S VGND VGND VPWR VPWR _24911_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32019_ _35986_/CLK _32019_/D VGND VGND VPWR VPWR _32019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25890_ _25013_/X _33365_/Q _25894_/S VGND VGND VPWR VPWR _25891_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24841_ _24841_/A VGND VGND VPWR VPWR _32903_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27560_ _27560_/A VGND VGND VPWR VPWR _34125_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24772_ _24772_/A VGND VGND VPWR VPWR _32870_/D sky130_fd_sc_hd__clkbuf_1
X_21984_ _21980_/X _21983_/X _21736_/X _21737_/X VGND VGND VPWR VPWR _21999_/B sky130_fd_sc_hd__o211a_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26511_ _26511_/A VGND VGND VPWR VPWR _33659_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35709_ _35709_/CLK _35709_/D VGND VGND VPWR VPWR _35709_/Q sky130_fd_sc_hd__dfxtp_1
X_23723_ _23834_/S VGND VGND VPWR VPWR _23742_/S sky130_fd_sc_hd__buf_4
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20935_ _20674_/X _20933_/X _20934_/X _20684_/X VGND VGND VPWR VPWR _20935_/X sky130_fd_sc_hd__a22o_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27491_ _26915_/X _34092_/Q _27509_/S VGND VGND VPWR VPWR _27492_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29230_ _29230_/A VGND VGND VPWR VPWR _34887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26442_ _26442_/A VGND VGND VPWR VPWR _33626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23654_ _23654_/A VGND VGND VPWR VPWR _32376_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20866_ _34515_/Q _32403_/Q _34387_/Q _34323_/Q _20766_/X _20767_/X VGND VGND VPWR
+ VPWR _20866_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22605_ _33797_/Q _33733_/Q _33669_/Q _33605_/Q _22502_/X _22503_/X VGND VGND VPWR
+ VPWR _22605_/X sky130_fd_sc_hd__mux4_1
X_29161_ _34865_/Q _29160_/X _29173_/S VGND VGND VPWR VPWR _29162_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26373_ _25128_/X _33594_/Q _26383_/S VGND VGND VPWR VPWR _26374_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23585_ _23696_/S VGND VGND VPWR VPWR _23604_/S sky130_fd_sc_hd__buf_4
X_20797_ _34769_/Q _34705_/Q _34641_/Q _34577_/Q _20675_/X _20676_/X VGND VGND VPWR
+ VPWR _20797_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28112_ _28112_/A VGND VGND VPWR VPWR _34385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25324_ _31680_/A _27561_/B VGND VGND VPWR VPWR _28643_/B sky130_fd_sc_hd__nor2_8
XFILLER_139_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22536_ _22530_/X _22535_/X _22467_/X VGND VGND VPWR VPWR _22537_/D sky130_fd_sc_hd__o21ba_1
X_29092_ input5/X VGND VGND VPWR VPWR _29092_/X sky130_fd_sc_hd__buf_4
XFILLER_122_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28043_ _26931_/X _34353_/Q _28051_/S VGND VGND VPWR VPWR _28044_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25255_ _25255_/A VGND VGND VPWR VPWR _33068_/D sky130_fd_sc_hd__clkbuf_1
X_22467_ _22467_/A VGND VGND VPWR VPWR _22467_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_183_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24206_ _24206_/A VGND VGND VPWR VPWR _32635_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21418_ _21414_/X _21417_/X _21375_/X VGND VGND VPWR VPWR _21440_/A sky130_fd_sc_hd__o21ba_1
X_25186_ input60/X VGND VGND VPWR VPWR _25186_/X sky130_fd_sc_hd__buf_2
X_22398_ _22148_/X _22394_/X _22397_/X _22153_/X VGND VGND VPWR VPWR _22398_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24137_ _24137_/A VGND VGND VPWR VPWR _32602_/D sky130_fd_sc_hd__clkbuf_1
X_21349_ _21310_/X _21347_/X _21348_/X _21314_/X VGND VGND VPWR VPWR _21349_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29994_ _29994_/A VGND VGND VPWR VPWR _35246_/D sky130_fd_sc_hd__clkbuf_1
X_24068_ _24068_/A VGND VGND VPWR VPWR _32570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28945_ _28945_/A VGND VGND VPWR VPWR _34780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23019_ input40/X VGND VGND VPWR VPWR _23019_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28876_ _26965_/X _34748_/Q _28882_/S VGND VGND VPWR VPWR _28877_/A sky130_fd_sc_hd__mux2_1
X_16890_ _32485_/Q _32357_/Q _32037_/Q _36005_/Q _16570_/X _16711_/X VGND VGND VPWR
+ VPWR _16890_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27827_ _34251_/Q _24434_/X _27831_/S VGND VGND VPWR VPWR _27828_/A sky130_fd_sc_hd__mux2_1
XTAP_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18560_ _33171_/Q _32531_/Q _35923_/Q _35859_/Q _18363_/X _18365_/X VGND VGND VPWR
+ VPWR _18560_/X sky130_fd_sc_hd__mux4_1
XTAP_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_24_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_24_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XTAP_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27758_ _34218_/Q _24332_/X _27760_/S VGND VGND VPWR VPWR _27759_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17511_ _35062_/Q _34998_/Q _34934_/Q _34870_/Q _17509_/X _17510_/X VGND VGND VPWR
+ VPWR _17511_/X sky130_fd_sc_hd__mux4_1
XTAP_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26709_ _33752_/Q _24276_/X _26727_/S VGND VGND VPWR VPWR _26710_/A sky130_fd_sc_hd__mux2_1
X_18491_ _20146_/A VGND VGND VPWR VPWR _18491_/X sky130_fd_sc_hd__buf_6
XTAP_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27689_ _27689_/A VGND VGND VPWR VPWR _34185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_530 _18184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_541 _20256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17442_ _17956_/A VGND VGND VPWR VPWR _17442_/X sky130_fd_sc_hd__buf_4
X_29428_ _23148_/X _34978_/Q _29446_/S VGND VGND VPWR VPWR _29429_/A sky130_fd_sc_hd__mux2_1
XANTENNA_552 _20142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_563 _18358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _35294_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_574 _20165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_585 _19452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_596 _19459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29359_ _29359_/A VGND VGND VPWR VPWR _34945_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17373_ _17846_/A VGND VGND VPWR VPWR _17373_/X sky130_fd_sc_hd__buf_4
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19112_ _33763_/Q _33699_/Q _33635_/Q _33571_/Q _18790_/X _18791_/X VGND VGND VPWR
+ VPWR _19112_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16324_ _16026_/X _16322_/X _16323_/X _16037_/X VGND VGND VPWR VPWR _16324_/X sky130_fd_sc_hd__a22o_1
XFILLER_242_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32370_ _36018_/CLK _32370_/D VGND VGND VPWR VPWR _32370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16255_ _17796_/A VGND VGND VPWR VPWR _16255_/X sky130_fd_sc_hd__buf_4
X_31321_ _35875_/Q input14/X _31337_/S VGND VGND VPWR VPWR _31322_/A sky130_fd_sc_hd__mux2_1
X_19043_ _19039_/X _19042_/X _18722_/X VGND VGND VPWR VPWR _19065_/A sky130_fd_sc_hd__o21ba_2
XFILLER_51_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31252_ _31252_/A VGND VGND VPWR VPWR _35842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34040_ _36152_/CLK _34040_/D VGND VGND VPWR VPWR _34040_/Q sky130_fd_sc_hd__dfxtp_1
X_16186_ _16026_/X _16184_/X _16185_/X _16037_/X VGND VGND VPWR VPWR _16186_/X sky130_fd_sc_hd__a22o_1
Xoutput206 _36231_/Q VGND VGND VPWR VPWR D2[57] sky130_fd_sc_hd__buf_2
XFILLER_182_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput217 _36183_/Q VGND VGND VPWR VPWR D2[9] sky130_fd_sc_hd__buf_2
XFILLER_138_1303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30203_ _30203_/A VGND VGND VPWR VPWR _35345_/D sky130_fd_sc_hd__clkbuf_1
Xoutput228 _32097_/Q VGND VGND VPWR VPWR D3[19] sky130_fd_sc_hd__buf_2
X_31183_ _31273_/S VGND VGND VPWR VPWR _31202_/S sky130_fd_sc_hd__buf_4
XFILLER_154_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput239 _32107_/Q VGND VGND VPWR VPWR D3[29] sky130_fd_sc_hd__buf_2
XFILLER_47_1219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30134_ _35313_/Q _29160_/X _30142_/S VGND VGND VPWR VPWR _30135_/A sky130_fd_sc_hd__mux2_1
X_19945_ _19802_/X _19943_/X _19944_/X _19805_/X VGND VGND VPWR VPWR _19945_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35991_ _35991_/CLK _35991_/D VGND VGND VPWR VPWR _35991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30065_ _35280_/Q _29058_/X _30079_/S VGND VGND VPWR VPWR _30066_/A sky130_fd_sc_hd__mux2_1
X_34942_ _35517_/CLK _34942_/D VGND VGND VPWR VPWR _34942_/Q sky130_fd_sc_hd__dfxtp_1
X_19876_ _35320_/Q _35256_/Q _35192_/Q _32312_/Q _19659_/X _19660_/X VGND VGND VPWR
+ VPWR _19876_/X sky130_fd_sc_hd__mux4_1
XFILLER_214_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_1279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18827_ _33755_/Q _33691_/Q _33627_/Q _33563_/Q _18790_/X _18791_/X VGND VGND VPWR
+ VPWR _18827_/X sky130_fd_sc_hd__mux4_1
X_34873_ _35386_/CLK _34873_/D VGND VGND VPWR VPWR _34873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33824_ _35745_/CLK _33824_/D VGND VGND VPWR VPWR _33824_/Q sky130_fd_sc_hd__dfxtp_1
X_18758_ _18758_/A VGND VGND VPWR VPWR _32088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17709_ _17705_/X _17706_/X _17707_/X _17708_/X VGND VGND VPWR VPWR _17709_/X sky130_fd_sc_hd__a22o_1
X_33755_ _34266_/CLK _33755_/D VGND VGND VPWR VPWR _33755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18689_ _18443_/X _18687_/X _18688_/X _18446_/X VGND VGND VPWR VPWR _18689_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30967_ _30967_/A VGND VGND VPWR VPWR _35707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20720_ _35791_/Q _32165_/Q _35663_/Q _35599_/Q _20645_/X _20646_/X VGND VGND VPWR
+ VPWR _20720_/X sky130_fd_sc_hd__mux4_1
X_32706_ _33026_/CLK _32706_/D VGND VGND VPWR VPWR _32706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33686_ _34260_/CLK _33686_/D VGND VGND VPWR VPWR _33686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30898_ _30898_/A VGND VGND VPWR VPWR _35674_/D sky130_fd_sc_hd__clkbuf_1
X_35425_ _35808_/CLK _35425_/D VGND VGND VPWR VPWR _35425_/Q sky130_fd_sc_hd__dfxtp_1
X_20651_ _22595_/A VGND VGND VPWR VPWR _20651_/X sky130_fd_sc_hd__clkbuf_4
X_32637_ _36092_/CLK _32637_/D VGND VGND VPWR VPWR _32637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35356_ _35869_/CLK _35356_/D VGND VGND VPWR VPWR _35356_/Q sky130_fd_sc_hd__dfxtp_1
X_23370_ _23370_/A VGND VGND VPWR VPWR _32244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20582_ _20659_/A VGND VGND VPWR VPWR _22503_/A sky130_fd_sc_hd__buf_12
X_32568_ _36024_/CLK _32568_/D VGND VGND VPWR VPWR _32568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34307_ _34310_/CLK _34307_/D VGND VGND VPWR VPWR _34307_/Q sky130_fd_sc_hd__dfxtp_1
X_22321_ _22321_/A VGND VGND VPWR VPWR _36220_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31519_ _23307_/X _35969_/Q _31535_/S VGND VGND VPWR VPWR _31520_/A sky130_fd_sc_hd__mux2_1
X_35287_ _36191_/CLK _35287_/D VGND VGND VPWR VPWR _35287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32499_ _36019_/CLK _32499_/D VGND VGND VPWR VPWR _32499_/Q sky130_fd_sc_hd__dfxtp_1
X_25040_ _25040_/A VGND VGND VPWR VPWR _32989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34238_ _34302_/CLK _34238_/D VGND VGND VPWR VPWR _34238_/Q sky130_fd_sc_hd__dfxtp_1
X_22252_ _33787_/Q _33723_/Q _33659_/Q _33595_/Q _22149_/X _22150_/X VGND VGND VPWR
+ VPWR _22252_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21203_ _32477_/Q _32349_/Q _32029_/Q _35997_/Q _21170_/X _20958_/X VGND VGND VPWR
+ VPWR _21203_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22183_ _22177_/X _22182_/X _22114_/X VGND VGND VPWR VPWR _22184_/D sky130_fd_sc_hd__o21ba_1
X_34169_ _36152_/CLK _34169_/D VGND VGND VPWR VPWR _34169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21134_ _32731_/Q _32667_/Q _32603_/Q _36059_/Q _20813_/X _20950_/X VGND VGND VPWR
+ VPWR _21134_/X sky130_fd_sc_hd__mux4_1
X_26991_ _26990_/X _33860_/Q _27006_/S VGND VGND VPWR VPWR _26992_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28730_ _28730_/A VGND VGND VPWR VPWR _34678_/D sky130_fd_sc_hd__clkbuf_1
X_21065_ _21061_/X _21064_/X _21022_/X VGND VGND VPWR VPWR _21087_/A sky130_fd_sc_hd__o21ba_1
X_25942_ _25942_/A VGND VGND VPWR VPWR _33389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20016_ _34556_/Q _32444_/Q _34428_/Q _34364_/Q _19878_/X _19879_/X VGND VGND VPWR
+ VPWR _20016_/X sky130_fd_sc_hd__mux4_1
X_25873_ _25873_/A VGND VGND VPWR VPWR _33357_/D sky130_fd_sc_hd__clkbuf_1
X_28661_ _26847_/X _34646_/Q _28663_/S VGND VGND VPWR VPWR _28662_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24824_ _24824_/A VGND VGND VPWR VPWR _32895_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27612_ _27612_/A VGND VGND VPWR VPWR _34148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28592_ _28592_/A VGND VGND VPWR VPWR _34613_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27543_ _26993_/X _34117_/Q _27551_/S VGND VGND VPWR VPWR _27544_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24755_ _24755_/A VGND VGND VPWR VPWR _32862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21967_ _21967_/A _21967_/B _21967_/C _21967_/D VGND VGND VPWR VPWR _21968_/A sky130_fd_sc_hd__or4_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23706_ _23706_/A VGND VGND VPWR VPWR _32399_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20918_ _20912_/X _20917_/X _20611_/X VGND VGND VPWR VPWR _20940_/A sky130_fd_sc_hd__o21ba_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27474_ _26891_/X _34084_/Q _27488_/S VGND VGND VPWR VPWR _27475_/A sky130_fd_sc_hd__mux2_1
X_24686_ _23031_/X _32831_/Q _24686_/S VGND VGND VPWR VPWR _24687_/A sky130_fd_sc_hd__mux2_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21898_ _21898_/A VGND VGND VPWR VPWR _36208_/D sky130_fd_sc_hd__buf_6
XFILLER_202_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29213_ input48/X VGND VGND VPWR VPWR _29213_/X sky130_fd_sc_hd__buf_4
XFILLER_9_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26425_ _26425_/A VGND VGND VPWR VPWR _33618_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23637_ _23637_/A VGND VGND VPWR VPWR _32368_/D sky130_fd_sc_hd__clkbuf_1
X_20849_ _20614_/X _20847_/X _20848_/X _20623_/X VGND VGND VPWR VPWR _20849_/X sky130_fd_sc_hd__a22o_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29144_ input24/X VGND VGND VPWR VPWR _29144_/X sky130_fd_sc_hd__clkbuf_4
X_26356_ _25103_/X _33586_/Q _26362_/S VGND VGND VPWR VPWR _26357_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23568_ _23568_/A VGND VGND VPWR VPWR _32335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25307_ _25307_/A VGND VGND VPWR VPWR _33093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22519_ _22369_/X _22517_/X _22518_/X _22373_/X VGND VGND VPWR VPWR _22519_/X sky130_fd_sc_hd__a22o_1
X_26287_ _25001_/X _33553_/Q _26299_/S VGND VGND VPWR VPWR _26288_/A sky130_fd_sc_hd__mux2_1
X_29075_ _29075_/A VGND VGND VPWR VPWR _34837_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23499_ _22985_/X _32304_/Q _23509_/S VGND VGND VPWR VPWR _23500_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16040_ _17842_/A VGND VGND VPWR VPWR _16040_/X sky130_fd_sc_hd__buf_2
XFILLER_10_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28026_ _26906_/X _34345_/Q _28030_/S VGND VGND VPWR VPWR _28027_/A sky130_fd_sc_hd__mux2_1
X_25238_ _25238_/A VGND VGND VPWR VPWR _33060_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25169_ _25168_/X _33031_/Q _25175_/S VGND VGND VPWR VPWR _25170_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17991_ _33220_/Q _32580_/Q _35972_/Q _35908_/Q _17780_/X _17781_/X VGND VGND VPWR
+ VPWR _17991_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29977_ _29977_/A VGND VGND VPWR VPWR _35238_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19730_ _19652_/X _19726_/X _19729_/X _19655_/X VGND VGND VPWR VPWR _19730_/X sky130_fd_sc_hd__a22o_1
X_28928_ _28928_/A VGND VGND VPWR VPWR _34772_/D sky130_fd_sc_hd__clkbuf_1
X_16942_ _16801_/X _16940_/X _16941_/X _16806_/X VGND VGND VPWR VPWR _16942_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19661_ _35314_/Q _35250_/Q _35186_/Q _32306_/Q _19659_/X _19660_/X VGND VGND VPWR
+ VPWR _19661_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16873_ _16873_/A VGND VGND VPWR VPWR _16873_/X sky130_fd_sc_hd__buf_4
X_28859_ _26940_/X _34740_/Q _28861_/S VGND VGND VPWR VPWR _28860_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18612_ _18436_/X _18610_/X _18611_/X _18441_/X VGND VGND VPWR VPWR _18612_/X sky130_fd_sc_hd__a22o_1
XTAP_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19592_ _19449_/X _19590_/X _19591_/X _19452_/X VGND VGND VPWR VPWR _19592_/X sky130_fd_sc_hd__a22o_1
X_31870_ _31870_/A VGND VGND VPWR VPWR _36135_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ _33491_/Q _33427_/Q _33363_/Q _33299_/Q _18298_/X _18299_/X VGND VGND VPWR
+ VPWR _18543_/X sky130_fd_sc_hd__mux4_1
XTAP_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30821_ _23270_/X _35638_/Q _30839_/S VGND VGND VPWR VPWR _30822_/A sky130_fd_sc_hd__mux2_1
XTAP_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33540_ _33545_/CLK _33540_/D VGND VGND VPWR VPWR _33540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18474_ _33745_/Q _33681_/Q _33617_/Q _33553_/Q _18437_/X _18438_/X VGND VGND VPWR
+ VPWR _18474_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30752_ _30752_/A VGND VGND VPWR VPWR _35605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_360 _36207_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_371 _36208_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_382 _36209_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17425_ _17347_/X _17423_/X _17424_/X _17350_/X VGND VGND VPWR VPWR _17425_/X sky130_fd_sc_hd__a22o_1
XANTENNA_393 _36209_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33471_ _34303_/CLK _33471_/D VGND VGND VPWR VPWR _33471_/Q sky130_fd_sc_hd__dfxtp_1
X_30683_ _35573_/Q _29172_/X _30683_/S VGND VGND VPWR VPWR _30684_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35210_ _35338_/CLK _35210_/D VGND VGND VPWR VPWR _35210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32422_ _35942_/CLK _32422_/D VGND VGND VPWR VPWR _32422_/Q sky130_fd_sc_hd__dfxtp_1
X_36190_ _36194_/CLK _36190_/D VGND VGND VPWR VPWR _36190_/Q sky130_fd_sc_hd__dfxtp_1
X_17356_ _17352_/X _17353_/X _17354_/X _17355_/X VGND VGND VPWR VPWR _17356_/X sky130_fd_sc_hd__a22o_1
XFILLER_207_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35141_ _35845_/CLK _35141_/D VGND VGND VPWR VPWR _35141_/Q sky130_fd_sc_hd__dfxtp_1
X_16307_ _16303_/X _16306_/X _16100_/X VGND VGND VPWR VPWR _16308_/D sky130_fd_sc_hd__o21ba_1
XFILLER_53_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32353_ _36001_/CLK _32353_/D VGND VGND VPWR VPWR _32353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17287_ _17283_/X _17286_/X _17147_/X VGND VGND VPWR VPWR _17297_/C sky130_fd_sc_hd__o21ba_1
XFILLER_174_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19026_ _34784_/Q _34720_/Q _34656_/Q _34592_/Q _18882_/X _18883_/X VGND VGND VPWR
+ VPWR _19026_/X sky130_fd_sc_hd__mux4_1
X_31304_ _35867_/Q input5/X _31316_/S VGND VGND VPWR VPWR _31305_/A sky130_fd_sc_hd__mux2_1
X_35072_ _35075_/CLK _35072_/D VGND VGND VPWR VPWR _35072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16238_ _16238_/A _16238_/B _16238_/C _16238_/D VGND VGND VPWR VPWR _16239_/A sky130_fd_sc_hd__or4_4
X_32284_ _35164_/CLK _32284_/D VGND VGND VPWR VPWR _32284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34023_ _34153_/CLK _34023_/D VGND VGND VPWR VPWR _34023_/Q sky130_fd_sc_hd__dfxtp_1
X_31235_ _31235_/A VGND VGND VPWR VPWR _35834_/D sky130_fd_sc_hd__clkbuf_1
X_16169_ _35024_/Q _34960_/Q _34896_/Q _34832_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _16169_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31166_ _31166_/A VGND VGND VPWR VPWR _35801_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19928_ _19708_/X _19926_/X _19927_/X _19714_/X VGND VGND VPWR VPWR _19928_/X sky130_fd_sc_hd__a22o_1
X_30117_ _35305_/Q _29135_/X _30121_/S VGND VGND VPWR VPWR _30118_/A sky130_fd_sc_hd__mux2_1
X_35974_ _35975_/CLK _35974_/D VGND VGND VPWR VPWR _35974_/Q sky130_fd_sc_hd__dfxtp_1
X_31097_ _35769_/Q _29185_/X _31109_/S VGND VGND VPWR VPWR _31098_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30048_ _30048_/A VGND VGND VPWR VPWR _35272_/D sky130_fd_sc_hd__clkbuf_1
X_34925_ _35757_/CLK _34925_/D VGND VGND VPWR VPWR _34925_/Q sky130_fd_sc_hd__dfxtp_1
X_19859_ _19855_/X _19856_/X _19857_/X _19858_/X VGND VGND VPWR VPWR _19859_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22870_ _35085_/Q _35021_/Q _34957_/Q _34893_/Q _20679_/X _20681_/X VGND VGND VPWR
+ VPWR _22870_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34856_ _34987_/CLK _34856_/D VGND VGND VPWR VPWR _34856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33807_ _35728_/CLK _33807_/D VGND VGND VPWR VPWR _33807_/Q sky130_fd_sc_hd__dfxtp_1
X_21821_ _21817_/X _21820_/X _21747_/X VGND VGND VPWR VPWR _21831_/C sky130_fd_sc_hd__o21ba_1
XFILLER_43_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34787_ _35928_/CLK _34787_/D VGND VGND VPWR VPWR _34787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31999_ _33946_/CLK _31999_/D VGND VGND VPWR VPWR _31999_/Q sky130_fd_sc_hd__dfxtp_1
X_24540_ _23019_/X _32763_/Q _24548_/S VGND VGND VPWR VPWR _24541_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33738_ _35977_/CLK _33738_/D VGND VGND VPWR VPWR _33738_/Q sky130_fd_sc_hd__dfxtp_1
X_21752_ _21752_/A VGND VGND VPWR VPWR _21752_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_224_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20703_ _20703_/A VGND VGND VPWR VPWR _36174_/D sky130_fd_sc_hd__clkbuf_1
X_24471_ _22917_/X _32730_/Q _24485_/S VGND VGND VPWR VPWR _24472_/A sky130_fd_sc_hd__mux2_1
X_33669_ _34309_/CLK _33669_/D VGND VGND VPWR VPWR _33669_/Q sky130_fd_sc_hd__dfxtp_1
X_21683_ _35050_/Q _34986_/Q _34922_/Q _34858_/Q _21403_/X _21404_/X VGND VGND VPWR
+ VPWR _21683_/X sky130_fd_sc_hd__mux4_1
X_26210_ _26210_/A VGND VGND VPWR VPWR _33516_/D sky130_fd_sc_hd__clkbuf_1
X_23422_ _23422_/A VGND VGND VPWR VPWR _32269_/D sky130_fd_sc_hd__clkbuf_1
X_35408_ _35793_/CLK _35408_/D VGND VGND VPWR VPWR _35408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20634_ _20659_/A VGND VGND VPWR VPWR _22430_/A sky130_fd_sc_hd__buf_12
X_27190_ _27190_/A VGND VGND VPWR VPWR _33949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26141_ _26141_/A VGND VGND VPWR VPWR _33484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35339_ _35339_/CLK _35339_/D VGND VGND VPWR VPWR _35339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23353_ _32236_/Q _23237_/X _23371_/S VGND VGND VPWR VPWR _23354_/A sky130_fd_sc_hd__mux2_1
X_20565_ _20561_/X _20564_/X _20153_/A VGND VGND VPWR VPWR _20573_/C sky130_fd_sc_hd__o21ba_1
X_22304_ _22300_/X _22301_/X _22302_/X _22303_/X VGND VGND VPWR VPWR _22304_/X sky130_fd_sc_hd__a22o_1
XFILLER_153_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26072_ _26072_/A VGND VGND VPWR VPWR _33451_/D sky130_fd_sc_hd__clkbuf_1
X_23284_ _32212_/Q _23283_/X _23301_/S VGND VGND VPWR VPWR _23285_/A sky130_fd_sc_hd__mux2_1
X_20496_ _33035_/Q _32971_/Q _32907_/Q _32843_/Q _18280_/X _18283_/X VGND VGND VPWR
+ VPWR _20496_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29900_ _35202_/Q _29213_/X _29914_/S VGND VGND VPWR VPWR _29901_/A sky130_fd_sc_hd__mux2_1
X_25023_ _25187_/S VGND VGND VPWR VPWR _25051_/S sky130_fd_sc_hd__buf_4
XFILLER_164_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22235_ _35770_/Q _35130_/Q _34490_/Q _33850_/Q _22093_/X _22094_/X VGND VGND VPWR
+ VPWR _22235_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29831_ _29831_/A VGND VGND VPWR VPWR _35169_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22166_ _22016_/X _22164_/X _22165_/X _22020_/X VGND VGND VPWR VPWR _22166_/X sky130_fd_sc_hd__a22o_1
XFILLER_79_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21117_ _35290_/Q _35226_/Q _35162_/Q _32282_/Q _20900_/X _20901_/X VGND VGND VPWR
+ VPWR _21117_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29762_ _29762_/A VGND VGND VPWR VPWR _35136_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26974_ input44/X VGND VGND VPWR VPWR _26974_/X sky130_fd_sc_hd__clkbuf_4
X_22097_ _35574_/Q _35510_/Q _35446_/Q _35382_/Q _21850_/X _21851_/X VGND VGND VPWR
+ VPWR _22097_/X sky130_fd_sc_hd__mux4_1
XTAP_6969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28713_ _28713_/A VGND VGND VPWR VPWR _34670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25925_ _25925_/A VGND VGND VPWR VPWR _33381_/D sky130_fd_sc_hd__clkbuf_1
X_21048_ _21754_/A VGND VGND VPWR VPWR _21048_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_59_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29693_ _35104_/Q _29107_/X _29695_/S VGND VGND VPWR VPWR _29694_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28644_ _28776_/S VGND VGND VPWR VPWR _28663_/S sky130_fd_sc_hd__buf_6
X_25856_ _25162_/X _33349_/Q _25864_/S VGND VGND VPWR VPWR _25857_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24807_ _23007_/X _32887_/Q _24823_/S VGND VGND VPWR VPWR _24808_/A sky130_fd_sc_hd__mux2_1
X_28575_ _26919_/X _34605_/Q _28591_/S VGND VGND VPWR VPWR _28576_/A sky130_fd_sc_hd__mux2_1
X_25787_ _25060_/X _33316_/Q _25801_/S VGND VGND VPWR VPWR _25788_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22999_ _22999_/A VGND VGND VPWR VPWR _32052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27526_ _26968_/X _34109_/Q _27530_/S VGND VGND VPWR VPWR _27527_/A sky130_fd_sc_hd__mux2_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24738_ _24738_/A VGND VGND VPWR VPWR _32854_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27457_ _26866_/X _34076_/Q _27467_/S VGND VGND VPWR VPWR _27458_/A sky130_fd_sc_hd__mux2_1
X_24669_ _24669_/A VGND VGND VPWR VPWR _32822_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17210_ _17055_/X _17208_/X _17209_/X _17061_/X VGND VGND VPWR VPWR _17210_/X sky130_fd_sc_hd__a22o_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26408_ _25180_/X _33611_/Q _26412_/S VGND VGND VPWR VPWR _26409_/A sky130_fd_sc_hd__mux2_1
X_18190_ _17908_/X _18188_/X _18189_/X _17911_/X VGND VGND VPWR VPWR _18190_/X sky130_fd_sc_hd__a22o_1
XFILLER_129_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27388_ _27388_/A VGND VGND VPWR VPWR _34043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1070 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17141_ _17995_/A VGND VGND VPWR VPWR _17141_/X sky130_fd_sc_hd__buf_4
X_29127_ _34854_/Q _29126_/X _29142_/S VGND VGND VPWR VPWR _29128_/A sky130_fd_sc_hd__mux2_1
X_26339_ _25078_/X _33578_/Q _26341_/S VGND VGND VPWR VPWR _26340_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17072_ _16994_/X _17070_/X _17071_/X _16997_/X VGND VGND VPWR VPWR _17072_/X sky130_fd_sc_hd__a22o_1
X_29058_ input23/X VGND VGND VPWR VPWR _29058_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_196_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16023_ _17906_/A VGND VGND VPWR VPWR _16023_/X sky130_fd_sc_hd__buf_2
X_28009_ _26881_/X _34337_/Q _28009_/S VGND VGND VPWR VPWR _28010_/A sky130_fd_sc_hd__mux2_1
X_31020_ _31020_/A VGND VGND VPWR VPWR _35732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17974_ _33540_/Q _33476_/Q _33412_/Q _33348_/Q _17829_/X _17830_/X VGND VGND VPWR
+ VPWR _17974_/X sky130_fd_sc_hd__mux4_1
X_19713_ _33268_/Q _36148_/Q _33140_/Q _33076_/Q _19711_/X _19712_/X VGND VGND VPWR
+ VPWR _19713_/X sky130_fd_sc_hd__mux4_1
X_16925_ _32998_/Q _32934_/Q _32870_/Q _32806_/Q _16636_/X _16637_/X VGND VGND VPWR
+ VPWR _16925_/X sky130_fd_sc_hd__mux4_1
X_32971_ _34251_/CLK _32971_/D VGND VGND VPWR VPWR _32971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_293_CLK clkbuf_6_51__f_CLK/X VGND VGND VPWR VPWR _36032_/CLK sky130_fd_sc_hd__clkbuf_16
X_34710_ _35669_/CLK _34710_/D VGND VGND VPWR VPWR _34710_/Q sky130_fd_sc_hd__dfxtp_1
X_31922_ _23303_/X _36160_/Q _31940_/S VGND VGND VPWR VPWR _31923_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19644_ _33010_/Q _32946_/Q _32882_/Q _32818_/Q _19642_/X _19643_/X VGND VGND VPWR
+ VPWR _19644_/X sky130_fd_sc_hd__mux4_1
X_35690_ _35818_/CLK _35690_/D VGND VGND VPWR VPWR _35690_/Q sky130_fd_sc_hd__dfxtp_1
X_16856_ _33252_/Q _36132_/Q _33124_/Q _33060_/Q _16705_/X _16706_/X VGND VGND VPWR
+ VPWR _16856_/X sky130_fd_sc_hd__mux4_1
X_34641_ _36220_/CLK _34641_/D VGND VGND VPWR VPWR _34641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19575_ _19355_/X _19573_/X _19574_/X _19361_/X VGND VGND VPWR VPWR _19575_/X sky130_fd_sc_hd__a22o_1
XFILLER_19_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31853_ _31853_/A VGND VGND VPWR VPWR _36127_/D sky130_fd_sc_hd__clkbuf_1
X_16787_ _17994_/A VGND VGND VPWR VPWR _16787_/X sky130_fd_sc_hd__buf_6
XFILLER_4_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18526_ _33170_/Q _32530_/Q _35922_/Q _35858_/Q _18363_/X _18365_/X VGND VGND VPWR
+ VPWR _18526_/X sky130_fd_sc_hd__mux4_1
X_30804_ _23244_/X _35630_/Q _30818_/S VGND VGND VPWR VPWR _30805_/A sky130_fd_sc_hd__mux2_1
X_34572_ _35981_/CLK _34572_/D VGND VGND VPWR VPWR _34572_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31784_ _36095_/Q input44/X _31784_/S VGND VGND VPWR VPWR _31785_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33523_ _33779_/CLK _33523_/D VGND VGND VPWR VPWR _33523_/Q sky130_fd_sc_hd__dfxtp_1
X_30735_ _30735_/A _30735_/B VGND VGND VPWR VPWR _30868_/S sky130_fd_sc_hd__nand2_8
X_18457_ _35728_/Q _35088_/Q _34448_/Q _33808_/Q _18349_/X _18351_/X VGND VGND VPWR
+ VPWR _18457_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_190 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17408_ _17901_/A VGND VGND VPWR VPWR _17408_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_166_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33454_ _34033_/CLK _33454_/D VGND VGND VPWR VPWR _33454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18388_ _20012_/A VGND VGND VPWR VPWR _18388_/X sky130_fd_sc_hd__buf_6
X_30666_ _30666_/A VGND VGND VPWR VPWR _35564_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32405_ _36196_/CLK _32405_/D VGND VGND VPWR VPWR _32405_/Q sky130_fd_sc_hd__dfxtp_1
X_36173_ _36173_/CLK _36173_/D VGND VGND VPWR VPWR _36173_/Q sky130_fd_sc_hd__dfxtp_1
X_17339_ _33266_/Q _36146_/Q _33138_/Q _33074_/Q _17058_/X _17059_/X VGND VGND VPWR
+ VPWR _17339_/X sky130_fd_sc_hd__mux4_1
XFILLER_186_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33385_ _33512_/CLK _33385_/D VGND VGND VPWR VPWR _33385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30597_ _30597_/A VGND VGND VPWR VPWR _35532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35124_ _35700_/CLK _35124_/D VGND VGND VPWR VPWR _35124_/Q sky130_fd_sc_hd__dfxtp_1
X_20350_ _35782_/Q _35142_/Q _34502_/Q _33862_/Q _20146_/X _20147_/X VGND VGND VPWR
+ VPWR _20350_/X sky130_fd_sc_hd__mux4_1
X_32336_ _36049_/CLK _32336_/D VGND VGND VPWR VPWR _32336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_918 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19009_ _19002_/X _19004_/X _19007_/X _19008_/X VGND VGND VPWR VPWR _19009_/X sky130_fd_sc_hd__a22o_1
X_35055_ _35953_/CLK _35055_/D VGND VGND VPWR VPWR _35055_/Q sky130_fd_sc_hd__dfxtp_1
X_32267_ _35273_/CLK _32267_/D VGND VGND VPWR VPWR _32267_/Q sky130_fd_sc_hd__dfxtp_1
X_20281_ _20061_/X _20279_/X _20280_/X _20067_/X VGND VGND VPWR VPWR _20281_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34006_ _34006_/CLK _34006_/D VGND VGND VPWR VPWR _34006_/Q sky130_fd_sc_hd__dfxtp_1
X_22020_ _22511_/A VGND VGND VPWR VPWR _22020_/X sky130_fd_sc_hd__clkbuf_4
X_31218_ _31218_/A VGND VGND VPWR VPWR _35826_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32198_ _35885_/CLK _32198_/D VGND VGND VPWR VPWR _32198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31149_ _31149_/A VGND VGND VPWR VPWR _35793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23971_ _23971_/A VGND VGND VPWR VPWR _32525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35957_ _35958_/CLK _35957_/D VGND VGND VPWR VPWR _35957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_284_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _32954_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25710_ _25710_/A VGND VGND VPWR VPWR _33280_/D sky130_fd_sc_hd__clkbuf_1
X_22922_ _22922_/A VGND VGND VPWR VPWR _32027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26690_ _33743_/Q _24249_/X _26706_/S VGND VGND VPWR VPWR _26691_/A sky130_fd_sc_hd__mux2_1
X_34908_ _35036_/CLK _34908_/D VGND VGND VPWR VPWR _34908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35888_ _35952_/CLK _35888_/D VGND VGND VPWR VPWR _35888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22853_ _33293_/Q _36173_/Q _33165_/Q _33101_/Q _20628_/X _21757_/A VGND VGND VPWR
+ VPWR _22853_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25641_ _33248_/Q _24301_/X _25643_/S VGND VGND VPWR VPWR _25642_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34839_ _34967_/CLK _34839_/D VGND VGND VPWR VPWR _34839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21804_ _34030_/Q _33966_/Q _33902_/Q _32238_/Q _21620_/X _21621_/X VGND VGND VPWR
+ VPWR _21804_/X sky130_fd_sc_hd__mux4_1
X_28360_ _28360_/A VGND VGND VPWR VPWR _34503_/D sky130_fd_sc_hd__clkbuf_1
X_25572_ _25572_/A VGND VGND VPWR VPWR _33216_/D sky130_fd_sc_hd__clkbuf_1
X_22784_ _22784_/A VGND VGND VPWR VPWR _36234_/D sky130_fd_sc_hd__clkbuf_1
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27311_ _34007_/Q _24273_/X _27311_/S VGND VGND VPWR VPWR _27312_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24523_ _22994_/X _32755_/Q _24527_/S VGND VGND VPWR VPWR _24524_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21735_ _21663_/X _21733_/X _21734_/X _21667_/X VGND VGND VPWR VPWR _21735_/X sky130_fd_sc_hd__a22o_1
XFILLER_243_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28291_ _28291_/A VGND VGND VPWR VPWR _34470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24454_ _22892_/X _32722_/Q _24464_/S VGND VGND VPWR VPWR _24455_/A sky130_fd_sc_hd__mux2_1
X_27242_ _26946_/X _33974_/Q _27260_/S VGND VGND VPWR VPWR _27243_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21666_ _33002_/Q _32938_/Q _32874_/Q _32810_/Q _21589_/X _21590_/X VGND VGND VPWR
+ VPWR _21666_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23405_ _32261_/Q _23319_/X _23413_/S VGND VGND VPWR VPWR _23406_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27173_ _27173_/A VGND VGND VPWR VPWR _33941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20617_ _20659_/A VGND VGND VPWR VPWR _22362_/A sky130_fd_sc_hd__buf_12
X_24385_ input40/X VGND VGND VPWR VPWR _24385_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_71_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21597_ _22458_/A VGND VGND VPWR VPWR _21597_/X sky130_fd_sc_hd__buf_4
X_26124_ _25159_/X _33476_/Q _26134_/S VGND VGND VPWR VPWR _26125_/A sky130_fd_sc_hd__mux2_1
X_23336_ input57/X VGND VGND VPWR VPWR _23336_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_197_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20548_ _33549_/Q _33485_/Q _33421_/Q _33357_/Q _18333_/X _18335_/X VGND VGND VPWR
+ VPWR _20548_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26055_ _25057_/X _33443_/Q _26071_/S VGND VGND VPWR VPWR _26056_/A sky130_fd_sc_hd__mux2_1
X_23267_ input33/X VGND VGND VPWR VPWR _23267_/X sky130_fd_sc_hd__clkbuf_4
X_20479_ _34570_/Q _32458_/Q _34442_/Q _34378_/Q _20231_/X _20232_/X VGND VGND VPWR
+ VPWR _20479_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25006_ _25006_/A VGND VGND VPWR VPWR _32978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22218_ _33786_/Q _33722_/Q _33658_/Q _33594_/Q _22149_/X _22150_/X VGND VGND VPWR
+ VPWR _22218_/X sky130_fd_sc_hd__mux4_1
XFILLER_234_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23198_ _23198_/A VGND VGND VPWR VPWR _32181_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29814_ _35161_/Q _29086_/X _29830_/S VGND VGND VPWR VPWR _29815_/A sky130_fd_sc_hd__mux2_1
XTAP_6733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22149_ _22502_/A VGND VGND VPWR VPWR _22149_/X sky130_fd_sc_hd__buf_4
XTAP_6744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29745_ _29745_/A VGND VGND VPWR VPWR _35128_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26957_ _26956_/X _33849_/Q _26975_/S VGND VGND VPWR VPWR _26958_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_275_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _33723_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_86_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16710_ _17908_/A VGND VGND VPWR VPWR _16710_/X sky130_fd_sc_hd__clkbuf_4
X_25908_ _25908_/A VGND VGND VPWR VPWR _33373_/D sky130_fd_sc_hd__clkbuf_1
X_17690_ _17686_/X _17689_/X _17481_/X VGND VGND VPWR VPWR _17720_/A sky130_fd_sc_hd__o21ba_1
X_29676_ _29787_/S VGND VGND VPWR VPWR _29695_/S sky130_fd_sc_hd__buf_4
X_26888_ input14/X VGND VGND VPWR VPWR _26888_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28627_ _26996_/X _34630_/Q _28633_/S VGND VGND VPWR VPWR _28628_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16641_ _17855_/A VGND VGND VPWR VPWR _16641_/X sky130_fd_sc_hd__buf_4
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25839_ _25137_/X _33341_/Q _25843_/S VGND VGND VPWR VPWR _25840_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19360_ _33258_/Q _36138_/Q _33130_/Q _33066_/Q _19358_/X _19359_/X VGND VGND VPWR
+ VPWR _19360_/X sky130_fd_sc_hd__mux4_1
X_28558_ _26894_/X _34597_/Q _28570_/S VGND VGND VPWR VPWR _28559_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16572_ _32988_/Q _32924_/Q _32860_/Q _32796_/Q _16283_/X _16284_/X VGND VGND VPWR
+ VPWR _16572_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18311_ _20134_/A VGND VGND VPWR VPWR _18311_/X sky130_fd_sc_hd__buf_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27509_ _26943_/X _34101_/Q _27509_/S VGND VGND VPWR VPWR _27510_/A sky130_fd_sc_hd__mux2_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19291_ _33000_/Q _32936_/Q _32872_/Q _32808_/Q _19289_/X _19290_/X VGND VGND VPWR
+ VPWR _19291_/X sky130_fd_sc_hd__mux4_1
X_28489_ _28489_/A VGND VGND VPWR VPWR _34564_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18242_ _18238_/X _18241_/X _17867_/A VGND VGND VPWR VPWR _18243_/D sky130_fd_sc_hd__o21ba_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30520_ _30520_/A VGND VGND VPWR VPWR _35495_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18173_ _33226_/Q _32586_/Q _35978_/Q _35914_/Q _16075_/X _16076_/X VGND VGND VPWR
+ VPWR _18173_/X sky130_fd_sc_hd__mux4_1
X_30451_ _23327_/X _35463_/Q _30455_/S VGND VGND VPWR VPWR _30452_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17124_ _17830_/A VGND VGND VPWR VPWR _17124_/X sky130_fd_sc_hd__buf_4
XFILLER_190_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33170_ _36114_/CLK _33170_/D VGND VGND VPWR VPWR _33170_/Q sky130_fd_sc_hd__dfxtp_1
X_30382_ _23217_/X _35430_/Q _30392_/S VGND VGND VPWR VPWR _30383_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32121_ _35950_/CLK _32121_/D VGND VGND VPWR VPWR _32121_/Q sky130_fd_sc_hd__dfxtp_2
X_17055_ _17901_/A VGND VGND VPWR VPWR _17055_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_143_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16006_ _16059_/A VGND VGND VPWR VPWR _17957_/A sky130_fd_sc_hd__buf_12
XFILLER_143_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32052_ _33013_/CLK _32052_/D VGND VGND VPWR VPWR _32052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31003_ _35725_/Q _29246_/X _31003_/S VGND VGND VPWR VPWR _31004_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35811_ _35811_/CLK _35811_/D VGND VGND VPWR VPWR _35811_/Q sky130_fd_sc_hd__dfxtp_1
X_17957_ _17957_/A VGND VGND VPWR VPWR _17957_/X sky130_fd_sc_hd__buf_4
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_266_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _36161_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_239_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35742_ _35935_/CLK _35742_/D VGND VGND VPWR VPWR _35742_/Q sky130_fd_sc_hd__dfxtp_1
X_16908_ _16801_/X _16906_/X _16907_/X _16806_/X VGND VGND VPWR VPWR _16908_/X sky130_fd_sc_hd__a22o_1
X_32954_ _32954_/CLK _32954_/D VGND VGND VPWR VPWR _32954_/Q sky130_fd_sc_hd__dfxtp_1
X_17888_ _35585_/Q _35521_/Q _35457_/Q _35393_/Q _17603_/X _17604_/X VGND VGND VPWR
+ VPWR _17888_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31905_ _23277_/X _36152_/Q _31919_/S VGND VGND VPWR VPWR _31906_/A sky130_fd_sc_hd__mux2_1
X_19627_ _19454_/X _19625_/X _19626_/X _19459_/X VGND VGND VPWR VPWR _19627_/X sky130_fd_sc_hd__a22o_1
X_16839_ _16835_/X _16838_/X _16808_/X VGND VGND VPWR VPWR _16840_/D sky130_fd_sc_hd__o21ba_1
X_35673_ _36063_/CLK _35673_/D VGND VGND VPWR VPWR _35673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32885_ _35829_/CLK _32885_/D VGND VGND VPWR VPWR _32885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34624_ _35328_/CLK _34624_/D VGND VGND VPWR VPWR _34624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1063 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31836_ _31836_/A VGND VGND VPWR VPWR _36119_/D sky130_fd_sc_hd__clkbuf_1
X_19558_ _19449_/X _19556_/X _19557_/X _19452_/X VGND VGND VPWR VPWR _19558_/X sky130_fd_sc_hd__a22o_1
X_18509_ _33490_/Q _33426_/Q _33362_/Q _33298_/Q _18298_/X _18299_/X VGND VGND VPWR
+ VPWR _18509_/X sky130_fd_sc_hd__mux4_1
XFILLER_206_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34555_ _34620_/CLK _34555_/D VGND VGND VPWR VPWR _34555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19489_ _34541_/Q _32429_/Q _34413_/Q _34349_/Q _19172_/X _19173_/X VGND VGND VPWR
+ VPWR _19489_/X sky130_fd_sc_hd__mux4_1
X_31767_ _31767_/A VGND VGND VPWR VPWR _36086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33506_ _34276_/CLK _33506_/D VGND VGND VPWR VPWR _33506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21520_ _32742_/Q _32678_/Q _32614_/Q _36070_/Q _21519_/X _21303_/X VGND VGND VPWR
+ VPWR _21520_/X sky130_fd_sc_hd__mux4_1
X_30718_ _30718_/A VGND VGND VPWR VPWR _35589_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34486_ _34809_/CLK _34486_/D VGND VGND VPWR VPWR _34486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_947 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31698_ _36054_/Q input63/X _31700_/S VGND VGND VPWR VPWR _31699_/A sky130_fd_sc_hd__mux2_1
X_36225_ _36228_/CLK _36225_/D VGND VGND VPWR VPWR _36225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21451_ _34020_/Q _33956_/Q _33892_/Q _32171_/Q _21267_/X _21268_/X VGND VGND VPWR
+ VPWR _21451_/X sky130_fd_sc_hd__mux4_1
X_33437_ _33946_/CLK _33437_/D VGND VGND VPWR VPWR _33437_/Q sky130_fd_sc_hd__dfxtp_1
X_30649_ _30649_/A VGND VGND VPWR VPWR _35556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20402_ _32776_/Q _32712_/Q _32648_/Q _36104_/Q _20278_/X _19173_/A VGND VGND VPWR
+ VPWR _20402_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36156_ _36156_/CLK _36156_/D VGND VGND VPWR VPWR _36156_/Q sky130_fd_sc_hd__dfxtp_1
X_24170_ _24170_/A VGND VGND VPWR VPWR _32618_/D sky130_fd_sc_hd__clkbuf_1
X_33368_ _36185_/CLK _33368_/D VGND VGND VPWR VPWR _33368_/Q sky130_fd_sc_hd__dfxtp_1
X_21382_ _21310_/X _21380_/X _21381_/X _21314_/X VGND VGND VPWR VPWR _21382_/X sky130_fd_sc_hd__a22o_1
XFILLER_200_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35107_ _35748_/CLK _35107_/D VGND VGND VPWR VPWR _35107_/Q sky130_fd_sc_hd__dfxtp_1
X_23121_ input3/X VGND VGND VPWR VPWR _23121_/X sky130_fd_sc_hd__buf_6
X_20333_ _20333_/A _20333_/B _20333_/C _20333_/D VGND VGND VPWR VPWR _20334_/A sky130_fd_sc_hd__or4_2
X_32319_ _35966_/CLK _32319_/D VGND VGND VPWR VPWR _32319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36087_ _36087_/CLK _36087_/D VGND VGND VPWR VPWR _36087_/Q sky130_fd_sc_hd__dfxtp_1
X_33299_ _36237_/CLK _33299_/D VGND VGND VPWR VPWR _33299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23052_ _23052_/A VGND VGND VPWR VPWR _32069_/D sky130_fd_sc_hd__clkbuf_1
X_35038_ _35038_/CLK _35038_/D VGND VGND VPWR VPWR _35038_/Q sky130_fd_sc_hd__dfxtp_1
X_20264_ _20155_/X _20262_/X _20263_/X _20158_/X VGND VGND VPWR VPWR _20264_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22003_ _21795_/X _22001_/X _22002_/X _21800_/X VGND VGND VPWR VPWR _22003_/X sky130_fd_sc_hd__a22o_1
XTAP_6029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27860_ _34266_/Q _24283_/X _27874_/S VGND VGND VPWR VPWR _27861_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20195_ _34561_/Q _32449_/Q _34433_/Q _34369_/Q _19878_/X _19879_/X VGND VGND VPWR
+ VPWR _20195_/X sky130_fd_sc_hd__mux4_1
XTAP_5306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26811_ _33801_/Q _24428_/X _26811_/S VGND VGND VPWR VPWR _26812_/A sky130_fd_sc_hd__mux2_1
XTAP_5328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27791_ _27791_/A VGND VGND VPWR VPWR _34233_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_257_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _36167_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29530_ _29530_/A VGND VGND VPWR VPWR _35026_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26742_ _33768_/Q _24326_/X _26748_/S VGND VGND VPWR VPWR _26743_/A sky130_fd_sc_hd__mux2_1
X_23954_ _23050_/X _32517_/Q _23962_/S VGND VGND VPWR VPWR _23955_/A sky130_fd_sc_hd__mux2_1
XTAP_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22905_ _22904_/X _32022_/Q _22908_/S VGND VGND VPWR VPWR _22906_/A sky130_fd_sc_hd__mux2_1
XTAP_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29461_ _23256_/X _34994_/Q _29467_/S VGND VGND VPWR VPWR _29462_/A sky130_fd_sc_hd__mux2_1
X_26673_ _25171_/X _33736_/Q _26675_/S VGND VGND VPWR VPWR _26674_/A sky130_fd_sc_hd__mux2_1
X_23885_ _22948_/X _32484_/Q _23899_/S VGND VGND VPWR VPWR _23886_/A sky130_fd_sc_hd__mux2_1
XANTENNA_904 _26412_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_915 _26968_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28412_ _26878_/X _34528_/Q _28414_/S VGND VGND VPWR VPWR _28413_/A sky130_fd_sc_hd__mux2_1
X_22836_ _34828_/Q _34764_/Q _34700_/Q _34636_/Q _22594_/X _22595_/X VGND VGND VPWR
+ VPWR _22836_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25624_ _25735_/S VGND VGND VPWR VPWR _25643_/S sky130_fd_sc_hd__buf_6
XANTENNA_926 _27781_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29392_ _23096_/X _34961_/Q _29404_/S VGND VGND VPWR VPWR _29393_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_937 _29070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_948 _29517_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_959 _29922_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28343_ _28343_/A VGND VGND VPWR VPWR _34495_/D sky130_fd_sc_hd__clkbuf_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22767_ _21754_/A _22765_/X _22766_/X _21759_/A VGND VGND VPWR VPWR _22767_/X sky130_fd_sc_hd__a22o_1
X_25555_ _25555_/A VGND VGND VPWR VPWR _33208_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21718_ _21718_/A _21718_/B _21718_/C _21718_/D VGND VGND VPWR VPWR _21719_/A sky130_fd_sc_hd__or4_4
X_24506_ _22969_/X _32747_/Q _24506_/S VGND VGND VPWR VPWR _24507_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28274_ _28274_/A VGND VGND VPWR VPWR _34462_/D sky130_fd_sc_hd__clkbuf_1
X_25486_ _25597_/S VGND VGND VPWR VPWR _25505_/S sky130_fd_sc_hd__buf_4
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22698_ _33544_/Q _33480_/Q _33416_/Q _33352_/Q _22429_/X _22430_/X VGND VGND VPWR
+ VPWR _22698_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1070 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27225_ _26922_/X _33966_/Q _27239_/S VGND VGND VPWR VPWR _27226_/A sky130_fd_sc_hd__mux2_1
X_24437_ input59/X VGND VGND VPWR VPWR _24437_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_205_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21649_ _34282_/Q _34218_/Q _34154_/Q _34090_/Q _21336_/X _21337_/X VGND VGND VPWR
+ VPWR _21649_/X sky130_fd_sc_hd__mux4_1
XFILLER_199_1439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27156_ _27426_/A _30465_/B VGND VGND VPWR VPWR _27289_/S sky130_fd_sc_hd__nand2_8
X_24368_ _24368_/A VGND VGND VPWR VPWR _32693_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_90 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23319_ input51/X VGND VGND VPWR VPWR _23319_/X sky130_fd_sc_hd__buf_4
X_26107_ _25134_/X _33468_/Q _26113_/S VGND VGND VPWR VPWR _26108_/A sky130_fd_sc_hd__mux2_1
X_27087_ _27087_/A VGND VGND VPWR VPWR _33900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24299_ _32671_/Q _24298_/X _24305_/S VGND VGND VPWR VPWR _24300_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26038_ _25032_/X _33435_/Q _26050_/S VGND VGND VPWR VPWR _26039_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_496_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _34973_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_234_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1303 _16557_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18860_ _34268_/Q _34204_/Q _34140_/Q _34076_/Q _18683_/X _18684_/X VGND VGND VPWR
+ VPWR _18860_/X sky130_fd_sc_hd__mux4_1
XTAP_6530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1314 _32121_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1325 _20256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1336 _19454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17811_ _35775_/Q _35135_/Q _34495_/Q _33855_/Q _17493_/X _17494_/X VGND VGND VPWR
+ VPWR _17811_/X sky130_fd_sc_hd__mux4_1
XTAP_6563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1347 _22446_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1358 _22904_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18791_ _20203_/A VGND VGND VPWR VPWR _18791_/X sky130_fd_sc_hd__buf_4
XTAP_6585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1369 _24407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27989_ _27989_/A VGND VGND VPWR VPWR _34327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_248_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _34306_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_5851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17742_ _33213_/Q _32573_/Q _35965_/Q _35901_/Q _17427_/X _17428_/X VGND VGND VPWR
+ VPWR _17742_/X sky130_fd_sc_hd__mux4_1
X_29728_ _29728_/A VGND VGND VPWR VPWR _35120_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29659_ _29659_/A VGND VGND VPWR VPWR _35087_/D sky130_fd_sc_hd__clkbuf_1
X_17673_ _17352_/X _17671_/X _17672_/X _17355_/X VGND VGND VPWR VPWR _17673_/X sky130_fd_sc_hd__a22o_1
XFILLER_35_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19412_ _35307_/Q _35243_/Q _35179_/Q _32299_/Q _19306_/X _19307_/X VGND VGND VPWR
+ VPWR _19412_/X sky130_fd_sc_hd__mux4_1
X_16624_ _16624_/A VGND VGND VPWR VPWR _31965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32670_ _34271_/CLK _32670_/D VGND VGND VPWR VPWR _32670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31621_ _31621_/A VGND VGND VPWR VPWR _36017_/D sky130_fd_sc_hd__clkbuf_1
X_19343_ _35049_/Q _34985_/Q _34921_/Q _34857_/Q _19103_/X _19104_/X VGND VGND VPWR
+ VPWR _19343_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16555_ _16448_/X _16553_/X _16554_/X _16453_/X VGND VGND VPWR VPWR _16555_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_420_CLK clkbuf_6_38__f_CLK/X VGND VGND VPWR VPWR _35250_/CLK sky130_fd_sc_hd__clkbuf_16
X_34340_ _35300_/CLK _34340_/D VGND VGND VPWR VPWR _34340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31552_ _31552_/A VGND VGND VPWR VPWR _35984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19274_ _19101_/X _19272_/X _19273_/X _19106_/X VGND VGND VPWR VPWR _19274_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16486_ _16482_/X _16485_/X _16455_/X VGND VGND VPWR VPWR _16487_/D sky130_fd_sc_hd__o21ba_1
X_18225_ _32524_/Q _32396_/Q _32076_/Q _36044_/Q _17982_/X _17007_/A VGND VGND VPWR
+ VPWR _18225_/X sky130_fd_sc_hd__mux4_1
X_30503_ _30503_/A VGND VGND VPWR VPWR _35487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34271_ _34271_/CLK _34271_/D VGND VGND VPWR VPWR _34271_/Q sky130_fd_sc_hd__dfxtp_1
X_31483_ _23250_/X _35952_/Q _31493_/S VGND VGND VPWR VPWR _31484_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36010_ _36075_/CLK _36010_/D VGND VGND VPWR VPWR _36010_/Q sky130_fd_sc_hd__dfxtp_1
X_33222_ _35975_/CLK _33222_/D VGND VGND VPWR VPWR _33222_/Q sky130_fd_sc_hd__dfxtp_1
X_18156_ _34314_/Q _34250_/Q _34186_/Q _34122_/Q _16045_/X _16046_/X VGND VGND VPWR
+ VPWR _18156_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30434_ _23300_/X _35455_/Q _30434_/S VGND VGND VPWR VPWR _30435_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_1162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17107_ _35563_/Q _35499_/Q _35435_/Q _35371_/Q _16897_/X _16898_/X VGND VGND VPWR
+ VPWR _17107_/X sky130_fd_sc_hd__mux4_1
X_33153_ _36159_/CLK _33153_/D VGND VGND VPWR VPWR _33153_/Q sky130_fd_sc_hd__dfxtp_1
X_18087_ _35335_/Q _35271_/Q _35207_/Q _32327_/Q _16088_/X _16090_/X VGND VGND VPWR
+ VPWR _18087_/X sky130_fd_sc_hd__mux4_1
X_30365_ _23136_/X _35422_/Q _30371_/S VGND VGND VPWR VPWR _30366_/A sky130_fd_sc_hd__mux2_1
X_32104_ _35808_/CLK _32104_/D VGND VGND VPWR VPWR _32104_/Q sky130_fd_sc_hd__dfxtp_1
X_17038_ _17034_/X _17037_/X _16794_/X VGND VGND VPWR VPWR _17046_/C sky130_fd_sc_hd__o21ba_1
X_33084_ _36156_/CLK _33084_/D VGND VGND VPWR VPWR _33084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30296_ _35390_/Q _29200_/X _30298_/S VGND VGND VPWR VPWR _30297_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_487_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _35744_/CLK sky130_fd_sc_hd__clkbuf_16
X_32035_ _36003_/CLK _32035_/D VGND VGND VPWR VPWR _32035_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_46__f_CLK clkbuf_5_23_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_46__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_113_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ _34527_/Q _32415_/Q _34399_/Q _34335_/Q _18819_/X _18820_/X VGND VGND VPWR
+ VPWR _18989_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_239_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _34819_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_112_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33986_ _34053_/CLK _33986_/D VGND VGND VPWR VPWR _33986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35725_ _35789_/CLK _35725_/D VGND VGND VPWR VPWR _35725_/Q sky130_fd_sc_hd__dfxtp_1
X_20951_ _32726_/Q _32662_/Q _32598_/Q _36054_/Q _20813_/X _20950_/X VGND VGND VPWR
+ VPWR _20951_/X sky130_fd_sc_hd__mux4_1
X_32937_ _36075_/CLK _32937_/D VGND VGND VPWR VPWR _32937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_836 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23670_ _32384_/Q _23303_/X _23688_/S VGND VGND VPWR VPWR _23671_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35656_ _35848_/CLK _35656_/D VGND VGND VPWR VPWR _35656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20882_ _32468_/Q _32340_/Q _32020_/Q _35988_/Q _20817_/X _22463_/A VGND VGND VPWR
+ VPWR _20882_/X sky130_fd_sc_hd__mux4_1
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32868_ _32994_/CLK _32868_/D VGND VGND VPWR VPWR _32868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22621_ _22300_/X _22619_/X _22620_/X _22303_/X VGND VGND VPWR VPWR _22621_/X sky130_fd_sc_hd__a22o_1
X_31819_ _23090_/X _36111_/Q _31835_/S VGND VGND VPWR VPWR _31820_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34607_ _35242_/CLK _34607_/D VGND VGND VPWR VPWR _34607_/Q sky130_fd_sc_hd__dfxtp_1
X_35587_ _35973_/CLK _35587_/D VGND VGND VPWR VPWR _35587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32799_ _35481_/CLK _32799_/D VGND VGND VPWR VPWR _32799_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_411_CLK clkbuf_6_33__f_CLK/X VGND VGND VPWR VPWR _34794_/CLK sky130_fd_sc_hd__clkbuf_16
X_25340_ _25340_/A VGND VGND VPWR VPWR _33108_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22552_ _22548_/X _22551_/X _22442_/X _22443_/X VGND VGND VPWR VPWR _22569_/B sky130_fd_sc_hd__o211a_1
X_34538_ _35179_/CLK _34538_/D VGND VGND VPWR VPWR _34538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21503_ _34789_/Q _34725_/Q _34661_/Q _34597_/Q _21182_/X _21183_/X VGND VGND VPWR
+ VPWR _21503_/X sky130_fd_sc_hd__mux4_1
XFILLER_210_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25271_ _25271_/A VGND VGND VPWR VPWR _33076_/D sky130_fd_sc_hd__clkbuf_1
X_22483_ _22369_/X _22481_/X _22482_/X _22373_/X VGND VGND VPWR VPWR _22483_/X sky130_fd_sc_hd__a22o_1
X_34469_ _35941_/CLK _34469_/D VGND VGND VPWR VPWR _34469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27010_ _27010_/A VGND VGND VPWR VPWR _33866_/D sky130_fd_sc_hd__clkbuf_1
X_24222_ _23044_/X _32643_/Q _24234_/S VGND VGND VPWR VPWR _24223_/A sky130_fd_sc_hd__mux2_1
X_36208_ _36211_/CLK _36208_/D VGND VGND VPWR VPWR _36208_/Q sky130_fd_sc_hd__dfxtp_1
X_21434_ _35299_/Q _35235_/Q _35171_/Q _32291_/Q _21253_/X _21254_/X VGND VGND VPWR
+ VPWR _21434_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24153_ _22941_/X _32610_/Q _24171_/S VGND VGND VPWR VPWR _24154_/A sky130_fd_sc_hd__mux2_1
X_36139_ _36139_/CLK _36139_/D VGND VGND VPWR VPWR _36139_/Q sky130_fd_sc_hd__dfxtp_1
X_21365_ _21365_/A _21365_/B _21365_/C _21365_/D VGND VGND VPWR VPWR _21366_/A sky130_fd_sc_hd__or4_2
XFILLER_206_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23104_ _23104_/A VGND VGND VPWR VPWR _32147_/D sky130_fd_sc_hd__clkbuf_1
X_20316_ _33029_/Q _32965_/Q _32901_/Q _32837_/Q _19995_/X _19996_/X VGND VGND VPWR
+ VPWR _20316_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24084_ _23041_/X _32578_/Q _24098_/S VGND VGND VPWR VPWR _24085_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28961_ _34788_/Q _24314_/X _28975_/S VGND VGND VPWR VPWR _28962_/A sky130_fd_sc_hd__mux2_1
X_21296_ _34272_/Q _34208_/Q _34144_/Q _34080_/Q _20983_/X _20984_/X VGND VGND VPWR
+ VPWR _21296_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_478_CLK clkbuf_6_9__f_CLK/X VGND VGND VPWR VPWR _35932_/CLK sky130_fd_sc_hd__clkbuf_16
X_23035_ _23075_/S VGND VGND VPWR VPWR _23063_/S sky130_fd_sc_hd__clkbuf_8
X_27912_ _34291_/Q _24360_/X _27916_/S VGND VGND VPWR VPWR _27913_/A sky130_fd_sc_hd__mux2_1
X_20247_ _33283_/Q _36163_/Q _33155_/Q _33091_/Q _20064_/X _20065_/X VGND VGND VPWR
+ VPWR _20247_/X sky130_fd_sc_hd__mux4_1
X_28892_ _28892_/A VGND VGND VPWR VPWR _34755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_1071 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27843_ _34258_/Q _24258_/X _27853_/S VGND VGND VPWR VPWR _27844_/A sky130_fd_sc_hd__mux2_1
XTAP_5125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20178_ _32769_/Q _32705_/Q _32641_/Q _36097_/Q _19925_/X _20062_/X VGND VGND VPWR
+ VPWR _20178_/X sky130_fd_sc_hd__mux4_1
XTAP_5136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27774_ _27774_/A VGND VGND VPWR VPWR _34225_/D sky130_fd_sc_hd__clkbuf_1
X_24986_ _24986_/A VGND VGND VPWR VPWR _32972_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29513_ _23339_/X _35019_/Q _29517_/S VGND VGND VPWR VPWR _29514_/A sky130_fd_sc_hd__mux2_1
XTAP_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26725_ _33760_/Q _24301_/X _26727_/S VGND VGND VPWR VPWR _26726_/A sky130_fd_sc_hd__mux2_1
X_23937_ _23025_/X _32509_/Q _23941_/S VGND VGND VPWR VPWR _23938_/A sky130_fd_sc_hd__mux2_1
XTAP_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_701 _22458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_712 _22465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29444_ _23231_/X _34986_/Q _29446_/S VGND VGND VPWR VPWR _29445_/A sky130_fd_sc_hd__mux2_1
XFILLER_233_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26656_ _26683_/S VGND VGND VPWR VPWR _26675_/S sky130_fd_sc_hd__buf_6
XANTENNA_723 _21759_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_734 _21223_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23868_ _22923_/X _32476_/Q _23878_/S VGND VGND VPWR VPWR _23869_/A sky130_fd_sc_hd__mux2_1
XANTENNA_745 _22217_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_756 _22470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25607_ _25607_/A VGND VGND VPWR VPWR _33231_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29375_ _29375_/A VGND VGND VPWR VPWR _34953_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_767 _22538_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22819_ _34060_/Q _33996_/Q _33932_/Q _32268_/Q _20658_/X _20660_/X VGND VGND VPWR
+ VPWR _22819_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_778 _22604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26587_ _25044_/X _33695_/Q _26591_/S VGND VGND VPWR VPWR _26588_/A sky130_fd_sc_hd__mux2_1
XANTENNA_789 _22664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23799_ _23022_/X _32444_/Q _23805_/S VGND VGND VPWR VPWR _23800_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_402_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _35819_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_241_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16340_ _16340_/A _16340_/B _16340_/C _16340_/D VGND VGND VPWR VPWR _16341_/A sky130_fd_sc_hd__or4_4
X_28326_ _34487_/Q _24373_/X _28342_/S VGND VGND VPWR VPWR _28327_/A sky130_fd_sc_hd__mux2_1
X_25538_ _25538_/A VGND VGND VPWR VPWR _33200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28257_ _28257_/A VGND VGND VPWR VPWR _34454_/D sky130_fd_sc_hd__clkbuf_1
X_16271_ _16271_/A VGND VGND VPWR VPWR _31955_/D sky130_fd_sc_hd__clkbuf_1
X_25469_ _25469_/A VGND VGND VPWR VPWR _33167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18010_ _17908_/X _18008_/X _18009_/X _17911_/X VGND VGND VPWR VPWR _18010_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27208_ _26897_/X _33958_/Q _27218_/S VGND VGND VPWR VPWR _27209_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_1192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28188_ _28236_/S VGND VGND VPWR VPWR _28207_/S sky130_fd_sc_hd__buf_4
XFILLER_218_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27139_ _27139_/A VGND VGND VPWR VPWR _33925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19961_ _19708_/X _19959_/X _19960_/X _19714_/X VGND VGND VPWR VPWR _19961_/X sky130_fd_sc_hd__a22o_1
X_30150_ _30150_/A VGND VGND VPWR VPWR _35320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_469_CLK clkbuf_6_8__f_CLK/X VGND VGND VPWR VPWR _35748_/CLK sky130_fd_sc_hd__clkbuf_16
X_18912_ _35549_/Q _35485_/Q _35421_/Q _35357_/Q _18844_/X _18845_/X VGND VGND VPWR
+ VPWR _18912_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19892_ _19888_/X _19891_/X _19781_/X VGND VGND VPWR VPWR _19916_/A sky130_fd_sc_hd__o21ba_1
XANTENNA_1100 _17368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30081_ _30192_/S VGND VGND VPWR VPWR _30100_/S sky130_fd_sc_hd__buf_4
XTAP_7061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1111 _32123_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1122 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1133 _17911_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18843_ _18588_/X _18841_/X _18842_/X _18591_/X VGND VGND VPWR VPWR _18843_/X sky130_fd_sc_hd__a22o_1
XFILLER_67_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1144 _20165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1155 _22503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1166 _22443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1177 _20908_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33840_ _35760_/CLK _33840_/D VGND VGND VPWR VPWR _33840_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1188 _22506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18774_ _35737_/Q _35097_/Q _34457_/Q _33817_/Q _18734_/X _18735_/X VGND VGND VPWR
+ VPWR _18774_/X sky130_fd_sc_hd__mux4_1
XTAP_5670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15986_ _17767_/A VGND VGND VPWR VPWR _17906_/A sky130_fd_sc_hd__buf_12
XANTENNA_1199 _23077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17725_ _33533_/Q _33469_/Q _33405_/Q _33341_/Q _17476_/X _17477_/X VGND VGND VPWR
+ VPWR _17725_/X sky130_fd_sc_hd__mux4_1
X_33771_ _34281_/CLK _33771_/D VGND VGND VPWR VPWR _33771_/Q sky130_fd_sc_hd__dfxtp_1
X_30983_ _35715_/Q _29216_/X _30995_/S VGND VGND VPWR VPWR _30984_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32722_ _36050_/CLK _32722_/D VGND VGND VPWR VPWR _32722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35510_ _35956_/CLK _35510_/D VGND VGND VPWR VPWR _35510_/Q sky130_fd_sc_hd__dfxtp_1
X_17656_ _34043_/Q _33979_/Q _33915_/Q _32251_/Q _17373_/X _17374_/X VGND VGND VPWR
+ VPWR _17656_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16607_ _17795_/A VGND VGND VPWR VPWR _16607_/X sky130_fd_sc_hd__buf_4
X_35441_ _35953_/CLK _35441_/D VGND VGND VPWR VPWR _35441_/Q sky130_fd_sc_hd__dfxtp_1
X_32653_ _36173_/CLK _32653_/D VGND VGND VPWR VPWR _32653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17587_ _34297_/Q _34233_/Q _34169_/Q _34105_/Q _17442_/X _17443_/X VGND VGND VPWR
+ VPWR _17587_/X sky130_fd_sc_hd__mux4_1
XFILLER_211_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31604_ _31604_/A VGND VGND VPWR VPWR _36009_/D sky130_fd_sc_hd__clkbuf_1
X_19326_ _33257_/Q _36137_/Q _33129_/Q _33065_/Q _19005_/X _19006_/X VGND VGND VPWR
+ VPWR _19326_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16538_ _32987_/Q _32923_/Q _32859_/Q _32795_/Q _16283_/X _16284_/X VGND VGND VPWR
+ VPWR _16538_/X sky130_fd_sc_hd__mux4_1
X_35372_ _35946_/CLK _35372_/D VGND VGND VPWR VPWR _35372_/Q sky130_fd_sc_hd__dfxtp_1
X_32584_ _35977_/CLK _32584_/D VGND VGND VPWR VPWR _32584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34323_ _36204_/CLK _34323_/D VGND VGND VPWR VPWR _34323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31535_ _23333_/X _35977_/Q _31535_/S VGND VGND VPWR VPWR _31536_/A sky130_fd_sc_hd__mux2_1
X_19257_ _32999_/Q _32935_/Q _32871_/Q _32807_/Q _18936_/X _18937_/X VGND VGND VPWR
+ VPWR _19257_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16469_ _32473_/Q _32345_/Q _32025_/Q _35993_/Q _16217_/X _16358_/X VGND VGND VPWR
+ VPWR _16469_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18208_ _16044_/X _18206_/X _18207_/X _16054_/X VGND VGND VPWR VPWR _18208_/X sky130_fd_sc_hd__a22o_1
X_34254_ _34256_/CLK _34254_/D VGND VGND VPWR VPWR _34254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31466_ _23223_/X _35944_/Q _31472_/S VGND VGND VPWR VPWR _31467_/A sky130_fd_sc_hd__mux2_1
X_19188_ _33253_/Q _36133_/Q _33125_/Q _33061_/Q _19005_/X _19006_/X VGND VGND VPWR
+ VPWR _19188_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33205_ _35958_/CLK _33205_/D VGND VGND VPWR VPWR _33205_/Q sky130_fd_sc_hd__dfxtp_1
X_18139_ _35849_/Q _32229_/Q _35721_/Q _35657_/Q _15989_/X _15991_/X VGND VGND VPWR
+ VPWR _18139_/X sky130_fd_sc_hd__mux4_1
X_30417_ _30417_/A VGND VGND VPWR VPWR _35446_/D sky130_fd_sc_hd__clkbuf_1
X_34185_ _34752_/CLK _34185_/D VGND VGND VPWR VPWR _34185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31397_ _31397_/A VGND VGND VPWR VPWR _35911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33136_ _36081_/CLK _33136_/D VGND VGND VPWR VPWR _33136_/Q sky130_fd_sc_hd__dfxtp_1
X_21150_ _34779_/Q _34715_/Q _34651_/Q _34587_/Q _20829_/X _20830_/X VGND VGND VPWR
+ VPWR _21150_/X sky130_fd_sc_hd__mux4_1
XFILLER_171_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30348_ _23111_/X _35414_/Q _30350_/S VGND VGND VPWR VPWR _30349_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20101_ _19855_/X _20099_/X _20100_/X _19858_/X VGND VGND VPWR VPWR _20101_/X sky130_fd_sc_hd__a22o_1
XFILLER_217_1030 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21081_ _35289_/Q _35225_/Q _35161_/Q _32281_/Q _20900_/X _20901_/X VGND VGND VPWR
+ VPWR _21081_/X sky130_fd_sc_hd__mux4_1
X_33067_ _36139_/CLK _33067_/D VGND VGND VPWR VPWR _33067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30279_ _30327_/S VGND VGND VPWR VPWR _30298_/S sky130_fd_sc_hd__buf_6
X_20032_ _33277_/Q _36157_/Q _33149_/Q _33085_/Q _19711_/X _19712_/X VGND VGND VPWR
+ VPWR _20032_/X sky130_fd_sc_hd__mux4_1
X_32018_ _36052_/CLK _32018_/D VGND VGND VPWR VPWR _32018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24840_ _23056_/X _32903_/Q _24844_/S VGND VGND VPWR VPWR _24841_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21983_ _21663_/X _21981_/X _21982_/X _21667_/X VGND VGND VPWR VPWR _21983_/X sky130_fd_sc_hd__a22o_1
X_24771_ _22954_/X _32870_/Q _24781_/S VGND VGND VPWR VPWR _24772_/A sky130_fd_sc_hd__mux2_1
X_33969_ _34222_/CLK _33969_/D VGND VGND VPWR VPWR _33969_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26510_ _25131_/X _33659_/Q _26518_/S VGND VGND VPWR VPWR _26511_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23722_ _23722_/A VGND VGND VPWR VPWR _32407_/D sky130_fd_sc_hd__clkbuf_1
X_35708_ _35772_/CLK _35708_/D VGND VGND VPWR VPWR _35708_/Q sky130_fd_sc_hd__dfxtp_1
X_20934_ _35285_/Q _35221_/Q _35157_/Q _32277_/Q _20900_/X _20901_/X VGND VGND VPWR
+ VPWR _20934_/X sky130_fd_sc_hd__mux4_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27490_ _27559_/S VGND VGND VPWR VPWR _27509_/S sky130_fd_sc_hd__clkbuf_8
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26441_ _25029_/X _33626_/Q _26455_/S VGND VGND VPWR VPWR _26442_/A sky130_fd_sc_hd__mux2_1
X_20865_ _20674_/X _20863_/X _20864_/X _20684_/X VGND VGND VPWR VPWR _20865_/X sky130_fd_sc_hd__a22o_1
X_23653_ _32376_/Q _23277_/X _23667_/S VGND VGND VPWR VPWR _23654_/A sky130_fd_sc_hd__mux2_1
X_35639_ _35831_/CLK _35639_/D VGND VGND VPWR VPWR _35639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22604_ _22604_/A VGND VGND VPWR VPWR _36228_/D sky130_fd_sc_hd__clkbuf_1
X_29160_ input29/X VGND VGND VPWR VPWR _29160_/X sky130_fd_sc_hd__buf_2
X_23584_ _23584_/A VGND VGND VPWR VPWR _32343_/D sky130_fd_sc_hd__clkbuf_1
X_26372_ _26372_/A VGND VGND VPWR VPWR _33593_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20796_ _20790_/X _20795_/X _20671_/X VGND VGND VPWR VPWR _20804_/C sky130_fd_sc_hd__o21ba_1
XFILLER_179_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28111_ _26832_/X _34385_/Q _28123_/S VGND VGND VPWR VPWR _28112_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22535_ _22460_/X _22533_/X _22534_/X _22465_/X VGND VGND VPWR VPWR _22535_/X sky130_fd_sc_hd__a22o_1
X_25323_ _25323_/A VGND VGND VPWR VPWR _33101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29091_ _29091_/A VGND VGND VPWR VPWR _34842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28042_ _28042_/A VGND VGND VPWR VPWR _34352_/D sky130_fd_sc_hd__clkbuf_1
X_22466_ _22460_/X _22461_/X _22464_/X _22465_/X VGND VGND VPWR VPWR _22466_/X sky130_fd_sc_hd__a22o_1
X_25254_ _25084_/X _33068_/Q _25272_/S VGND VGND VPWR VPWR _25255_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24205_ _23019_/X _32635_/Q _24213_/S VGND VGND VPWR VPWR _24206_/A sky130_fd_sc_hd__mux2_1
X_21417_ _21096_/X _21415_/X _21416_/X _21099_/X VGND VGND VPWR VPWR _21417_/X sky130_fd_sc_hd__a22o_1
X_25185_ _25185_/A VGND VGND VPWR VPWR _33036_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22397_ _34303_/Q _34239_/Q _34175_/Q _34111_/Q _22395_/X _22396_/X VGND VGND VPWR
+ VPWR _22397_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24136_ _22917_/X _32602_/Q _24150_/S VGND VGND VPWR VPWR _24137_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21348_ _32993_/Q _32929_/Q _32865_/Q _32801_/Q _21236_/X _21237_/X VGND VGND VPWR
+ VPWR _21348_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29993_ _35246_/Q _29151_/X _30007_/S VGND VGND VPWR VPWR _29994_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24067_ _23016_/X _32570_/Q _24077_/S VGND VGND VPWR VPWR _24068_/A sky130_fd_sc_hd__mux2_1
X_28944_ _34780_/Q _24289_/X _28954_/S VGND VGND VPWR VPWR _28945_/A sky130_fd_sc_hd__mux2_1
X_21279_ _35807_/Q _32183_/Q _35679_/Q _35615_/Q _21207_/X _21208_/X VGND VGND VPWR
+ VPWR _21279_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23018_ _23018_/A VGND VGND VPWR VPWR _32058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28875_ _28875_/A VGND VGND VPWR VPWR _34747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27826_ _27826_/A VGND VGND VPWR VPWR _34250_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27757_ _27757_/A VGND VGND VPWR VPWR _34217_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24969_ _23047_/X _32964_/Q _24979_/S VGND VGND VPWR VPWR _24970_/A sky130_fd_sc_hd__mux2_1
XTAP_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17510_ _17863_/A VGND VGND VPWR VPWR _17510_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26708_ _26819_/S VGND VGND VPWR VPWR _26727_/S sky130_fd_sc_hd__buf_4
XTAP_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18490_ _18344_/X _18488_/X _18489_/X _18354_/X VGND VGND VPWR VPWR _18490_/X sky130_fd_sc_hd__a22o_1
XTAP_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27688_ _34185_/Q _24428_/X _27688_/S VGND VGND VPWR VPWR _27689_/A sky130_fd_sc_hd__mux2_1
XTAP_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_520 _17970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_531 _18214_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_542 _20257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29427_ _29517_/S VGND VGND VPWR VPWR _29446_/S sky130_fd_sc_hd__buf_4
XFILLER_79_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17441_ _33781_/Q _33717_/Q _33653_/Q _33589_/Q _17196_/X _17197_/X VGND VGND VPWR
+ VPWR _17441_/X sky130_fd_sc_hd__mux4_1
XANTENNA_553 _20143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26639_ _26639_/A VGND VGND VPWR VPWR _33719_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_564 _20147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_575 _20165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_586 _19454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29358_ _23307_/X _34945_/Q _29374_/S VGND VGND VPWR VPWR _29359_/A sky130_fd_sc_hd__mux2_1
XANTENNA_597 _20167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17372_ _33523_/Q _33459_/Q _33395_/Q _33331_/Q _17123_/X _17124_/X VGND VGND VPWR
+ VPWR _17372_/X sky130_fd_sc_hd__mux4_1
X_19111_ _19111_/A VGND VGND VPWR VPWR _32098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16323_ _32981_/Q _32917_/Q _32853_/Q _32789_/Q _16283_/X _16284_/X VGND VGND VPWR
+ VPWR _16323_/X sky130_fd_sc_hd__mux4_1
X_28309_ _34479_/Q _24348_/X _28321_/S VGND VGND VPWR VPWR _28310_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29289_ _29289_/A VGND VGND VPWR VPWR _34912_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31320_ _31320_/A VGND VGND VPWR VPWR _35874_/D sky130_fd_sc_hd__clkbuf_1
X_19042_ _18796_/X _19040_/X _19041_/X _18799_/X VGND VGND VPWR VPWR _19042_/X sky130_fd_sc_hd__a22o_1
X_16254_ _17795_/A VGND VGND VPWR VPWR _16254_/X sky130_fd_sc_hd__buf_6
XFILLER_71_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31251_ _35842_/Q input48/X _31265_/S VGND VGND VPWR VPWR _31252_/A sky130_fd_sc_hd__mux2_1
X_16185_ _32977_/Q _32913_/Q _32849_/Q _32785_/Q _16033_/X _16035_/X VGND VGND VPWR
+ VPWR _16185_/X sky130_fd_sc_hd__mux4_1
Xoutput207 _36232_/Q VGND VGND VPWR VPWR D2[58] sky130_fd_sc_hd__buf_2
X_30202_ _35345_/Q _29061_/X _30214_/S VGND VGND VPWR VPWR _30203_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput218 _32078_/Q VGND VGND VPWR VPWR D3[0] sky130_fd_sc_hd__buf_2
XFILLER_182_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput229 _32079_/Q VGND VGND VPWR VPWR D3[1] sky130_fd_sc_hd__buf_2
X_31182_ _31182_/A VGND VGND VPWR VPWR _35809_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30133_ _30133_/A VGND VGND VPWR VPWR _35312_/D sky130_fd_sc_hd__clkbuf_1
X_19944_ _35322_/Q _35258_/Q _35194_/Q _32314_/Q _19659_/X _19660_/X VGND VGND VPWR
+ VPWR _19944_/X sky130_fd_sc_hd__mux4_1
X_35990_ _35991_/CLK _35990_/D VGND VGND VPWR VPWR _35990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30064_ _30064_/A VGND VGND VPWR VPWR _35279_/D sky130_fd_sc_hd__clkbuf_1
X_34941_ _35989_/CLK _34941_/D VGND VGND VPWR VPWR _34941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19875_ _34808_/Q _34744_/Q _34680_/Q _34616_/Q _19588_/X _19589_/X VGND VGND VPWR
+ VPWR _19875_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18826_ _18826_/A VGND VGND VPWR VPWR _32090_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34872_ _35257_/CLK _34872_/D VGND VGND VPWR VPWR _34872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33823_ _35745_/CLK _33823_/D VGND VGND VPWR VPWR _33823_/Q sky130_fd_sc_hd__dfxtp_1
X_18757_ _18757_/A _18757_/B _18757_/C _18757_/D VGND VGND VPWR VPWR _18758_/A sky130_fd_sc_hd__or4_2
XFILLER_97_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17708_ _17865_/A VGND VGND VPWR VPWR _17708_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_224_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33754_ _34266_/CLK _33754_/D VGND VGND VPWR VPWR _33754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18688_ _34007_/Q _33943_/Q _33879_/Q _32151_/Q _18614_/X _18615_/X VGND VGND VPWR
+ VPWR _18688_/X sky130_fd_sc_hd__mux4_1
X_30966_ _35707_/Q _29191_/X _30974_/S VGND VGND VPWR VPWR _30967_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32705_ _36159_/CLK _32705_/D VGND VGND VPWR VPWR _32705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17639_ _17352_/X _17637_/X _17638_/X _17355_/X VGND VGND VPWR VPWR _17639_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33685_ _33685_/CLK _33685_/D VGND VGND VPWR VPWR _33685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30897_ _35674_/Q _29089_/X _30911_/S VGND VGND VPWR VPWR _30898_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32636_ _36092_/CLK _32636_/D VGND VGND VPWR VPWR _32636_/Q sky130_fd_sc_hd__dfxtp_1
X_20650_ _22362_/A VGND VGND VPWR VPWR _22595_/A sky130_fd_sc_hd__buf_12
X_35424_ _35808_/CLK _35424_/D VGND VGND VPWR VPWR _35424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19309_ _19096_/X _19305_/X _19308_/X _19099_/X VGND VGND VPWR VPWR _19309_/X sky130_fd_sc_hd__a22o_1
X_35355_ _35869_/CLK _35355_/D VGND VGND VPWR VPWR _35355_/Q sky130_fd_sc_hd__dfxtp_1
X_20581_ input72/X VGND VGND VPWR VPWR _20659_/A sky130_fd_sc_hd__buf_8
XFILLER_220_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32567_ _36023_/CLK _32567_/D VGND VGND VPWR VPWR _32567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22320_ _22320_/A _22320_/B _22320_/C _22320_/D VGND VGND VPWR VPWR _22321_/A sky130_fd_sc_hd__or4_4
X_34306_ _34306_/CLK _34306_/D VGND VGND VPWR VPWR _34306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31518_ _31518_/A VGND VGND VPWR VPWR _35968_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35286_ _35286_/CLK _35286_/D VGND VGND VPWR VPWR _35286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32498_ _36019_/CLK _32498_/D VGND VGND VPWR VPWR _32498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22251_ _22251_/A VGND VGND VPWR VPWR _36218_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34237_ _34302_/CLK _34237_/D VGND VGND VPWR VPWR _34237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31449_ _23142_/X _35936_/Q _31451_/S VGND VGND VPWR VPWR _31450_/A sky130_fd_sc_hd__mux2_1
X_21202_ _20949_/X _21200_/X _21201_/X _20955_/X VGND VGND VPWR VPWR _21202_/X sky130_fd_sc_hd__a22o_1
XFILLER_219_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22182_ _22107_/X _22180_/X _22181_/X _22112_/X VGND VGND VPWR VPWR _22182_/X sky130_fd_sc_hd__a22o_1
X_34168_ _36152_/CLK _34168_/D VGND VGND VPWR VPWR _34168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21133_ _21129_/X _21132_/X _21022_/X VGND VGND VPWR VPWR _21157_/A sky130_fd_sc_hd__o21ba_1
X_33119_ _36124_/CLK _33119_/D VGND VGND VPWR VPWR _33119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26990_ input50/X VGND VGND VPWR VPWR _26990_/X sky130_fd_sc_hd__buf_4
XFILLER_133_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34099_ _34291_/CLK _34099_/D VGND VGND VPWR VPWR _34099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21064_ _20743_/X _21062_/X _21063_/X _20746_/X VGND VGND VPWR VPWR _21064_/X sky130_fd_sc_hd__a22o_1
X_25941_ _25088_/X _33389_/Q _25957_/S VGND VGND VPWR VPWR _25942_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20015_ _19802_/X _20011_/X _20014_/X _19805_/X VGND VGND VPWR VPWR _20015_/X sky130_fd_sc_hd__a22o_1
XFILLER_154_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28660_ _28660_/A VGND VGND VPWR VPWR _34645_/D sky130_fd_sc_hd__clkbuf_1
X_25872_ _25186_/X _33357_/Q _25872_/S VGND VGND VPWR VPWR _25873_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27611_ _34148_/Q _24314_/X _27625_/S VGND VGND VPWR VPWR _27612_/A sky130_fd_sc_hd__mux2_1
X_24823_ _23031_/X _32895_/Q _24823_/S VGND VGND VPWR VPWR _24824_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28591_ _26943_/X _34613_/Q _28591_/S VGND VGND VPWR VPWR _28592_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27542_ _27542_/A VGND VGND VPWR VPWR _34116_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24754_ _22929_/X _32862_/Q _24760_/S VGND VGND VPWR VPWR _24755_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21966_ _21962_/X _21965_/X _21761_/X VGND VGND VPWR VPWR _21967_/D sky130_fd_sc_hd__o21ba_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23705_ _22883_/X _32399_/Q _23721_/S VGND VGND VPWR VPWR _23706_/A sky130_fd_sc_hd__mux2_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20917_ _20743_/X _20913_/X _20916_/X _20746_/X VGND VGND VPWR VPWR _20917_/X sky130_fd_sc_hd__a22o_1
XFILLER_27_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27473_ _27473_/A VGND VGND VPWR VPWR _34083_/D sky130_fd_sc_hd__clkbuf_1
X_24685_ _24685_/A VGND VGND VPWR VPWR _32830_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21897_ _21897_/A _21897_/B _21897_/C _21897_/D VGND VGND VPWR VPWR _21898_/A sky130_fd_sc_hd__or4_1
XFILLER_203_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29212_ _29212_/A VGND VGND VPWR VPWR _34881_/D sky130_fd_sc_hd__clkbuf_1
X_26424_ _25004_/X _33618_/Q _26434_/S VGND VGND VPWR VPWR _26425_/A sky130_fd_sc_hd__mux2_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20848_ _33235_/Q _36115_/Q _33107_/Q _33043_/Q _20620_/X _20621_/X VGND VGND VPWR
+ VPWR _20848_/X sky130_fd_sc_hd__mux4_1
X_23636_ _32368_/Q _23250_/X _23646_/S VGND VGND VPWR VPWR _23637_/A sky130_fd_sc_hd__mux2_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29143_ _29143_/A VGND VGND VPWR VPWR _34859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26355_ _26355_/A VGND VGND VPWR VPWR _33585_/D sky130_fd_sc_hd__clkbuf_1
X_20779_ _20743_/X _20777_/X _20778_/X _20746_/X VGND VGND VPWR VPWR _20779_/X sky130_fd_sc_hd__a22o_1
XFILLER_204_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23567_ _32335_/Q _23090_/X _23583_/S VGND VGND VPWR VPWR _23568_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25306_ _25162_/X _33093_/Q _25314_/S VGND VGND VPWR VPWR _25307_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22518_ _33026_/Q _32962_/Q _32898_/Q _32834_/Q _22295_/X _22296_/X VGND VGND VPWR
+ VPWR _22518_/X sky130_fd_sc_hd__mux4_1
X_29074_ _34837_/Q _29073_/X _29080_/S VGND VGND VPWR VPWR _29075_/A sky130_fd_sc_hd__mux2_1
X_26286_ _26286_/A VGND VGND VPWR VPWR _33552_/D sky130_fd_sc_hd__clkbuf_1
X_23498_ _23498_/A VGND VGND VPWR VPWR _32303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28025_ _28025_/A VGND VGND VPWR VPWR _34344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22449_ _22300_/X _22445_/X _22448_/X _22303_/X VGND VGND VPWR VPWR _22449_/X sky130_fd_sc_hd__a22o_1
X_25237_ _25060_/X _33060_/Q _25251_/S VGND VGND VPWR VPWR _25238_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25168_ input53/X VGND VGND VPWR VPWR _25168_/X sky130_fd_sc_hd__clkbuf_4
X_24119_ _22892_/X _32594_/Q _24129_/S VGND VGND VPWR VPWR _24120_/A sky130_fd_sc_hd__mux2_1
X_17990_ _35588_/Q _35524_/Q _35460_/Q _35396_/Q _17956_/X _17957_/X VGND VGND VPWR
+ VPWR _17990_/X sky130_fd_sc_hd__mux4_1
X_25099_ _25099_/A VGND VGND VPWR VPWR _33008_/D sky130_fd_sc_hd__clkbuf_1
X_29976_ _35238_/Q _29126_/X _29986_/S VGND VGND VPWR VPWR _29977_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28927_ _34772_/Q _24264_/X _28933_/S VGND VGND VPWR VPWR _28928_/A sky130_fd_sc_hd__mux2_1
X_16941_ _35046_/Q _34982_/Q _34918_/Q _34854_/Q _16803_/X _16804_/X VGND VGND VPWR
+ VPWR _16941_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19660_ _20013_/A VGND VGND VPWR VPWR _19660_/X sky130_fd_sc_hd__buf_4
X_16872_ _17712_/A VGND VGND VPWR VPWR _16872_/X sky130_fd_sc_hd__clkbuf_8
X_28858_ _28858_/A VGND VGND VPWR VPWR _34739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18611_ _34261_/Q _34197_/Q _34133_/Q _34069_/Q _18305_/X _18307_/X VGND VGND VPWR
+ VPWR _18611_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27809_ _34242_/Q _24407_/X _27823_/S VGND VGND VPWR VPWR _27810_/A sky130_fd_sc_hd__mux2_1
XTAP_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19591_ _35312_/Q _35248_/Q _35184_/Q _32304_/Q _19306_/X _19307_/X VGND VGND VPWR
+ VPWR _19591_/X sky130_fd_sc_hd__mux4_1
X_28789_ _28789_/A VGND VGND VPWR VPWR _34706_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ _18436_/X _18540_/X _18541_/X _18441_/X VGND VGND VPWR VPWR _18542_/X sky130_fd_sc_hd__a22o_1
XTAP_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30820_ _30868_/S VGND VGND VPWR VPWR _30839_/S sky130_fd_sc_hd__clkbuf_8
XTAP_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30751_ _23108_/X _35605_/Q _30755_/S VGND VGND VPWR VPWR _30752_/A sky130_fd_sc_hd__mux2_1
X_18473_ _18473_/A VGND VGND VPWR VPWR _32080_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_350 _36205_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_361 _36207_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_372 _36208_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17424_ _35764_/Q _35124_/Q _34484_/Q _33844_/Q _17140_/X _17141_/X VGND VGND VPWR
+ VPWR _17424_/X sky130_fd_sc_hd__mux4_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33470_ _34303_/CLK _33470_/D VGND VGND VPWR VPWR _33470_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_383 _36209_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30682_ _30682_/A VGND VGND VPWR VPWR _35572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_394 _36210_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32421_ _35942_/CLK _32421_/D VGND VGND VPWR VPWR _32421_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _17865_/A VGND VGND VPWR VPWR _17355_/X sky130_fd_sc_hd__buf_4
XFILLER_18_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35140_ _35780_/CLK _35140_/D VGND VGND VPWR VPWR _35140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16306_ _16087_/X _16304_/X _16305_/X _16097_/X VGND VGND VPWR VPWR _16306_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32352_ _36001_/CLK _32352_/D VGND VGND VPWR VPWR _32352_/Q sky130_fd_sc_hd__dfxtp_1
X_17286_ _16999_/X _17284_/X _17285_/X _17002_/X VGND VGND VPWR VPWR _17286_/X sky130_fd_sc_hd__a22o_1
XFILLER_201_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19025_ _19019_/X _19024_/X _18741_/X VGND VGND VPWR VPWR _19033_/C sky130_fd_sc_hd__o21ba_1
X_31303_ _31303_/A VGND VGND VPWR VPWR _35866_/D sky130_fd_sc_hd__clkbuf_1
X_16237_ _16233_/X _16236_/X _16100_/X VGND VGND VPWR VPWR _16238_/D sky130_fd_sc_hd__o21ba_1
X_35071_ _35982_/CLK _35071_/D VGND VGND VPWR VPWR _35071_/Q sky130_fd_sc_hd__dfxtp_1
X_32283_ _36201_/CLK _32283_/D VGND VGND VPWR VPWR _32283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34022_ _34087_/CLK _34022_/D VGND VGND VPWR VPWR _34022_/Q sky130_fd_sc_hd__dfxtp_1
X_31234_ _35834_/Q input39/X _31244_/S VGND VGND VPWR VPWR _31235_/A sky130_fd_sc_hd__mux2_1
X_16168_ _34512_/Q _32400_/Q _34384_/Q _34320_/Q _16166_/X _16167_/X VGND VGND VPWR
+ VPWR _16168_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31165_ _35801_/Q input3/X _31181_/S VGND VGND VPWR VPWR _31166_/A sky130_fd_sc_hd__mux2_1
X_16099_ input70/X input69/X VGND VGND VPWR VPWR _17867_/A sky130_fd_sc_hd__or2b_4
XFILLER_173_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30116_ _30116_/A VGND VGND VPWR VPWR _35304_/D sky130_fd_sc_hd__clkbuf_1
X_19927_ _33274_/Q _36154_/Q _33146_/Q _33082_/Q _19711_/X _19712_/X VGND VGND VPWR
+ VPWR _19927_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35973_ _35973_/CLK _35973_/D VGND VGND VPWR VPWR _35973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31096_ _31096_/A VGND VGND VPWR VPWR _35768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30047_ _35272_/Q _29231_/X _30049_/S VGND VGND VPWR VPWR _30048_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34924_ _35313_/CLK _34924_/D VGND VGND VPWR VPWR _34924_/Q sky130_fd_sc_hd__dfxtp_1
X_19858_ _20211_/A VGND VGND VPWR VPWR _19858_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_151_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18809_ _35802_/Q _32177_/Q _35674_/Q _35610_/Q _18554_/X _18555_/X VGND VGND VPWR
+ VPWR _18809_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34855_ _35943_/CLK _34855_/D VGND VGND VPWR VPWR _34855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19789_ _20142_/A VGND VGND VPWR VPWR _19789_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_3_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33806_ _35727_/CLK _33806_/D VGND VGND VPWR VPWR _33806_/Q sky130_fd_sc_hd__dfxtp_1
X_21820_ _21599_/X _21818_/X _21819_/X _21602_/X VGND VGND VPWR VPWR _21820_/X sky130_fd_sc_hd__a22o_1
X_34786_ _35300_/CLK _34786_/D VGND VGND VPWR VPWR _34786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31998_ _33946_/CLK _31998_/D VGND VGND VPWR VPWR _31998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21751_ _35308_/Q _35244_/Q _35180_/Q _32300_/Q _21606_/X _21607_/X VGND VGND VPWR
+ VPWR _21751_/X sky130_fd_sc_hd__mux4_1
X_33737_ _34817_/CLK _33737_/D VGND VGND VPWR VPWR _33737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30949_ _35699_/Q _29166_/X _30953_/S VGND VGND VPWR VPWR _30950_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20702_ _20702_/A _20702_/B _20702_/C _20702_/D VGND VGND VPWR VPWR _20703_/A sky130_fd_sc_hd__or4_4
XFILLER_19_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24470_ _24470_/A VGND VGND VPWR VPWR _32729_/D sky130_fd_sc_hd__clkbuf_1
X_21682_ _34538_/Q _32426_/Q _34410_/Q _34346_/Q _21472_/X _21473_/X VGND VGND VPWR
+ VPWR _21682_/X sky130_fd_sc_hd__mux4_1
X_33668_ _33795_/CLK _33668_/D VGND VGND VPWR VPWR _33668_/Q sky130_fd_sc_hd__dfxtp_1
X_35407_ _35791_/CLK _35407_/D VGND VGND VPWR VPWR _35407_/Q sky130_fd_sc_hd__dfxtp_1
X_23421_ _32269_/Q _23345_/X _23421_/S VGND VGND VPWR VPWR _23422_/A sky130_fd_sc_hd__mux2_1
X_20633_ _22429_/A VGND VGND VPWR VPWR _20633_/X sky130_fd_sc_hd__buf_4
XFILLER_149_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32619_ _36075_/CLK _32619_/D VGND VGND VPWR VPWR _32619_/Q sky130_fd_sc_hd__dfxtp_1
X_33599_ _33729_/CLK _33599_/D VGND VGND VPWR VPWR _33599_/Q sky130_fd_sc_hd__dfxtp_1
X_26140_ _25183_/X _33484_/Q _26142_/S VGND VGND VPWR VPWR _26141_/A sky130_fd_sc_hd__mux2_1
X_23352_ _23421_/S VGND VGND VPWR VPWR _23371_/S sky130_fd_sc_hd__buf_4
X_35338_ _35338_/CLK _35338_/D VGND VGND VPWR VPWR _35338_/Q sky130_fd_sc_hd__dfxtp_1
X_20564_ _18297_/X _20562_/X _20563_/X _18303_/X VGND VGND VPWR VPWR _20564_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22303_ _22458_/A VGND VGND VPWR VPWR _22303_/X sky130_fd_sc_hd__buf_4
XFILLER_149_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23283_ input39/X VGND VGND VPWR VPWR _23283_/X sky130_fd_sc_hd__clkbuf_4
X_26071_ _25081_/X _33451_/Q _26071_/S VGND VGND VPWR VPWR _26072_/A sky130_fd_sc_hd__mux2_1
X_35269_ _35333_/CLK _35269_/D VGND VGND VPWR VPWR _35269_/Q sky130_fd_sc_hd__dfxtp_1
X_20495_ _32523_/Q _32395_/Q _32075_/Q _36043_/Q _20282_/X _19307_/A VGND VGND VPWR
+ VPWR _20495_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_23_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_23_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_106_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22234_ _35834_/Q _32212_/Q _35706_/Q _35642_/Q _21913_/X _21914_/X VGND VGND VPWR
+ VPWR _22234_/X sky130_fd_sc_hd__mux4_1
X_25022_ input2/X VGND VGND VPWR VPWR _25022_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_118_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29830_ _35169_/Q _29110_/X _29830_/S VGND VGND VPWR VPWR _29831_/A sky130_fd_sc_hd__mux2_1
XFILLER_234_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22165_ _33016_/Q _32952_/Q _32888_/Q _32824_/Q _21942_/X _21943_/X VGND VGND VPWR
+ VPWR _22165_/X sky130_fd_sc_hd__mux4_1
XTAP_6904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21116_ _34778_/Q _34714_/Q _34650_/Q _34586_/Q _20829_/X _20830_/X VGND VGND VPWR
+ VPWR _21116_/X sky130_fd_sc_hd__mux4_1
XTAP_6937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29761_ _35136_/Q _29206_/X _29779_/S VGND VGND VPWR VPWR _29762_/A sky130_fd_sc_hd__mux2_1
XTAP_6948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26973_ _26973_/A VGND VGND VPWR VPWR _33854_/D sky130_fd_sc_hd__clkbuf_1
X_22096_ _21947_/X _22092_/X _22095_/X _21950_/X VGND VGND VPWR VPWR _22096_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28712_ _26922_/X _34670_/Q _28726_/S VGND VGND VPWR VPWR _28713_/A sky130_fd_sc_hd__mux2_1
X_25924_ _25063_/X _33381_/Q _25936_/S VGND VGND VPWR VPWR _25925_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21047_ _21043_/X _21044_/X _21045_/X _21046_/X VGND VGND VPWR VPWR _21047_/X sky130_fd_sc_hd__a22o_1
X_29692_ _29692_/A VGND VGND VPWR VPWR _35103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28643_ _28778_/B _28643_/B VGND VGND VPWR VPWR _28776_/S sky130_fd_sc_hd__nand2_8
XFILLER_130_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25855_ _25855_/A VGND VGND VPWR VPWR _33348_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24806_ _24806_/A VGND VGND VPWR VPWR _32886_/D sky130_fd_sc_hd__clkbuf_1
X_28574_ _28574_/A VGND VGND VPWR VPWR _34604_/D sky130_fd_sc_hd__clkbuf_1
X_25786_ _25786_/A VGND VGND VPWR VPWR _33315_/D sky130_fd_sc_hd__clkbuf_1
X_22998_ _22997_/X _32052_/Q _23001_/S VGND VGND VPWR VPWR _22999_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27525_ _27525_/A VGND VGND VPWR VPWR _34108_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_991 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24737_ _22904_/X _32854_/Q _24739_/S VGND VGND VPWR VPWR _24738_/A sky130_fd_sc_hd__mux2_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21949_ _35762_/Q _35122_/Q _34482_/Q _33842_/Q _21740_/X _21741_/X VGND VGND VPWR
+ VPWR _21949_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27456_ _27456_/A VGND VGND VPWR VPWR _34075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24668_ _23003_/X _32822_/Q _24686_/S VGND VGND VPWR VPWR _24669_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26407_ _26407_/A VGND VGND VPWR VPWR _33610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23619_ _32360_/Q _23223_/X _23625_/S VGND VGND VPWR VPWR _23620_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27387_ _34043_/Q _24385_/X _27395_/S VGND VGND VPWR VPWR _27388_/A sky130_fd_sc_hd__mux2_1
X_24599_ _24599_/A VGND VGND VPWR VPWR _32789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17140_ _17994_/A VGND VGND VPWR VPWR _17140_/X sky130_fd_sc_hd__buf_6
X_29126_ input17/X VGND VGND VPWR VPWR _29126_/X sky130_fd_sc_hd__buf_2
XFILLER_204_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26338_ _26338_/A VGND VGND VPWR VPWR _33577_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29057_ _29057_/A VGND VGND VPWR VPWR _34831_/D sky130_fd_sc_hd__clkbuf_1
X_17071_ _35754_/Q _35114_/Q _34474_/Q _33834_/Q _16787_/X _16788_/X VGND VGND VPWR
+ VPWR _17071_/X sky130_fd_sc_hd__mux4_1
X_26269_ _25174_/X _33545_/Q _26269_/S VGND VGND VPWR VPWR _26270_/A sky130_fd_sc_hd__mux2_1
X_16022_ _33230_/Q _36110_/Q _33102_/Q _33038_/Q _16020_/X _16021_/X VGND VGND VPWR
+ VPWR _16022_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28008_ _28008_/A VGND VGND VPWR VPWR _34336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_1099 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17973_ _17901_/X _17971_/X _17972_/X _17906_/X VGND VGND VPWR VPWR _17973_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29959_ _35230_/Q _29101_/X _29965_/S VGND VGND VPWR VPWR _29960_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16924_ _32486_/Q _32358_/Q _32038_/Q _36006_/Q _16923_/X _16711_/X VGND VGND VPWR
+ VPWR _16924_/X sky130_fd_sc_hd__mux4_1
X_19712_ _20070_/A VGND VGND VPWR VPWR _19712_/X sky130_fd_sc_hd__clkbuf_4
X_32970_ _35979_/CLK _32970_/D VGND VGND VPWR VPWR _32970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31921_ _31948_/S VGND VGND VPWR VPWR _31940_/S sky130_fd_sc_hd__buf_6
X_16855_ _32740_/Q _32676_/Q _32612_/Q _36068_/Q _16566_/X _16703_/X VGND VGND VPWR
+ VPWR _16855_/X sky130_fd_sc_hd__mux4_1
X_19643_ _20130_/A VGND VGND VPWR VPWR _19643_/X sky130_fd_sc_hd__buf_4
XFILLER_226_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34640_ _36216_/CLK _34640_/D VGND VGND VPWR VPWR _34640_/Q sky130_fd_sc_hd__dfxtp_1
X_19574_ _33264_/Q _36144_/Q _33136_/Q _33072_/Q _19358_/X _19359_/X VGND VGND VPWR
+ VPWR _19574_/X sky130_fd_sc_hd__mux4_1
X_31852_ _23139_/X _36127_/Q _31856_/S VGND VGND VPWR VPWR _31853_/A sky130_fd_sc_hd__mux2_1
X_16786_ _35810_/Q _32186_/Q _35682_/Q _35618_/Q _16607_/X _16608_/X VGND VGND VPWR
+ VPWR _16786_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18525_ _35538_/Q _35474_/Q _35410_/Q _35346_/Q _18491_/X _18492_/X VGND VGND VPWR
+ VPWR _18525_/X sky130_fd_sc_hd__mux4_1
X_30803_ _30803_/A VGND VGND VPWR VPWR _35629_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34571_ _35147_/CLK _34571_/D VGND VGND VPWR VPWR _34571_/Q sky130_fd_sc_hd__dfxtp_1
X_31783_ _31783_/A VGND VGND VPWR VPWR _36094_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30734_ _30734_/A VGND VGND VPWR VPWR _35597_/D sky130_fd_sc_hd__clkbuf_1
X_18456_ _35792_/Q _32166_/Q _35664_/Q _35600_/Q _18345_/X _18346_/X VGND VGND VPWR
+ VPWR _18456_/X sky130_fd_sc_hd__mux4_1
X_33522_ _33775_/CLK _33522_/D VGND VGND VPWR VPWR _33522_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_180 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_191 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17407_ _17403_/X _17406_/X _17128_/X VGND VGND VPWR VPWR _17439_/A sky130_fd_sc_hd__o21ba_1
XFILLER_226_1471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33453_ _34293_/CLK _33453_/D VGND VGND VPWR VPWR _33453_/Q sky130_fd_sc_hd__dfxtp_1
X_18387_ _19454_/A VGND VGND VPWR VPWR _18387_/X sky130_fd_sc_hd__buf_4
X_30665_ _35564_/Q _29144_/X _30683_/S VGND VGND VPWR VPWR _30666_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32404_ _34775_/CLK _32404_/D VGND VGND VPWR VPWR _32404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17338_ _32754_/Q _32690_/Q _32626_/Q _36082_/Q _17272_/X _17056_/X VGND VGND VPWR
+ VPWR _17338_/X sky130_fd_sc_hd__mux4_1
X_36172_ _36172_/CLK _36172_/D VGND VGND VPWR VPWR _36172_/Q sky130_fd_sc_hd__dfxtp_1
X_33384_ _33512_/CLK _33384_/D VGND VGND VPWR VPWR _33384_/Q sky130_fd_sc_hd__dfxtp_1
X_30596_ _23342_/X _35532_/Q _30598_/S VGND VGND VPWR VPWR _30597_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32335_ _36041_/CLK _32335_/D VGND VGND VPWR VPWR _32335_/Q sky130_fd_sc_hd__dfxtp_1
X_35123_ _35829_/CLK _35123_/D VGND VGND VPWR VPWR _35123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17269_ _34032_/Q _33968_/Q _33904_/Q _32240_/Q _17020_/X _17021_/X VGND VGND VPWR
+ VPWR _17269_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19008_ _20206_/A VGND VGND VPWR VPWR _19008_/X sky130_fd_sc_hd__clkbuf_4
X_35054_ _35054_/CLK _35054_/D VGND VGND VPWR VPWR _35054_/Q sky130_fd_sc_hd__dfxtp_1
X_32266_ _35851_/CLK _32266_/D VGND VGND VPWR VPWR _32266_/Q sky130_fd_sc_hd__dfxtp_1
X_20280_ _33284_/Q _36164_/Q _33156_/Q _33092_/Q _20064_/X _20065_/X VGND VGND VPWR
+ VPWR _20280_/X sky130_fd_sc_hd__mux4_1
XFILLER_161_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34005_ _35280_/CLK _34005_/D VGND VGND VPWR VPWR _34005_/Q sky130_fd_sc_hd__dfxtp_1
X_31217_ _35826_/Q input30/X _31223_/S VGND VGND VPWR VPWR _31218_/A sky130_fd_sc_hd__mux2_1
X_32197_ _35950_/CLK _32197_/D VGND VGND VPWR VPWR _32197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31148_ _35793_/Q input34/X _31160_/S VGND VGND VPWR VPWR _31149_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23970_ _23074_/X _32525_/Q _23970_/S VGND VGND VPWR VPWR _23971_/A sky130_fd_sc_hd__mux2_1
XTAP_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31079_ _31079_/A VGND VGND VPWR VPWR _35760_/D sky130_fd_sc_hd__clkbuf_1
X_35956_ _35956_/CLK _35956_/D VGND VGND VPWR VPWR _35956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22921_ _22920_/X _32027_/Q _22939_/S VGND VGND VPWR VPWR _22922_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34907_ _35166_/CLK _34907_/D VGND VGND VPWR VPWR _34907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35887_ _35951_/CLK _35887_/D VGND VGND VPWR VPWR _35887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25640_ _25640_/A VGND VGND VPWR VPWR _33247_/D sky130_fd_sc_hd__clkbuf_1
X_22852_ _32781_/Q _32717_/Q _32653_/Q _36109_/Q _22578_/X _21473_/A VGND VGND VPWR
+ VPWR _22852_/X sky130_fd_sc_hd__mux4_1
X_34838_ _35028_/CLK _34838_/D VGND VGND VPWR VPWR _34838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21803_ _33518_/Q _33454_/Q _33390_/Q _33326_/Q _21723_/X _21724_/X VGND VGND VPWR
+ VPWR _21803_/X sky130_fd_sc_hd__mux4_1
X_25571_ _33216_/Q _24400_/X _25589_/S VGND VGND VPWR VPWR _25572_/A sky130_fd_sc_hd__mux2_1
X_22783_ _22783_/A _22783_/B _22783_/C _22783_/D VGND VGND VPWR VPWR _22784_/A sky130_fd_sc_hd__or4_4
X_34769_ _35280_/CLK _34769_/D VGND VGND VPWR VPWR _34769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27310_ _27310_/A VGND VGND VPWR VPWR _34006_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24522_ _24522_/A VGND VGND VPWR VPWR _32754_/D sky130_fd_sc_hd__clkbuf_1
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28290_ _34470_/Q _24320_/X _28300_/S VGND VGND VPWR VPWR _28291_/A sky130_fd_sc_hd__mux2_1
X_21734_ _33004_/Q _32940_/Q _32876_/Q _32812_/Q _21589_/X _21590_/X VGND VGND VPWR
+ VPWR _21734_/X sky130_fd_sc_hd__mux4_1
XFILLER_212_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27241_ _27289_/S VGND VGND VPWR VPWR _27260_/S sky130_fd_sc_hd__buf_4
X_24453_ _24453_/A VGND VGND VPWR VPWR _32721_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21665_ _32490_/Q _32362_/Q _32042_/Q _36010_/Q _21523_/X _21664_/X VGND VGND VPWR
+ VPWR _21665_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23404_ _23404_/A VGND VGND VPWR VPWR _32260_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27172_ _26844_/X _33941_/Q _27176_/S VGND VGND VPWR VPWR _27173_/A sky130_fd_sc_hd__mux2_1
X_20616_ _22578_/A VGND VGND VPWR VPWR _22462_/A sky130_fd_sc_hd__buf_12
X_24384_ _24384_/A VGND VGND VPWR VPWR _32698_/D sky130_fd_sc_hd__clkbuf_1
X_21596_ _35752_/Q _35112_/Q _34472_/Q _33832_/Q _21387_/X _21388_/X VGND VGND VPWR
+ VPWR _21596_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26123_ _26123_/A VGND VGND VPWR VPWR _33475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23335_ _23335_/A VGND VGND VPWR VPWR _32229_/D sky130_fd_sc_hd__clkbuf_1
X_20547_ _18314_/X _20545_/X _20546_/X _18323_/X VGND VGND VPWR VPWR _20547_/X sky130_fd_sc_hd__a22o_1
XFILLER_165_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26054_ _26054_/A VGND VGND VPWR VPWR _33442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20478_ _18344_/X _20476_/X _20477_/X _18354_/X VGND VGND VPWR VPWR _20478_/X sky130_fd_sc_hd__a22o_1
XFILLER_3_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23266_ _23266_/A VGND VGND VPWR VPWR _32206_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25005_ _25004_/X _32978_/Q _25020_/S VGND VGND VPWR VPWR _25006_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22217_ _22217_/A VGND VGND VPWR VPWR _36217_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23197_ _32181_/Q _23136_/X _23206_/S VGND VGND VPWR VPWR _23198_/A sky130_fd_sc_hd__mux2_1
XTAP_6701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22148_ _22501_/A VGND VGND VPWR VPWR _22148_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29813_ _29813_/A VGND VGND VPWR VPWR _35160_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26956_ input38/X VGND VGND VPWR VPWR _26956_/X sky130_fd_sc_hd__clkbuf_4
X_29744_ _35128_/Q _29182_/X _29758_/S VGND VGND VPWR VPWR _29745_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22079_ _34038_/Q _33974_/Q _33910_/Q _32246_/Q _21973_/X _21974_/X VGND VGND VPWR
+ VPWR _22079_/X sky130_fd_sc_hd__mux4_1
XTAP_6789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25907_ _25038_/X _33373_/Q _25915_/S VGND VGND VPWR VPWR _25908_/A sky130_fd_sc_hd__mux2_1
X_29675_ _29675_/A VGND VGND VPWR VPWR _35095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26887_ _26887_/A VGND VGND VPWR VPWR _33826_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28626_ _28626_/A VGND VGND VPWR VPWR _34629_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16640_ _16634_/X _16639_/X _16430_/X _16431_/X VGND VGND VPWR VPWR _16661_/B sky130_fd_sc_hd__o211a_2
X_25838_ _25838_/A VGND VGND VPWR VPWR _33340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28557_ _28557_/A VGND VGND VPWR VPWR _34596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16571_ _32476_/Q _32348_/Q _32028_/Q _35996_/Q _16570_/X _16358_/X VGND VGND VPWR
+ VPWR _16571_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25769_ _25769_/A VGND VGND VPWR VPWR _33307_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18310_ input81/X input82/X VGND VGND VPWR VPWR _20134_/A sky130_fd_sc_hd__or2b_4
XFILLER_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27508_ _27508_/A VGND VGND VPWR VPWR _34100_/D sky130_fd_sc_hd__clkbuf_1
X_19290_ _20130_/A VGND VGND VPWR VPWR _19290_/X sky130_fd_sc_hd__buf_6
X_28488_ _26990_/X _34564_/Q _28498_/S VGND VGND VPWR VPWR _28489_/A sky130_fd_sc_hd__mux2_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18241_ _16056_/X _18239_/X _18240_/X _16068_/X VGND VGND VPWR VPWR _18241_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27439_ _27439_/A VGND VGND VPWR VPWR _34067_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1019 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18172_ _35594_/Q _35530_/Q _35466_/Q _35402_/Q _17956_/X _17957_/X VGND VGND VPWR
+ VPWR _18172_/X sky130_fd_sc_hd__mux4_1
X_30450_ _30450_/A VGND VGND VPWR VPWR _35462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29109_ _29109_/A VGND VGND VPWR VPWR _34848_/D sky130_fd_sc_hd__clkbuf_1
X_17123_ _17829_/A VGND VGND VPWR VPWR _17123_/X sky130_fd_sc_hd__buf_4
XFILLER_102_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30381_ _30381_/A VGND VGND VPWR VPWR _35429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32120_ _35814_/CLK _32120_/D VGND VGND VPWR VPWR _32120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17054_ _17050_/X _17053_/X _16775_/X VGND VGND VPWR VPWR _17086_/A sky130_fd_sc_hd__o21ba_1
XFILLER_125_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16005_ _17956_/A VGND VGND VPWR VPWR _16005_/X sky130_fd_sc_hd__clkbuf_8
X_32051_ _36019_/CLK _32051_/D VGND VGND VPWR VPWR _32051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31002_ _31002_/A VGND VGND VPWR VPWR _35724_/D sky130_fd_sc_hd__clkbuf_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35810_ _35811_/CLK _35810_/D VGND VGND VPWR VPWR _35810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17956_ _17956_/A VGND VGND VPWR VPWR _17956_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35741_ _35869_/CLK _35741_/D VGND VGND VPWR VPWR _35741_/Q sky130_fd_sc_hd__dfxtp_1
X_16907_ _35045_/Q _34981_/Q _34917_/Q _34853_/Q _16803_/X _16804_/X VGND VGND VPWR
+ VPWR _16907_/X sky130_fd_sc_hd__mux4_1
X_17887_ _17700_/X _17885_/X _17886_/X _17703_/X VGND VGND VPWR VPWR _17887_/X sky130_fd_sc_hd__a22o_1
X_32953_ _36090_/CLK _32953_/D VGND VGND VPWR VPWR _32953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31904_ _31904_/A VGND VGND VPWR VPWR _36151_/D sky130_fd_sc_hd__clkbuf_1
X_19626_ _35057_/Q _34993_/Q _34929_/Q _34865_/Q _19456_/X _19457_/X VGND VGND VPWR
+ VPWR _19626_/X sky130_fd_sc_hd__mux4_1
X_16838_ _16801_/X _16836_/X _16837_/X _16806_/X VGND VGND VPWR VPWR _16838_/X sky130_fd_sc_hd__a22o_1
X_35672_ _35675_/CLK _35672_/D VGND VGND VPWR VPWR _35672_/Q sky130_fd_sc_hd__dfxtp_1
X_32884_ _35765_/CLK _32884_/D VGND VGND VPWR VPWR _32884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34623_ _35837_/CLK _34623_/D VGND VGND VPWR VPWR _34623_/Q sky130_fd_sc_hd__dfxtp_1
X_31835_ _23114_/X _36119_/Q _31835_/S VGND VGND VPWR VPWR _31836_/A sky130_fd_sc_hd__mux2_1
X_19557_ _35311_/Q _35247_/Q _35183_/Q _32303_/Q _19306_/X _19307_/X VGND VGND VPWR
+ VPWR _19557_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16769_ _16489_/X _16767_/X _16768_/X _16494_/X VGND VGND VPWR VPWR _16769_/X sky130_fd_sc_hd__a22o_1
XFILLER_213_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18508_ _18436_/X _18506_/X _18507_/X _18441_/X VGND VGND VPWR VPWR _18508_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34554_ _35771_/CLK _34554_/D VGND VGND VPWR VPWR _34554_/Q sky130_fd_sc_hd__dfxtp_1
X_31766_ _36086_/Q input35/X _31784_/S VGND VGND VPWR VPWR _31767_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19488_ _19449_/X _19486_/X _19487_/X _19452_/X VGND VGND VPWR VPWR _19488_/X sky130_fd_sc_hd__a22o_1
X_30717_ _35589_/Q _29222_/X _30725_/S VGND VGND VPWR VPWR _30718_/A sky130_fd_sc_hd__mux2_1
X_33505_ _34145_/CLK _33505_/D VGND VGND VPWR VPWR _33505_/Q sky130_fd_sc_hd__dfxtp_1
X_18439_ _33744_/Q _33680_/Q _33616_/Q _33552_/Q _18437_/X _18438_/X VGND VGND VPWR
+ VPWR _18439_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31697_ _31697_/A VGND VGND VPWR VPWR _36053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34485_ _35828_/CLK _34485_/D VGND VGND VPWR VPWR _34485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36224_ _36228_/CLK _36224_/D VGND VGND VPWR VPWR _36224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21450_ _33508_/Q _33444_/Q _33380_/Q _33316_/Q _21370_/X _21371_/X VGND VGND VPWR
+ VPWR _21450_/X sky130_fd_sc_hd__mux4_1
X_30648_ _35556_/Q _29120_/X _30662_/S VGND VGND VPWR VPWR _30649_/A sky130_fd_sc_hd__mux2_1
X_33436_ _34074_/CLK _33436_/D VGND VGND VPWR VPWR _33436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20401_ _20397_/X _20400_/X _20134_/X VGND VGND VPWR VPWR _20423_/A sky130_fd_sc_hd__o21ba_2
XFILLER_120_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33367_ _36228_/CLK _33367_/D VGND VGND VPWR VPWR _33367_/Q sky130_fd_sc_hd__dfxtp_1
X_36155_ _36156_/CLK _36155_/D VGND VGND VPWR VPWR _36155_/Q sky130_fd_sc_hd__dfxtp_1
X_21381_ _32994_/Q _32930_/Q _32866_/Q _32802_/Q _21236_/X _21237_/X VGND VGND VPWR
+ VPWR _21381_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30579_ _30579_/A VGND VGND VPWR VPWR _35523_/D sky130_fd_sc_hd__clkbuf_1
X_20332_ _20328_/X _20331_/X _20167_/X VGND VGND VPWR VPWR _20333_/D sky130_fd_sc_hd__o21ba_1
XFILLER_174_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23120_ _23120_/A VGND VGND VPWR VPWR _32152_/D sky130_fd_sc_hd__clkbuf_1
X_35106_ _35876_/CLK _35106_/D VGND VGND VPWR VPWR _35106_/Q sky130_fd_sc_hd__dfxtp_1
X_32318_ _36105_/CLK _32318_/D VGND VGND VPWR VPWR _32318_/Q sky130_fd_sc_hd__dfxtp_1
X_33298_ _33940_/CLK _33298_/D VGND VGND VPWR VPWR _33298_/Q sky130_fd_sc_hd__dfxtp_1
X_36086_ _36086_/CLK _36086_/D VGND VGND VPWR VPWR _36086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1086 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23051_ _23050_/X _32069_/Q _23063_/S VGND VGND VPWR VPWR _23052_/A sky130_fd_sc_hd__mux2_1
X_20263_ _35331_/Q _35267_/Q _35203_/Q _32323_/Q _20012_/X _20013_/X VGND VGND VPWR
+ VPWR _20263_/X sky130_fd_sc_hd__mux4_1
X_32249_ _36154_/CLK _32249_/D VGND VGND VPWR VPWR _32249_/Q sky130_fd_sc_hd__dfxtp_1
X_35037_ _35038_/CLK _35037_/D VGND VGND VPWR VPWR _35037_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22002_ _34292_/Q _34228_/Q _34164_/Q _34100_/Q _21689_/X _21690_/X VGND VGND VPWR
+ VPWR _22002_/X sky130_fd_sc_hd__mux4_1
XTAP_6019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20194_ _20155_/X _20192_/X _20193_/X _20158_/X VGND VGND VPWR VPWR _20194_/X sky130_fd_sc_hd__a22o_1
XFILLER_153_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26810_ _26810_/A VGND VGND VPWR VPWR _33800_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27790_ _34233_/Q _24379_/X _27802_/S VGND VGND VPWR VPWR _27791_/A sky130_fd_sc_hd__mux2_1
XFILLER_233_1272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26741_ _26741_/A VGND VGND VPWR VPWR _33767_/D sky130_fd_sc_hd__clkbuf_1
X_23953_ _23953_/A VGND VGND VPWR VPWR _32516_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35939_ _35940_/CLK _35939_/D VGND VGND VPWR VPWR _35939_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_1002 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22904_ input63/X VGND VGND VPWR VPWR _22904_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29460_ _29460_/A VGND VGND VPWR VPWR _34993_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26672_ _26672_/A VGND VGND VPWR VPWR _33735_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23884_ _23884_/A VGND VGND VPWR VPWR _32483_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_905 _26819_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28411_ _28411_/A VGND VGND VPWR VPWR _34527_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_916 _26993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25623_ _25623_/A VGND VGND VPWR VPWR _33239_/D sky130_fd_sc_hd__clkbuf_1
X_22835_ _22831_/X _22834_/X _22453_/A VGND VGND VPWR VPWR _22843_/C sky130_fd_sc_hd__o21ba_1
X_29391_ _29391_/A VGND VGND VPWR VPWR _34960_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_927 _27966_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_938 _29079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_949 _29652_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28342_ _34495_/Q _24397_/X _28342_/S VGND VGND VPWR VPWR _28343_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25554_ _33208_/Q _24376_/X _25568_/S VGND VGND VPWR VPWR _25555_/A sky130_fd_sc_hd__mux2_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22766_ _33034_/Q _32970_/Q _32906_/Q _32842_/Q _20580_/X _20583_/X VGND VGND VPWR
+ VPWR _22766_/X sky130_fd_sc_hd__mux4_1
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24505_ _24505_/A VGND VGND VPWR VPWR _32746_/D sky130_fd_sc_hd__clkbuf_1
X_28273_ _34462_/Q _24295_/X _28279_/S VGND VGND VPWR VPWR _28274_/A sky130_fd_sc_hd__mux2_1
X_21717_ _21713_/X _21716_/X _21408_/X VGND VGND VPWR VPWR _21718_/D sky130_fd_sc_hd__o21ba_1
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25485_ _25485_/A VGND VGND VPWR VPWR _33175_/D sky130_fd_sc_hd__clkbuf_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22697_ _22501_/X _22695_/X _22696_/X _22506_/X VGND VGND VPWR VPWR _22697_/X sky130_fd_sc_hd__a22o_1
XFILLER_227_1098 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27224_ _27224_/A VGND VGND VPWR VPWR _33965_/D sky130_fd_sc_hd__clkbuf_1
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24436_ _24436_/A VGND VGND VPWR VPWR _32715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21648_ _33770_/Q _33706_/Q _33642_/Q _33578_/Q _21443_/X _21444_/X VGND VGND VPWR
+ VPWR _21648_/X sky130_fd_sc_hd__mux4_1
XFILLER_227_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27155_ _27155_/A VGND VGND VPWR VPWR _33933_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_193_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _36105_/CLK sky130_fd_sc_hd__clkbuf_16
X_24367_ _32693_/Q _24366_/X _24367_/S VGND VGND VPWR VPWR _24368_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_80 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21579_ _34280_/Q _34216_/Q _34152_/Q _34088_/Q _21336_/X _21337_/X VGND VGND VPWR
+ VPWR _21579_/X sky130_fd_sc_hd__mux4_1
XANTENNA_91 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26106_ _26106_/A VGND VGND VPWR VPWR _33467_/D sky130_fd_sc_hd__clkbuf_1
X_23318_ _23318_/A VGND VGND VPWR VPWR _32223_/D sky130_fd_sc_hd__clkbuf_1
X_27086_ _26915_/X _33900_/Q _27104_/S VGND VGND VPWR VPWR _27087_/A sky130_fd_sc_hd__mux2_1
X_24298_ input9/X VGND VGND VPWR VPWR _24298_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_181_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26037_ _26037_/A VGND VGND VPWR VPWR _33434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23249_ _23249_/A VGND VGND VPWR VPWR _32200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1304 _16591_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1315 _32124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_1058 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1326 _20134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1337 _20167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17810_ _35839_/Q _32218_/Q _35711_/Q _35647_/Q _17666_/X _17667_/X VGND VGND VPWR
+ VPWR _17810_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1348 _22447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18790_ _20202_/A VGND VGND VPWR VPWR _18790_/X sky130_fd_sc_hd__buf_6
XTAP_5830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27988_ _26850_/X _34327_/Q _27988_/S VGND VGND VPWR VPWR _27989_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1359 _22938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_999 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17741_ _35581_/Q _35517_/Q _35453_/Q _35389_/Q _17603_/X _17604_/X VGND VGND VPWR
+ VPWR _17741_/X sky130_fd_sc_hd__mux4_1
XFILLER_248_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29727_ _35120_/Q _29157_/X _29737_/S VGND VGND VPWR VPWR _29728_/A sky130_fd_sc_hd__mux2_1
X_26939_ _26939_/A VGND VGND VPWR VPWR _33843_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17672_ _33211_/Q _32571_/Q _35963_/Q _35899_/Q _17427_/X _17428_/X VGND VGND VPWR
+ VPWR _17672_/X sky130_fd_sc_hd__mux4_1
X_29658_ _35087_/Q _29055_/X _29674_/S VGND VGND VPWR VPWR _29659_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19411_ _34795_/Q _34731_/Q _34667_/Q _34603_/Q _19235_/X _19236_/X VGND VGND VPWR
+ VPWR _19411_/X sky130_fd_sc_hd__mux4_1
X_16623_ _16623_/A _16623_/B _16623_/C _16623_/D VGND VGND VPWR VPWR _16624_/A sky130_fd_sc_hd__or4_1
X_28609_ _28609_/A VGND VGND VPWR VPWR _34621_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29589_ _29589_/A VGND VGND VPWR VPWR _35054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31620_ _36017_/Q input29/X _31628_/S VGND VGND VPWR VPWR _31621_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16554_ _35035_/Q _34971_/Q _34907_/Q _34843_/Q _16450_/X _16451_/X VGND VGND VPWR
+ VPWR _16554_/X sky130_fd_sc_hd__mux4_1
X_19342_ _34537_/Q _32425_/Q _34409_/Q _34345_/Q _19172_/X _19173_/X VGND VGND VPWR
+ VPWR _19342_/X sky130_fd_sc_hd__mux4_1
XFILLER_188_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31551_ _35984_/Q input23/X _31565_/S VGND VGND VPWR VPWR _31552_/A sky130_fd_sc_hd__mux2_1
X_19273_ _35047_/Q _34983_/Q _34919_/Q _34855_/Q _19103_/X _19104_/X VGND VGND VPWR
+ VPWR _19273_/X sky130_fd_sc_hd__mux4_1
X_16485_ _16448_/X _16483_/X _16484_/X _16453_/X VGND VGND VPWR VPWR _16485_/X sky130_fd_sc_hd__a22o_1
XFILLER_245_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18224_ _17149_/A _18222_/X _18223_/X _17152_/A VGND VGND VPWR VPWR _18224_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30502_ _23139_/X _35487_/Q _30506_/S VGND VGND VPWR VPWR _30503_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34270_ _34777_/CLK _34270_/D VGND VGND VPWR VPWR _34270_/Q sky130_fd_sc_hd__dfxtp_1
X_31482_ _31482_/A VGND VGND VPWR VPWR _35951_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33221_ _35973_/CLK _33221_/D VGND VGND VPWR VPWR _33221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18155_ _33802_/Q _33738_/Q _33674_/Q _33610_/Q _17902_/X _17903_/X VGND VGND VPWR
+ VPWR _18155_/X sky130_fd_sc_hd__mux4_1
X_30433_ _30433_/A VGND VGND VPWR VPWR _35454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_184_CLK clkbuf_leaf_66_CLK/A VGND VGND VPWR VPWR _35989_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_141_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17106_ _16994_/X _17104_/X _17105_/X _16997_/X VGND VGND VPWR VPWR _17106_/X sky130_fd_sc_hd__a22o_1
X_33152_ _36160_/CLK _33152_/D VGND VGND VPWR VPWR _33152_/Q sky130_fd_sc_hd__dfxtp_1
X_18086_ _34823_/Q _34759_/Q _34695_/Q _34631_/Q _17994_/X _17995_/X VGND VGND VPWR
+ VPWR _18086_/X sky130_fd_sc_hd__mux4_1
X_30364_ _30364_/A VGND VGND VPWR VPWR _35421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32103_ _35552_/CLK _32103_/D VGND VGND VPWR VPWR _32103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17037_ _16999_/X _17035_/X _17036_/X _17002_/X VGND VGND VPWR VPWR _17037_/X sky130_fd_sc_hd__a22o_1
X_33083_ _33083_/CLK _33083_/D VGND VGND VPWR VPWR _33083_/Q sky130_fd_sc_hd__dfxtp_1
X_30295_ _30295_/A VGND VGND VPWR VPWR _35389_/D sky130_fd_sc_hd__clkbuf_1
X_32034_ _36003_/CLK _32034_/D VGND VGND VPWR VPWR _32034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18988_ _18743_/X _18986_/X _18987_/X _18746_/X VGND VGND VPWR VPWR _18988_/X sky130_fd_sc_hd__a22o_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17939_ _33795_/Q _33731_/Q _33667_/Q _33603_/Q _17902_/X _17903_/X VGND VGND VPWR
+ VPWR _17939_/X sky130_fd_sc_hd__mux4_1
XFILLER_227_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33985_ _34305_/CLK _33985_/D VGND VGND VPWR VPWR _33985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35724_ _35853_/CLK _35724_/D VGND VGND VPWR VPWR _35724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20950_ _22362_/A VGND VGND VPWR VPWR _20950_/X sky130_fd_sc_hd__buf_4
X_32936_ _36075_/CLK _32936_/D VGND VGND VPWR VPWR _32936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19609_ _32497_/Q _32369_/Q _32049_/Q _36017_/Q _19576_/X _19364_/X VGND VGND VPWR
+ VPWR _19609_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35655_ _35848_/CLK _35655_/D VGND VGND VPWR VPWR _35655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20881_ _20614_/X _20879_/X _20880_/X _20623_/X VGND VGND VPWR VPWR _20881_/X sky130_fd_sc_hd__a22o_1
X_32867_ _32994_/CLK _32867_/D VGND VGND VPWR VPWR _32867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22620_ _35781_/Q _35141_/Q _34501_/Q _33861_/Q _22446_/X _22447_/X VGND VGND VPWR
+ VPWR _22620_/X sky130_fd_sc_hd__mux4_1
XFILLER_198_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34606_ _35304_/CLK _34606_/D VGND VGND VPWR VPWR _34606_/Q sky130_fd_sc_hd__dfxtp_1
X_31818_ _31818_/A VGND VGND VPWR VPWR _36110_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35586_ _35909_/CLK _35586_/D VGND VGND VPWR VPWR _35586_/Q sky130_fd_sc_hd__dfxtp_1
X_32798_ _35481_/CLK _32798_/D VGND VGND VPWR VPWR _32798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22551_ _22369_/X _22549_/X _22550_/X _22373_/X VGND VGND VPWR VPWR _22551_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34537_ _35944_/CLK _34537_/D VGND VGND VPWR VPWR _34537_/Q sky130_fd_sc_hd__dfxtp_1
X_31749_ _36078_/Q input26/X _31763_/S VGND VGND VPWR VPWR _31750_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21502_ _21496_/X _21501_/X _21394_/X VGND VGND VPWR VPWR _21510_/C sky130_fd_sc_hd__o21ba_1
X_25270_ _25109_/X _33076_/Q _25272_/S VGND VGND VPWR VPWR _25271_/A sky130_fd_sc_hd__mux2_1
X_22482_ _33025_/Q _32961_/Q _32897_/Q _32833_/Q _22295_/X _22296_/X VGND VGND VPWR
+ VPWR _22482_/X sky130_fd_sc_hd__mux4_1
XFILLER_167_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34468_ _35941_/CLK _34468_/D VGND VGND VPWR VPWR _34468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36207_ _36211_/CLK _36207_/D VGND VGND VPWR VPWR _36207_/Q sky130_fd_sc_hd__dfxtp_1
X_24221_ _24221_/A VGND VGND VPWR VPWR _32642_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33419_ _33548_/CLK _33419_/D VGND VGND VPWR VPWR _33419_/Q sky130_fd_sc_hd__dfxtp_1
X_21433_ _34787_/Q _34723_/Q _34659_/Q _34595_/Q _21182_/X _21183_/X VGND VGND VPWR
+ VPWR _21433_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_175_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _35984_/CLK sky130_fd_sc_hd__clkbuf_16
X_34399_ _35039_/CLK _34399_/D VGND VGND VPWR VPWR _34399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21364_ _21360_/X _21363_/X _21055_/X VGND VGND VPWR VPWR _21365_/D sky130_fd_sc_hd__o21ba_1
X_24152_ _24242_/S VGND VGND VPWR VPWR _24171_/S sky130_fd_sc_hd__buf_4
X_36138_ _36139_/CLK _36138_/D VGND VGND VPWR VPWR _36138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23103_ _32147_/Q _23102_/X _23115_/S VGND VGND VPWR VPWR _23104_/A sky130_fd_sc_hd__mux2_1
X_20315_ _32517_/Q _32389_/Q _32069_/Q _36037_/Q _20282_/X _20070_/X VGND VGND VPWR
+ VPWR _20315_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24083_ _24083_/A VGND VGND VPWR VPWR _32577_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28960_ _28960_/A VGND VGND VPWR VPWR _34787_/D sky130_fd_sc_hd__clkbuf_1
X_36069_ _36069_/CLK _36069_/D VGND VGND VPWR VPWR _36069_/Q sky130_fd_sc_hd__dfxtp_1
X_21295_ _33760_/Q _33696_/Q _33632_/Q _33568_/Q _21090_/X _21091_/X VGND VGND VPWR
+ VPWR _21295_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20246_ _32771_/Q _32707_/Q _32643_/Q _36099_/Q _19925_/X _20062_/X VGND VGND VPWR
+ VPWR _20246_/X sky130_fd_sc_hd__mux4_1
X_23034_ input46/X VGND VGND VPWR VPWR _23034_/X sky130_fd_sc_hd__clkbuf_4
X_27911_ _27911_/A VGND VGND VPWR VPWR _34290_/D sky130_fd_sc_hd__clkbuf_1
X_28891_ _26987_/X _34755_/Q _28903_/S VGND VGND VPWR VPWR _28892_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_1053 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27842_ _27842_/A VGND VGND VPWR VPWR _34257_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20177_ _20173_/X _20176_/X _20134_/X VGND VGND VPWR VPWR _20199_/A sky130_fd_sc_hd__o21ba_1
XTAP_5115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27773_ _34225_/Q _24354_/X _27781_/S VGND VGND VPWR VPWR _27774_/A sky130_fd_sc_hd__mux2_1
X_24985_ _23071_/X _32972_/Q _24987_/S VGND VGND VPWR VPWR _24986_/A sky130_fd_sc_hd__mux2_1
XTAP_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29512_ _29512_/A VGND VGND VPWR VPWR _35018_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26724_ _26724_/A VGND VGND VPWR VPWR _33759_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23936_ _23936_/A VGND VGND VPWR VPWR _32508_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_702 _22447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29443_ _29443_/A VGND VGND VPWR VPWR _34985_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26655_ _26655_/A VGND VGND VPWR VPWR _33727_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_713 _22465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23867_ _23867_/A VGND VGND VPWR VPWR _32475_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_724 _21759_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_735 _21223_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_746 _22283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25606_ _33231_/Q _24249_/X _25622_/S VGND VGND VPWR VPWR _25607_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29374_ _23333_/X _34953_/Q _29374_/S VGND VGND VPWR VPWR _29375_/A sky130_fd_sc_hd__mux2_1
XANTENNA_757 _22470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22818_ _33548_/Q _33484_/Q _33420_/Q _33356_/Q _20633_/X _20635_/X VGND VGND VPWR
+ VPWR _22818_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26586_ _26586_/A VGND VGND VPWR VPWR _33694_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_768 _22538_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23798_ _23798_/A VGND VGND VPWR VPWR _32443_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_779 _22604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28325_ _28325_/A VGND VGND VPWR VPWR _34486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25537_ _33200_/Q _24351_/X _25547_/S VGND VGND VPWR VPWR _25538_/A sky130_fd_sc_hd__mux2_1
X_22749_ _34569_/Q _32457_/Q _34441_/Q _34377_/Q _22531_/X _22532_/X VGND VGND VPWR
+ VPWR _22749_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16270_ _16270_/A _16270_/B _16270_/C _16270_/D VGND VGND VPWR VPWR _16271_/A sky130_fd_sc_hd__or4_4
X_28256_ _34454_/Q _24270_/X _28258_/S VGND VGND VPWR VPWR _28257_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25468_ _33167_/Q _24249_/X _25484_/S VGND VGND VPWR VPWR _25469_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_52__f_CLK clkbuf_5_26_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_52__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_27207_ _27207_/A VGND VGND VPWR VPWR _33957_/D sky130_fd_sc_hd__clkbuf_1
X_24419_ input52/X VGND VGND VPWR VPWR _24419_/X sky130_fd_sc_hd__buf_6
XFILLER_200_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_166_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _35978_/CLK sky130_fd_sc_hd__clkbuf_16
X_28187_ _28187_/A VGND VGND VPWR VPWR _34421_/D sky130_fd_sc_hd__clkbuf_1
X_25399_ _25399_/A VGND VGND VPWR VPWR _33136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27138_ _26993_/X _33925_/Q _27146_/S VGND VGND VPWR VPWR _27139_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19960_ _33275_/Q _36155_/Q _33147_/Q _33083_/Q _19711_/X _19712_/X VGND VGND VPWR
+ VPWR _19960_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27069_ _26891_/X _33892_/Q _27083_/S VGND VGND VPWR VPWR _27070_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18911_ _18588_/X _18909_/X _18910_/X _18591_/X VGND VGND VPWR VPWR _18911_/X sky130_fd_sc_hd__a22o_1
XTAP_7040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30080_ _30080_/A VGND VGND VPWR VPWR _35287_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19891_ _19855_/X _19889_/X _19890_/X _19858_/X VGND VGND VPWR VPWR _19891_/X sky130_fd_sc_hd__a22o_1
XTAP_7062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1101 _17368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1112 _32127_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1123 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18842_ _35739_/Q _35099_/Q _34459_/Q _33819_/Q _18734_/X _18735_/X VGND VGND VPWR
+ VPWR _18842_/X sky130_fd_sc_hd__mux4_1
XTAP_7095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1134 _17911_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1145 _19449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1156 _22503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1167 _22595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1178 _21099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15985_ input67/X input68/X VGND VGND VPWR VPWR _17767_/A sky130_fd_sc_hd__nor2_4
X_18773_ _35801_/Q _32176_/Q _35673_/Q _35609_/Q _18554_/X _18555_/X VGND VGND VPWR
+ VPWR _18773_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1189 _22508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17724_ _17548_/X _17722_/X _17723_/X _17553_/X VGND VGND VPWR VPWR _17724_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30982_ _30982_/A VGND VGND VPWR VPWR _35714_/D sky130_fd_sc_hd__clkbuf_1
X_33770_ _34281_/CLK _33770_/D VGND VGND VPWR VPWR _33770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32721_ _36050_/CLK _32721_/D VGND VGND VPWR VPWR _32721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17655_ _33531_/Q _33467_/Q _33403_/Q _33339_/Q _17476_/X _17477_/X VGND VGND VPWR
+ VPWR _17655_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_1249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35440_ _36013_/CLK _35440_/D VGND VGND VPWR VPWR _35440_/Q sky130_fd_sc_hd__dfxtp_1
X_16606_ _16602_/X _16605_/X _16430_/X _16431_/X VGND VGND VPWR VPWR _16623_/B sky130_fd_sc_hd__o211a_1
X_32652_ _36109_/CLK _32652_/D VGND VGND VPWR VPWR _32652_/Q sky130_fd_sc_hd__dfxtp_1
X_17586_ _33785_/Q _33721_/Q _33657_/Q _33593_/Q _17549_/X _17550_/X VGND VGND VPWR
+ VPWR _17586_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16537_ _32475_/Q _32347_/Q _32027_/Q _35995_/Q _16217_/X _16358_/X VGND VGND VPWR
+ VPWR _16537_/X sky130_fd_sc_hd__mux4_1
X_31603_ _36009_/Q input20/X _31607_/S VGND VGND VPWR VPWR _31604_/A sky130_fd_sc_hd__mux2_1
X_19325_ _32745_/Q _32681_/Q _32617_/Q _36073_/Q _19219_/X _19003_/X VGND VGND VPWR
+ VPWR _19325_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32583_ _36168_/CLK _32583_/D VGND VGND VPWR VPWR _32583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35371_ _35819_/CLK _35371_/D VGND VGND VPWR VPWR _35371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34322_ _35028_/CLK _34322_/D VGND VGND VPWR VPWR _34322_/Q sky130_fd_sc_hd__dfxtp_1
X_31534_ _31534_/A VGND VGND VPWR VPWR _35976_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16468_ _16349_/X _16466_/X _16467_/X _16355_/X VGND VGND VPWR VPWR _16468_/X sky130_fd_sc_hd__a22o_1
X_19256_ _32487_/Q _32359_/Q _32039_/Q _36007_/Q _19223_/X _19011_/X VGND VGND VPWR
+ VPWR _19256_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18207_ _35339_/Q _35275_/Q _35211_/Q _32331_/Q _16088_/X _16090_/X VGND VGND VPWR
+ VPWR _18207_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_157_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _35273_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_223_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34253_ _34317_/CLK _34253_/D VGND VGND VPWR VPWR _34253_/Q sky130_fd_sc_hd__dfxtp_1
X_31465_ _31465_/A VGND VGND VPWR VPWR _35943_/D sky130_fd_sc_hd__clkbuf_1
X_19187_ _32741_/Q _32677_/Q _32613_/Q _36069_/Q _18866_/X _19003_/X VGND VGND VPWR
+ VPWR _19187_/X sky130_fd_sc_hd__mux4_1
X_16399_ _35735_/Q _35095_/Q _34455_/Q _33815_/Q _16049_/X _16051_/X VGND VGND VPWR
+ VPWR _16399_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18138_ _18134_/X _18137_/X _17842_/X _17843_/X VGND VGND VPWR VPWR _18153_/B sky130_fd_sc_hd__o211a_1
X_33204_ _35956_/CLK _33204_/D VGND VGND VPWR VPWR _33204_/Q sky130_fd_sc_hd__dfxtp_1
X_30416_ _23270_/X _35446_/Q _30434_/S VGND VGND VPWR VPWR _30417_/A sky130_fd_sc_hd__mux2_1
X_34184_ _34312_/CLK _34184_/D VGND VGND VPWR VPWR _34184_/Q sky130_fd_sc_hd__dfxtp_1
X_31396_ _35911_/Q input53/X _31400_/S VGND VGND VPWR VPWR _31397_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18069_ _34055_/Q _33991_/Q _33927_/Q _32263_/Q _16058_/X _16060_/X VGND VGND VPWR
+ VPWR _18069_/X sky130_fd_sc_hd__mux4_1
X_30347_ _30347_/A VGND VGND VPWR VPWR _35413_/D sky130_fd_sc_hd__clkbuf_1
X_33135_ _36081_/CLK _33135_/D VGND VGND VPWR VPWR _33135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20100_ _34047_/Q _33983_/Q _33919_/Q _32255_/Q _20026_/X _20027_/X VGND VGND VPWR
+ VPWR _20100_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21080_ _34777_/Q _34713_/Q _34649_/Q _34585_/Q _20829_/X _20830_/X VGND VGND VPWR
+ VPWR _21080_/X sky130_fd_sc_hd__mux4_1
X_33066_ _36139_/CLK _33066_/D VGND VGND VPWR VPWR _33066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30278_ _30278_/A VGND VGND VPWR VPWR _35381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_1042 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32017_ _36049_/CLK _32017_/D VGND VGND VPWR VPWR _32017_/Q sky130_fd_sc_hd__dfxtp_1
X_20031_ _32765_/Q _32701_/Q _32637_/Q _36093_/Q _19925_/X _19709_/X VGND VGND VPWR
+ VPWR _20031_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24770_ _24770_/A VGND VGND VPWR VPWR _32869_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33968_ _34286_/CLK _33968_/D VGND VGND VPWR VPWR _33968_/Q sky130_fd_sc_hd__dfxtp_1
X_21982_ _33011_/Q _32947_/Q _32883_/Q _32819_/Q _21942_/X _21943_/X VGND VGND VPWR
+ VPWR _21982_/X sky130_fd_sc_hd__mux4_1
XFILLER_187_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23721_ _22907_/X _32407_/Q _23721_/S VGND VGND VPWR VPWR _23722_/A sky130_fd_sc_hd__mux2_1
X_35707_ _35707_/CLK _35707_/D VGND VGND VPWR VPWR _35707_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20933_ _34773_/Q _34709_/Q _34645_/Q _34581_/Q _20829_/X _20830_/X VGND VGND VPWR
+ VPWR _20933_/X sky130_fd_sc_hd__mux4_1
X_32919_ _35991_/CLK _32919_/D VGND VGND VPWR VPWR _32919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33899_ _36136_/CLK _33899_/D VGND VGND VPWR VPWR _33899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26440_ _26440_/A VGND VGND VPWR VPWR _33625_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23652_ _23652_/A VGND VGND VPWR VPWR _32375_/D sky130_fd_sc_hd__clkbuf_1
X_35638_ _35638_/CLK _35638_/D VGND VGND VPWR VPWR _35638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20864_ _35283_/Q _35219_/Q _35155_/Q _32275_/Q _20679_/X _20681_/X VGND VGND VPWR
+ VPWR _20864_/X sky130_fd_sc_hd__mux4_1
XFILLER_126_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22603_ _22603_/A _22603_/B _22603_/C _22603_/D VGND VGND VPWR VPWR _22604_/A sky130_fd_sc_hd__or4_4
X_26371_ _25125_/X _33593_/Q _26383_/S VGND VGND VPWR VPWR _26372_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23583_ _32343_/Q _23114_/X _23583_/S VGND VGND VPWR VPWR _23584_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_396_CLK clkbuf_6_34__f_CLK/X VGND VGND VPWR VPWR _35885_/CLK sky130_fd_sc_hd__clkbuf_16
X_35569_ _35953_/CLK _35569_/D VGND VGND VPWR VPWR _35569_/Q sky130_fd_sc_hd__dfxtp_1
X_20795_ _20656_/X _20793_/X _20794_/X _20668_/X VGND VGND VPWR VPWR _20795_/X sky130_fd_sc_hd__a22o_1
XFILLER_169_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28110_ _28110_/A VGND VGND VPWR VPWR _34384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25322_ _25186_/X _33101_/Q _25322_/S VGND VGND VPWR VPWR _25323_/A sky130_fd_sc_hd__mux2_1
X_22534_ _35074_/Q _35010_/Q _34946_/Q _34882_/Q _22462_/X _22463_/X VGND VGND VPWR
+ VPWR _22534_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29090_ _34842_/Q _29089_/X _29111_/S VGND VGND VPWR VPWR _29091_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28041_ _26928_/X _34352_/Q _28051_/S VGND VGND VPWR VPWR _28042_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25253_ _25322_/S VGND VGND VPWR VPWR _25272_/S sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_148_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _35338_/CLK sky130_fd_sc_hd__clkbuf_16
X_22465_ _22465_/A VGND VGND VPWR VPWR _22465_/X sky130_fd_sc_hd__buf_4
XFILLER_183_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24204_ _24204_/A VGND VGND VPWR VPWR _32634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21416_ _34019_/Q _33955_/Q _33891_/Q _32163_/Q _21267_/X _21268_/X VGND VGND VPWR
+ VPWR _21416_/X sky130_fd_sc_hd__mux4_1
X_25184_ _25183_/X _33036_/Q _25187_/S VGND VGND VPWR VPWR _25185_/A sky130_fd_sc_hd__mux2_1
X_22396_ _22396_/A VGND VGND VPWR VPWR _22396_/X sky130_fd_sc_hd__buf_4
XFILLER_108_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24135_ _24135_/A VGND VGND VPWR VPWR _32601_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21347_ _32481_/Q _32353_/Q _32033_/Q _36001_/Q _21170_/X _21311_/X VGND VGND VPWR
+ VPWR _21347_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29992_ _29992_/A VGND VGND VPWR VPWR _35245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24066_ _24066_/A VGND VGND VPWR VPWR _32569_/D sky130_fd_sc_hd__clkbuf_1
X_28943_ _28943_/A VGND VGND VPWR VPWR _34779_/D sky130_fd_sc_hd__clkbuf_1
X_21278_ _21274_/X _21277_/X _21030_/X _21031_/X VGND VGND VPWR VPWR _21293_/B sky130_fd_sc_hd__o211a_1
XFILLER_78_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23017_ _23016_/X _32058_/Q _23032_/S VGND VGND VPWR VPWR _23018_/A sky130_fd_sc_hd__mux2_1
X_20229_ _35330_/Q _35266_/Q _35202_/Q _32322_/Q _20012_/X _20013_/X VGND VGND VPWR
+ VPWR _20229_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_320_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _35575_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_235_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28874_ _26962_/X _34747_/Q _28882_/S VGND VGND VPWR VPWR _28875_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27825_ _34250_/Q _24431_/X _27831_/S VGND VGND VPWR VPWR _27826_/A sky130_fd_sc_hd__mux2_1
XTAP_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24968_ _24968_/A VGND VGND VPWR VPWR _32963_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27756_ _34217_/Q _24329_/X _27760_/S VGND VGND VPWR VPWR _27757_/A sky130_fd_sc_hd__mux2_1
XTAP_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26707_ _26707_/A VGND VGND VPWR VPWR _33751_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23919_ _23919_/A VGND VGND VPWR VPWR _32500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27687_ _27687_/A VGND VGND VPWR VPWR _34184_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_510 _17938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24899_ _24899_/A VGND VGND VPWR VPWR _32930_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_521 _17970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _17440_/A VGND VGND VPWR VPWR _31988_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_532 _20203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29426_ _29426_/A VGND VGND VPWR VPWR _34977_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26638_ _25119_/X _33719_/Q _26654_/S VGND VGND VPWR VPWR _26639_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_543 _20134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_554 _20143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_565 _20147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_576 _20165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_587 _19454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17371_ _17195_/X _17369_/X _17370_/X _17200_/X VGND VGND VPWR VPWR _17371_/X sky130_fd_sc_hd__a22o_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26569_ _26569_/A VGND VGND VPWR VPWR _33686_/D sky130_fd_sc_hd__clkbuf_1
X_29357_ _29357_/A VGND VGND VPWR VPWR _34944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_387_CLK clkbuf_6_41__f_CLK/X VGND VGND VPWR VPWR _34997_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_242_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_598 _20167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16322_ _32469_/Q _32341_/Q _32021_/Q _35989_/Q _16217_/X _17863_/A VGND VGND VPWR
+ VPWR _16322_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19110_ _19110_/A _19110_/B _19110_/C _19110_/D VGND VGND VPWR VPWR _19111_/A sky130_fd_sc_hd__or4_2
XFILLER_186_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28308_ _28308_/A VGND VGND VPWR VPWR _34478_/D sky130_fd_sc_hd__clkbuf_1
X_29288_ _23142_/X _34912_/Q _29290_/S VGND VGND VPWR VPWR _29289_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19041_ _34017_/Q _33953_/Q _33889_/Q _32161_/Q _18967_/X _18968_/X VGND VGND VPWR
+ VPWR _19041_/X sky130_fd_sc_hd__mux4_1
X_28239_ _28371_/S VGND VGND VPWR VPWR _28258_/S sky130_fd_sc_hd__buf_4
X_16253_ _16249_/X _16252_/X _16040_/X _16042_/X VGND VGND VPWR VPWR _16270_/B sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_139_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _35917_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31250_ _31250_/A VGND VGND VPWR VPWR _35841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16184_ _32465_/Q _32337_/Q _32017_/Q _35985_/Q _16028_/X _17863_/A VGND VGND VPWR
+ VPWR _16184_/X sky130_fd_sc_hd__mux4_1
X_30201_ _30201_/A VGND VGND VPWR VPWR _35344_/D sky130_fd_sc_hd__clkbuf_1
Xoutput208 _36233_/Q VGND VGND VPWR VPWR D2[59] sky130_fd_sc_hd__buf_2
XFILLER_177_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31181_ _35809_/Q input11/X _31181_/S VGND VGND VPWR VPWR _31182_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput219 _32088_/Q VGND VGND VPWR VPWR D3[10] sky130_fd_sc_hd__buf_2
XFILLER_173_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30132_ _35312_/Q _29157_/X _30142_/S VGND VGND VPWR VPWR _30133_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19943_ _34810_/Q _34746_/Q _34682_/Q _34618_/Q _19941_/X _19942_/X VGND VGND VPWR
+ VPWR _19943_/X sky130_fd_sc_hd__mux4_1
X_30063_ _35279_/Q _29055_/X _30079_/S VGND VGND VPWR VPWR _30064_/A sky130_fd_sc_hd__mux2_1
X_34940_ _35515_/CLK _34940_/D VGND VGND VPWR VPWR _34940_/Q sky130_fd_sc_hd__dfxtp_1
X_19874_ _19870_/X _19873_/X _19800_/X VGND VGND VPWR VPWR _19884_/C sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_311_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _35319_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18825_ _18825_/A _18825_/B _18825_/C _18825_/D VGND VGND VPWR VPWR _18826_/A sky130_fd_sc_hd__or4_2
XTAP_6180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34871_ _35257_/CLK _34871_/D VGND VGND VPWR VPWR _34871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33822_ _35743_/CLK _33822_/D VGND VGND VPWR VPWR _33822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18756_ _18747_/X _18754_/X _18755_/X VGND VGND VPWR VPWR _18757_/D sky130_fd_sc_hd__o21ba_1
XTAP_5490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17707_ _33212_/Q _32572_/Q _35964_/Q _35900_/Q _17427_/X _17428_/X VGND VGND VPWR
+ VPWR _17707_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33753_ _35799_/CLK _33753_/D VGND VGND VPWR VPWR _33753_/Q sky130_fd_sc_hd__dfxtp_1
X_18687_ _33495_/Q _33431_/Q _33367_/Q _33303_/Q _18298_/X _18299_/X VGND VGND VPWR
+ VPWR _18687_/X sky130_fd_sc_hd__mux4_1
X_30965_ _30965_/A VGND VGND VPWR VPWR _35706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32704_ _36098_/CLK _32704_/D VGND VGND VPWR VPWR _32704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17638_ _33210_/Q _32570_/Q _35962_/Q _35898_/Q _17427_/X _17428_/X VGND VGND VPWR
+ VPWR _17638_/X sky130_fd_sc_hd__mux4_1
X_33684_ _33685_/CLK _33684_/D VGND VGND VPWR VPWR _33684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30896_ _30896_/A VGND VGND VPWR VPWR _35673_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35423_ _35744_/CLK _35423_/D VGND VGND VPWR VPWR _35423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32635_ _33083_/CLK _32635_/D VGND VGND VPWR VPWR _32635_/Q sky130_fd_sc_hd__dfxtp_1
X_17569_ _35768_/Q _35128_/Q _34488_/Q _33848_/Q _17493_/X _17494_/X VGND VGND VPWR
+ VPWR _17569_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_378_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _35952_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19308_ _35304_/Q _35240_/Q _35176_/Q _32296_/Q _19306_/X _19307_/X VGND VGND VPWR
+ VPWR _19308_/X sky130_fd_sc_hd__mux4_1
X_20580_ _22502_/A VGND VGND VPWR VPWR _20580_/X sky130_fd_sc_hd__buf_8
XFILLER_177_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35354_ _35929_/CLK _35354_/D VGND VGND VPWR VPWR _35354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32566_ _36022_/CLK _32566_/D VGND VGND VPWR VPWR _32566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34305_ _34305_/CLK _34305_/D VGND VGND VPWR VPWR _34305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_917 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31517_ _23303_/X _35968_/Q _31535_/S VGND VGND VPWR VPWR _31518_/A sky130_fd_sc_hd__mux2_1
X_19239_ _19096_/X _19237_/X _19238_/X _19099_/X VGND VGND VPWR VPWR _19239_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35285_ _36191_/CLK _35285_/D VGND VGND VPWR VPWR _35285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32497_ _36078_/CLK _32497_/D VGND VGND VPWR VPWR _32497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34236_ _36157_/CLK _34236_/D VGND VGND VPWR VPWR _34236_/Q sky130_fd_sc_hd__dfxtp_1
X_22250_ _22250_/A _22250_/B _22250_/C _22250_/D VGND VGND VPWR VPWR _22251_/A sky130_fd_sc_hd__or4_4
X_31448_ _31448_/A VGND VGND VPWR VPWR _35935_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21201_ _33245_/Q _36125_/Q _33117_/Q _33053_/Q _20952_/X _20953_/X VGND VGND VPWR
+ VPWR _21201_/X sky130_fd_sc_hd__mux4_1
X_22181_ _35064_/Q _35000_/Q _34936_/Q _34872_/Q _22109_/X _22110_/X VGND VGND VPWR
+ VPWR _22181_/X sky130_fd_sc_hd__mux4_1
X_31379_ _35903_/Q input44/X _31379_/S VGND VGND VPWR VPWR _31380_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34167_ _34295_/CLK _34167_/D VGND VGND VPWR VPWR _34167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21132_ _21096_/X _21130_/X _21131_/X _21099_/X VGND VGND VPWR VPWR _21132_/X sky130_fd_sc_hd__a22o_1
X_33118_ _36127_/CLK _33118_/D VGND VGND VPWR VPWR _33118_/Q sky130_fd_sc_hd__dfxtp_1
X_34098_ _34286_/CLK _34098_/D VGND VGND VPWR VPWR _34098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21063_ _34009_/Q _33945_/Q _33881_/Q _32153_/Q _20914_/X _20915_/X VGND VGND VPWR
+ VPWR _21063_/X sky130_fd_sc_hd__mux4_1
X_25940_ _25940_/A VGND VGND VPWR VPWR _33388_/D sky130_fd_sc_hd__clkbuf_1
X_33049_ _35863_/CLK _33049_/D VGND VGND VPWR VPWR _33049_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_302_CLK clkbuf_6_50__f_CLK/X VGND VGND VPWR VPWR _35771_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20014_ _35324_/Q _35260_/Q _35196_/Q _32316_/Q _20012_/X _20013_/X VGND VGND VPWR
+ VPWR _20014_/X sky130_fd_sc_hd__mux4_1
XFILLER_115_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25871_ _25871_/A VGND VGND VPWR VPWR _33356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24822_ _24822_/A VGND VGND VPWR VPWR _32894_/D sky130_fd_sc_hd__clkbuf_1
X_27610_ _27610_/A VGND VGND VPWR VPWR _34147_/D sky130_fd_sc_hd__clkbuf_1
X_28590_ _28590_/A VGND VGND VPWR VPWR _34612_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27541_ _26990_/X _34116_/Q _27551_/S VGND VGND VPWR VPWR _27542_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24753_ _24753_/A VGND VGND VPWR VPWR _32861_/D sky130_fd_sc_hd__clkbuf_1
X_21965_ _21754_/X _21963_/X _21964_/X _21759_/X VGND VGND VPWR VPWR _21965_/X sky130_fd_sc_hd__a22o_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23704_ _23704_/A VGND VGND VPWR VPWR _32398_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ _34005_/Q _33941_/Q _33877_/Q _32149_/Q _20914_/X _20915_/X VGND VGND VPWR
+ VPWR _20916_/X sky130_fd_sc_hd__mux4_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27472_ _26888_/X _34083_/Q _27488_/S VGND VGND VPWR VPWR _27473_/A sky130_fd_sc_hd__mux2_1
X_24684_ _23028_/X _32830_/Q _24686_/S VGND VGND VPWR VPWR _24685_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21896_ _21892_/X _21895_/X _21761_/X VGND VGND VPWR VPWR _21897_/D sky130_fd_sc_hd__o21ba_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26423_ _26423_/A VGND VGND VPWR VPWR _33617_/D sky130_fd_sc_hd__clkbuf_1
X_29211_ _34881_/Q _29210_/X _29235_/S VGND VGND VPWR VPWR _29212_/A sky130_fd_sc_hd__mux2_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23635_ _23635_/A VGND VGND VPWR VPWR _32367_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20847_ _32723_/Q _32659_/Q _32595_/Q _36051_/Q _20813_/X _22313_/A VGND VGND VPWR
+ VPWR _20847_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_369_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _36081_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_243_1433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29142_ _34859_/Q _29141_/X _29142_/S VGND VGND VPWR VPWR _29143_/A sky130_fd_sc_hd__mux2_1
X_26354_ _25100_/X _33585_/Q _26362_/S VGND VGND VPWR VPWR _26355_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23566_ _23566_/A VGND VGND VPWR VPWR _32334_/D sky130_fd_sc_hd__clkbuf_1
X_20778_ _34001_/Q _33937_/Q _33873_/Q _32145_/Q _20708_/X _20709_/X VGND VGND VPWR
+ VPWR _20778_/X sky130_fd_sc_hd__mux4_1
X_25305_ _25305_/A VGND VGND VPWR VPWR _33092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22517_ _32514_/Q _32386_/Q _32066_/Q _36034_/Q _22229_/X _22370_/X VGND VGND VPWR
+ VPWR _22517_/X sky130_fd_sc_hd__mux4_1
X_29073_ input62/X VGND VGND VPWR VPWR _29073_/X sky130_fd_sc_hd__buf_4
XFILLER_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26285_ _24998_/X _33552_/Q _26299_/S VGND VGND VPWR VPWR _26286_/A sky130_fd_sc_hd__mux2_1
X_23497_ _22982_/X _32303_/Q _23509_/S VGND VGND VPWR VPWR _23498_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28024_ _26903_/X _34344_/Q _28030_/S VGND VGND VPWR VPWR _28025_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25236_ _25236_/A VGND VGND VPWR VPWR _33059_/D sky130_fd_sc_hd__clkbuf_1
X_22448_ _35776_/Q _35136_/Q _34496_/Q _33856_/Q _22446_/X _22447_/X VGND VGND VPWR
+ VPWR _22448_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25167_ _25167_/A VGND VGND VPWR VPWR _33030_/D sky130_fd_sc_hd__clkbuf_1
X_22379_ _35582_/Q _35518_/Q _35454_/Q _35390_/Q _22203_/X _22204_/X VGND VGND VPWR
+ VPWR _22379_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24118_ _24118_/A VGND VGND VPWR VPWR _32593_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25098_ _25097_/X _33008_/Q _25113_/S VGND VGND VPWR VPWR _25099_/A sky130_fd_sc_hd__mux2_1
X_29975_ _29975_/A VGND VGND VPWR VPWR _35237_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28926_ _28926_/A VGND VGND VPWR VPWR _34771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24049_ _24049_/A VGND VGND VPWR VPWR _32561_/D sky130_fd_sc_hd__clkbuf_1
X_16940_ _34534_/Q _32422_/Q _34406_/Q _34342_/Q _16872_/X _16873_/X VGND VGND VPWR
+ VPWR _16940_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16871_ _16796_/X _16869_/X _16870_/X _16799_/X VGND VGND VPWR VPWR _16871_/X sky130_fd_sc_hd__a22o_1
X_28857_ _26937_/X _34739_/Q _28861_/S VGND VGND VPWR VPWR _28858_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18610_ _33749_/Q _33685_/Q _33621_/Q _33557_/Q _18437_/X _18438_/X VGND VGND VPWR
+ VPWR _18610_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27808_ _27808_/A VGND VGND VPWR VPWR _34241_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19590_ _34800_/Q _34736_/Q _34672_/Q _34608_/Q _19588_/X _19589_/X VGND VGND VPWR
+ VPWR _19590_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28788_ _26835_/X _34706_/Q _28798_/S VGND VGND VPWR VPWR _28789_/A sky130_fd_sc_hd__mux2_1
XTAP_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18541_ _34259_/Q _34195_/Q _34131_/Q _34067_/Q _18305_/X _18307_/X VGND VGND VPWR
+ VPWR _18541_/X sky130_fd_sc_hd__mux4_1
XTAP_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27739_ _34209_/Q _24304_/X _27739_/S VGND VGND VPWR VPWR _27740_/A sky130_fd_sc_hd__mux2_1
XTAP_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18472_ _18472_/A _18472_/B _18472_/C _18472_/D VGND VGND VPWR VPWR _18473_/A sky130_fd_sc_hd__or4_4
X_30750_ _30750_/A VGND VGND VPWR VPWR _35604_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_340 _36205_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_351 _36206_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_362 _36207_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29409_ _23121_/X _34969_/Q _29425_/S VGND VGND VPWR VPWR _29410_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17423_ _35828_/Q _32206_/Q _35700_/Q _35636_/Q _17313_/X _17314_/X VGND VGND VPWR
+ VPWR _17423_/X sky130_fd_sc_hd__mux4_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_373 _36208_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30681_ _35572_/Q _29169_/X _30683_/S VGND VGND VPWR VPWR _30682_/A sky130_fd_sc_hd__mux2_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_384 _36209_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_395 _36210_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32420_ _35239_/CLK _32420_/D VGND VGND VPWR VPWR _32420_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _33202_/Q _32562_/Q _35954_/Q _35890_/Q _17074_/X _17075_/X VGND VGND VPWR
+ VPWR _17354_/X sky130_fd_sc_hd__mux4_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16305_ _35028_/Q _34964_/Q _34900_/Q _34836_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _16305_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17285_ _33200_/Q _32560_/Q _35952_/Q _35888_/Q _17074_/X _17075_/X VGND VGND VPWR
+ VPWR _17285_/X sky130_fd_sc_hd__mux4_1
X_32351_ _36129_/CLK _32351_/D VGND VGND VPWR VPWR _32351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16236_ _16087_/X _16234_/X _16235_/X _16097_/X VGND VGND VPWR VPWR _16236_/X sky130_fd_sc_hd__a22o_1
X_19024_ _18946_/X _19020_/X _19023_/X _18949_/X VGND VGND VPWR VPWR _19024_/X sky130_fd_sc_hd__a22o_1
X_31302_ _35866_/Q input4/X _31316_/S VGND VGND VPWR VPWR _31303_/A sky130_fd_sc_hd__mux2_1
X_35070_ _35326_/CLK _35070_/D VGND VGND VPWR VPWR _35070_/Q sky130_fd_sc_hd__dfxtp_1
X_32282_ _35226_/CLK _32282_/D VGND VGND VPWR VPWR _32282_/Q sky130_fd_sc_hd__dfxtp_1
X_31233_ _31233_/A VGND VGND VPWR VPWR _35833_/D sky130_fd_sc_hd__clkbuf_1
X_34021_ _34087_/CLK _34021_/D VGND VGND VPWR VPWR _34021_/Q sky130_fd_sc_hd__dfxtp_1
X_16167_ _16873_/A VGND VGND VPWR VPWR _16167_/X sky130_fd_sc_hd__buf_6
XFILLER_154_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31164_ _31164_/A VGND VGND VPWR VPWR _35800_/D sky130_fd_sc_hd__clkbuf_1
X_16098_ _16087_/X _16091_/X _16095_/X _16097_/X VGND VGND VPWR VPWR _16098_/X sky130_fd_sc_hd__a22o_1
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30115_ _35304_/Q _29132_/X _30121_/S VGND VGND VPWR VPWR _30116_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19926_ _32762_/Q _32698_/Q _32634_/Q _36090_/Q _19925_/X _19709_/X VGND VGND VPWR
+ VPWR _19926_/X sky130_fd_sc_hd__mux4_1
XFILLER_218_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35972_ _35973_/CLK _35972_/D VGND VGND VPWR VPWR _35972_/Q sky130_fd_sc_hd__dfxtp_1
X_31095_ _35768_/Q _29182_/X _31109_/S VGND VGND VPWR VPWR _31096_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30046_ _30046_/A VGND VGND VPWR VPWR _35271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34923_ _34987_/CLK _34923_/D VGND VGND VPWR VPWR _34923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19857_ _34040_/Q _33976_/Q _33912_/Q _32248_/Q _19673_/X _19674_/X VGND VGND VPWR
+ VPWR _19857_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18808_ _18804_/X _18807_/X _18730_/X _18731_/X VGND VGND VPWR VPWR _18825_/B sky130_fd_sc_hd__o211a_1
X_34854_ _35239_/CLK _34854_/D VGND VGND VPWR VPWR _34854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19788_ _19716_/X _19786_/X _19787_/X _19720_/X VGND VGND VPWR VPWR _19788_/X sky130_fd_sc_hd__a22o_1
XFILLER_216_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33805_ _34317_/CLK _33805_/D VGND VGND VPWR VPWR _33805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18739_ _33176_/Q _32536_/Q _35928_/Q _35864_/Q _18668_/X _18669_/X VGND VGND VPWR
+ VPWR _18739_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34785_ _35098_/CLK _34785_/D VGND VGND VPWR VPWR _34785_/Q sky130_fd_sc_hd__dfxtp_1
X_31997_ _34205_/CLK _31997_/D VGND VGND VPWR VPWR _31997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33736_ _34243_/CLK _33736_/D VGND VGND VPWR VPWR _33736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21750_ _34796_/Q _34732_/Q _34668_/Q _34604_/Q _21535_/X _21536_/X VGND VGND VPWR
+ VPWR _21750_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30948_ _30948_/A VGND VGND VPWR VPWR _35698_/D sky130_fd_sc_hd__clkbuf_1
X_20701_ _20685_/X _20698_/X _20700_/X VGND VGND VPWR VPWR _20702_/D sky130_fd_sc_hd__o21ba_1
XFILLER_145_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33667_ _33795_/CLK _33667_/D VGND VGND VPWR VPWR _33667_/Q sky130_fd_sc_hd__dfxtp_1
X_21681_ _21396_/X _21679_/X _21680_/X _21399_/X VGND VGND VPWR VPWR _21681_/X sky130_fd_sc_hd__a22o_1
XFILLER_211_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30879_ _30879_/A VGND VGND VPWR VPWR _35665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35406_ _35791_/CLK _35406_/D VGND VGND VPWR VPWR _35406_/Q sky130_fd_sc_hd__dfxtp_1
X_23420_ _23420_/A VGND VGND VPWR VPWR _32268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20632_ _20657_/A VGND VGND VPWR VPWR _22429_/A sky130_fd_sc_hd__buf_12
XFILLER_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32618_ _36139_/CLK _32618_/D VGND VGND VPWR VPWR _32618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33598_ _33729_/CLK _33598_/D VGND VGND VPWR VPWR _33598_/Q sky130_fd_sc_hd__dfxtp_1
X_35337_ _35337_/CLK _35337_/D VGND VGND VPWR VPWR _35337_/Q sky130_fd_sc_hd__dfxtp_1
X_23351_ _23351_/A VGND VGND VPWR VPWR _32235_/D sky130_fd_sc_hd__clkbuf_1
X_20563_ _33229_/Q _32589_/Q _35981_/Q _35917_/Q _18375_/X _18376_/X VGND VGND VPWR
+ VPWR _20563_/X sky130_fd_sc_hd__mux4_1
X_32549_ _35942_/CLK _32549_/D VGND VGND VPWR VPWR _32549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22302_ _35772_/Q _35132_/Q _34492_/Q _33852_/Q _22093_/X _22094_/X VGND VGND VPWR
+ VPWR _22302_/X sky130_fd_sc_hd__mux4_1
X_26070_ _26070_/A VGND VGND VPWR VPWR _33450_/D sky130_fd_sc_hd__clkbuf_1
X_35268_ _35332_/CLK _35268_/D VGND VGND VPWR VPWR _35268_/Q sky130_fd_sc_hd__dfxtp_1
X_23282_ _23282_/A VGND VGND VPWR VPWR _32211_/D sky130_fd_sc_hd__clkbuf_1
X_20494_ _19449_/A _20492_/X _20493_/X _19452_/A VGND VGND VPWR VPWR _20494_/X sky130_fd_sc_hd__a22o_1
X_25021_ _25021_/A VGND VGND VPWR VPWR _32983_/D sky130_fd_sc_hd__clkbuf_1
X_22233_ _22228_/X _22232_/X _22089_/X _22090_/X VGND VGND VPWR VPWR _22250_/B sky130_fd_sc_hd__o211a_1
X_34219_ _34282_/CLK _34219_/D VGND VGND VPWR VPWR _34219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35199_ _35581_/CLK _35199_/D VGND VGND VPWR VPWR _35199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22164_ _32504_/Q _32376_/Q _32056_/Q _36024_/Q _21876_/X _22017_/X VGND VGND VPWR
+ VPWR _22164_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21115_ _21111_/X _21114_/X _21041_/X VGND VGND VPWR VPWR _21125_/C sky130_fd_sc_hd__o21ba_1
XTAP_6938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29760_ _29787_/S VGND VGND VPWR VPWR _29779_/S sky130_fd_sc_hd__buf_4
XFILLER_120_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26972_ _26971_/X _33854_/Q _26975_/S VGND VGND VPWR VPWR _26973_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22095_ _35766_/Q _35126_/Q _34486_/Q _33846_/Q _22093_/X _22094_/X VGND VGND VPWR
+ VPWR _22095_/X sky130_fd_sc_hd__mux4_1
XTAP_6949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28711_ _28711_/A VGND VGND VPWR VPWR _34669_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25923_ _25923_/A VGND VGND VPWR VPWR _33380_/D sky130_fd_sc_hd__clkbuf_1
X_21046_ _21752_/A VGND VGND VPWR VPWR _21046_/X sky130_fd_sc_hd__clkbuf_4
X_29691_ _35103_/Q _29104_/X _29695_/S VGND VGND VPWR VPWR _29692_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28642_ _28642_/A VGND VGND VPWR VPWR _34637_/D sky130_fd_sc_hd__clkbuf_1
X_25854_ _25159_/X _33348_/Q _25864_/S VGND VGND VPWR VPWR _25855_/A sky130_fd_sc_hd__mux2_1
XFILLER_247_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24805_ _23003_/X _32886_/Q _24823_/S VGND VGND VPWR VPWR _24806_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25785_ _25057_/X _33315_/Q _25801_/S VGND VGND VPWR VPWR _25786_/A sky130_fd_sc_hd__mux2_1
X_28573_ _26915_/X _34604_/Q _28591_/S VGND VGND VPWR VPWR _28574_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22997_ input32/X VGND VGND VPWR VPWR _22997_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27524_ _26965_/X _34108_/Q _27530_/S VGND VGND VPWR VPWR _27525_/A sky130_fd_sc_hd__mux2_1
X_24736_ _24736_/A VGND VGND VPWR VPWR _32853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21948_ _35826_/Q _32203_/Q _35698_/Q _35634_/Q _21913_/X _21914_/X VGND VGND VPWR
+ VPWR _21948_/X sky130_fd_sc_hd__mux4_1
XFILLER_243_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27455_ _26863_/X _34075_/Q _27467_/S VGND VGND VPWR VPWR _27456_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24667_ _24715_/S VGND VGND VPWR VPWR _24686_/S sky130_fd_sc_hd__buf_4
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21879_ _21663_/X _21877_/X _21878_/X _21667_/X VGND VGND VPWR VPWR _21879_/X sky130_fd_sc_hd__a22o_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26406_ _25177_/X _33610_/Q _26412_/S VGND VGND VPWR VPWR _26407_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23618_ _23618_/A VGND VGND VPWR VPWR _32359_/D sky130_fd_sc_hd__clkbuf_1
X_27386_ _27386_/A VGND VGND VPWR VPWR _34042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24598_ _22901_/X _32789_/Q _24602_/S VGND VGND VPWR VPWR _24599_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26337_ _25075_/X _33577_/Q _26341_/S VGND VGND VPWR VPWR _26338_/A sky130_fd_sc_hd__mux2_1
X_29125_ _29125_/A VGND VGND VPWR VPWR _34853_/D sky130_fd_sc_hd__clkbuf_1
X_23549_ _23059_/X _32328_/Q _23551_/S VGND VGND VPWR VPWR _23550_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29056_ _34831_/Q _29055_/X _29080_/S VGND VGND VPWR VPWR _29057_/A sky130_fd_sc_hd__mux2_1
X_17070_ _35818_/Q _32195_/Q _35690_/Q _35626_/Q _16960_/X _16961_/X VGND VGND VPWR
+ VPWR _17070_/X sky130_fd_sc_hd__mux4_1
X_26268_ _26268_/A VGND VGND VPWR VPWR _33544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16021_ _17903_/A VGND VGND VPWR VPWR _16021_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25219_ _25219_/A VGND VGND VPWR VPWR _33051_/D sky130_fd_sc_hd__clkbuf_1
X_28007_ _26878_/X _34336_/Q _28009_/S VGND VGND VPWR VPWR _28008_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26199_ _26199_/A VGND VGND VPWR VPWR _33511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_70_CLK clkbuf_leaf_73_CLK/A VGND VGND VPWR VPWR _36118_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_87_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17972_ _34308_/Q _34244_/Q _34180_/Q _34116_/Q _17795_/X _17796_/X VGND VGND VPWR
+ VPWR _17972_/X sky130_fd_sc_hd__mux4_1
X_29958_ _29958_/A VGND VGND VPWR VPWR _35229_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1040 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19711_ _20282_/A VGND VGND VPWR VPWR _19711_/X sky130_fd_sc_hd__buf_4
X_28909_ _27014_/X _34764_/Q _28911_/S VGND VGND VPWR VPWR _28910_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16923_ _17982_/A VGND VGND VPWR VPWR _16923_/X sky130_fd_sc_hd__buf_6
XFILLER_104_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29889_ _35197_/Q _29197_/X _29893_/S VGND VGND VPWR VPWR _29890_/A sky130_fd_sc_hd__mux2_1
X_31920_ _31920_/A VGND VGND VPWR VPWR _36159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19642_ _20129_/A VGND VGND VPWR VPWR _19642_/X sky130_fd_sc_hd__buf_4
X_16854_ _16848_/X _16853_/X _16775_/X VGND VGND VPWR VPWR _16878_/A sky130_fd_sc_hd__o21ba_1
XFILLER_4_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19573_ _32752_/Q _32688_/Q _32624_/Q _36080_/Q _19572_/X _19356_/X VGND VGND VPWR
+ VPWR _19573_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31851_ _31851_/A VGND VGND VPWR VPWR _36126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16785_ _16779_/X _16782_/X _16783_/X _16784_/X VGND VGND VPWR VPWR _16810_/B sky130_fd_sc_hd__o211a_1
XFILLER_168_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18524_ _18344_/X _18522_/X _18523_/X _18354_/X VGND VGND VPWR VPWR _18524_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30802_ _23241_/X _35629_/Q _30818_/S VGND VGND VPWR VPWR _30803_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34570_ _35787_/CLK _34570_/D VGND VGND VPWR VPWR _34570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31782_ _36094_/Q input43/X _31784_/S VGND VGND VPWR VPWR _31783_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33521_ _34033_/CLK _33521_/D VGND VGND VPWR VPWR _33521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30733_ _35597_/Q _29246_/X _30733_/S VGND VGND VPWR VPWR _30734_/A sky130_fd_sc_hd__mux2_1
X_18455_ _18451_/X _18454_/X _18340_/X _18342_/X VGND VGND VPWR VPWR _18472_/B sky130_fd_sc_hd__o211a_2
XFILLER_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_170 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17406_ _17202_/X _17404_/X _17405_/X _17205_/X VGND VGND VPWR VPWR _17406_/X sky130_fd_sc_hd__a22o_1
X_33452_ _34293_/CLK _33452_/D VGND VGND VPWR VPWR _33452_/Q sky130_fd_sc_hd__dfxtp_1
X_18386_ _20069_/A VGND VGND VPWR VPWR _19454_/A sky130_fd_sc_hd__buf_12
X_30664_ _30733_/S VGND VGND VPWR VPWR _30683_/S sky130_fd_sc_hd__buf_6
XFILLER_57_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32403_ _36211_/CLK _32403_/D VGND VGND VPWR VPWR _32403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36171_ _36171_/CLK _36171_/D VGND VGND VPWR VPWR _36171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17337_ _17333_/X _17336_/X _17128_/X VGND VGND VPWR VPWR _17367_/A sky130_fd_sc_hd__o21ba_1
X_30595_ _30595_/A VGND VGND VPWR VPWR _35531_/D sky130_fd_sc_hd__clkbuf_1
X_33383_ _35991_/CLK _33383_/D VGND VGND VPWR VPWR _33383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35122_ _35826_/CLK _35122_/D VGND VGND VPWR VPWR _35122_/Q sky130_fd_sc_hd__dfxtp_1
X_32334_ _36041_/CLK _32334_/D VGND VGND VPWR VPWR _32334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17268_ _33520_/Q _33456_/Q _33392_/Q _33328_/Q _17123_/X _17124_/X VGND VGND VPWR
+ VPWR _17268_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19007_ _33248_/Q _36128_/Q _33120_/Q _33056_/Q _19005_/X _19006_/X VGND VGND VPWR
+ VPWR _19007_/X sky130_fd_sc_hd__mux4_1
X_16219_ _32978_/Q _32914_/Q _32850_/Q _32786_/Q _16033_/X _16035_/X VGND VGND VPWR
+ VPWR _16219_/X sky130_fd_sc_hd__mux4_1
X_35053_ _35757_/CLK _35053_/D VGND VGND VPWR VPWR _35053_/Q sky130_fd_sc_hd__dfxtp_1
X_32265_ _34816_/CLK _32265_/D VGND VGND VPWR VPWR _32265_/Q sky130_fd_sc_hd__dfxtp_1
X_17199_ _34286_/Q _34222_/Q _34158_/Q _34094_/Q _17089_/X _17090_/X VGND VGND VPWR
+ VPWR _17199_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_61_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _34278_/CLK sky130_fd_sc_hd__clkbuf_16
X_34004_ _34004_/CLK _34004_/D VGND VGND VPWR VPWR _34004_/Q sky130_fd_sc_hd__dfxtp_1
X_31216_ _31216_/A VGND VGND VPWR VPWR _35825_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32196_ _35819_/CLK _32196_/D VGND VGND VPWR VPWR _32196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31147_ _31147_/A VGND VGND VPWR VPWR _35792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19909_ _34809_/Q _34745_/Q _34681_/Q _34617_/Q _19588_/X _19589_/X VGND VGND VPWR
+ VPWR _19909_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_6_29__f_CLK clkbuf_5_14_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_29__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_216_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31078_ _35760_/Q _29157_/X _31088_/S VGND VGND VPWR VPWR _31079_/A sky130_fd_sc_hd__mux2_1
X_35955_ _35955_/CLK _35955_/D VGND VGND VPWR VPWR _35955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30029_ _30029_/A VGND VGND VPWR VPWR _35263_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34906_ _34970_/CLK _34906_/D VGND VGND VPWR VPWR _34906_/Q sky130_fd_sc_hd__dfxtp_1
X_22920_ input5/X VGND VGND VPWR VPWR _22920_/X sky130_fd_sc_hd__buf_4
XFILLER_60_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35886_ _35950_/CLK _35886_/D VGND VGND VPWR VPWR _35886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22851_ _22847_/X _22850_/X _22434_/A VGND VGND VPWR VPWR _22873_/A sky130_fd_sc_hd__o21ba_1
X_34837_ _36196_/CLK _34837_/D VGND VGND VPWR VPWR _34837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21802_ _22508_/A VGND VGND VPWR VPWR _21802_/X sky130_fd_sc_hd__clkbuf_4
X_25570_ _25597_/S VGND VGND VPWR VPWR _25589_/S sky130_fd_sc_hd__buf_4
X_22782_ _22778_/X _22781_/X _22467_/A VGND VGND VPWR VPWR _22783_/D sky130_fd_sc_hd__o21ba_1
X_34768_ _35280_/CLK _34768_/D VGND VGND VPWR VPWR _34768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24521_ _22991_/X _32754_/Q _24527_/S VGND VGND VPWR VPWR _24522_/A sky130_fd_sc_hd__mux2_1
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21733_ _32492_/Q _32364_/Q _32044_/Q _36012_/Q _21523_/X _21664_/X VGND VGND VPWR
+ VPWR _21733_/X sky130_fd_sc_hd__mux4_1
X_33719_ _34293_/CLK _33719_/D VGND VGND VPWR VPWR _33719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34699_ _35339_/CLK _34699_/D VGND VGND VPWR VPWR _34699_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27240_ _27240_/A VGND VGND VPWR VPWR _33973_/D sky130_fd_sc_hd__clkbuf_1
X_24452_ _22889_/X _32721_/Q _24464_/S VGND VGND VPWR VPWR _24453_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21664_ _22370_/A VGND VGND VPWR VPWR _21664_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_71_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23403_ _32260_/Q _23316_/X _23413_/S VGND VGND VPWR VPWR _23404_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27171_ _27171_/A VGND VGND VPWR VPWR _33940_/D sky130_fd_sc_hd__clkbuf_1
X_20615_ _20657_/A VGND VGND VPWR VPWR _22578_/A sky130_fd_sc_hd__buf_12
XFILLER_177_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24383_ _32698_/Q _24382_/X _24398_/S VGND VGND VPWR VPWR _24384_/A sky130_fd_sc_hd__mux2_1
X_21595_ _35816_/Q _32192_/Q _35688_/Q _35624_/Q _21560_/X _21561_/X VGND VGND VPWR
+ VPWR _21595_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26122_ _25156_/X _33475_/Q _26134_/S VGND VGND VPWR VPWR _26123_/A sky130_fd_sc_hd__mux2_1
X_23334_ _32229_/Q _23333_/X _23334_/S VGND VGND VPWR VPWR _23335_/A sky130_fd_sc_hd__mux2_1
X_20546_ _34317_/Q _34253_/Q _34189_/Q _34125_/Q _18345_/X _18346_/X VGND VGND VPWR
+ VPWR _20546_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26053_ _25053_/X _33442_/Q _26071_/S VGND VGND VPWR VPWR _26054_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23265_ _32206_/Q _23264_/X _23268_/S VGND VGND VPWR VPWR _23266_/A sky130_fd_sc_hd__mux2_1
X_20477_ _35338_/Q _35274_/Q _35210_/Q _32330_/Q _18388_/X _18390_/X VGND VGND VPWR
+ VPWR _20477_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_52_CLK clkbuf_leaf_57_CLK/A VGND VGND VPWR VPWR _32860_/CLK sky130_fd_sc_hd__clkbuf_16
X_25004_ input45/X VGND VGND VPWR VPWR _25004_/X sky130_fd_sc_hd__buf_4
X_22216_ _22216_/A _22216_/B _22216_/C _22216_/D VGND VGND VPWR VPWR _22217_/A sky130_fd_sc_hd__or4_4
XFILLER_118_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23196_ _23196_/A VGND VGND VPWR VPWR _32180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29812_ _35160_/Q _29082_/X _29830_/S VGND VGND VPWR VPWR _29813_/A sky130_fd_sc_hd__mux2_1
X_22147_ _22147_/A VGND VGND VPWR VPWR _36215_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29743_ _29743_/A VGND VGND VPWR VPWR _35127_/D sky130_fd_sc_hd__clkbuf_1
X_26955_ _26955_/A VGND VGND VPWR VPWR _33848_/D sky130_fd_sc_hd__clkbuf_1
X_22078_ _33526_/Q _33462_/Q _33398_/Q _33334_/Q _22076_/X _22077_/X VGND VGND VPWR
+ VPWR _22078_/X sky130_fd_sc_hd__mux4_1
XTAP_6779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21029_ _20957_/X _21027_/X _21028_/X _20961_/X VGND VGND VPWR VPWR _21029_/X sky130_fd_sc_hd__a22o_1
X_25906_ _25906_/A VGND VGND VPWR VPWR _33372_/D sky130_fd_sc_hd__clkbuf_1
X_29674_ _35095_/Q _29079_/X _29674_/S VGND VGND VPWR VPWR _29675_/A sky130_fd_sc_hd__mux2_1
X_26886_ _26884_/X _33826_/Q _26913_/S VGND VGND VPWR VPWR _26887_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28625_ _26993_/X _34629_/Q _28633_/S VGND VGND VPWR VPWR _28626_/A sky130_fd_sc_hd__mux2_1
X_25837_ _25134_/X _33340_/Q _25843_/S VGND VGND VPWR VPWR _25838_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28556_ _26891_/X _34596_/Q _28570_/S VGND VGND VPWR VPWR _28557_/A sky130_fd_sc_hd__mux2_1
X_16570_ _17982_/A VGND VGND VPWR VPWR _16570_/X sky130_fd_sc_hd__buf_6
X_25768_ _25032_/X _33307_/Q _25780_/S VGND VGND VPWR VPWR _25769_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27507_ _26940_/X _34100_/Q _27509_/S VGND VGND VPWR VPWR _27508_/A sky130_fd_sc_hd__mux2_1
X_24719_ _31815_/B _31410_/B VGND VGND VPWR VPWR _24852_/S sky130_fd_sc_hd__nand2_8
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28487_ _28487_/A VGND VGND VPWR VPWR _34563_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25699_ _25699_/A VGND VGND VPWR VPWR _33275_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18240_ _35084_/Q _35020_/Q _34956_/Q _34892_/Q _16079_/X _16081_/X VGND VGND VPWR
+ VPWR _18240_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27438_ _26838_/X _34067_/Q _27446_/S VGND VGND VPWR VPWR _27439_/A sky130_fd_sc_hd__mux2_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18171_ _15977_/X _18169_/X _18170_/X _15987_/X VGND VGND VPWR VPWR _18171_/X sky130_fd_sc_hd__a22o_1
X_27369_ _27369_/A VGND VGND VPWR VPWR _34034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29108_ _34848_/Q _29107_/X _29111_/S VGND VGND VPWR VPWR _29109_/A sky130_fd_sc_hd__mux2_1
X_17122_ _16842_/X _17120_/X _17121_/X _16847_/X VGND VGND VPWR VPWR _17122_/X sky130_fd_sc_hd__a22o_1
X_30380_ _23199_/X _35429_/Q _30392_/S VGND VGND VPWR VPWR _30381_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17053_ _16849_/X _17051_/X _17052_/X _16852_/X VGND VGND VPWR VPWR _17053_/X sky130_fd_sc_hd__a22o_1
X_29039_ _29039_/A VGND VGND VPWR VPWR _34825_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_43_CLK clkbuf_6_6__f_CLK/X VGND VGND VPWR VPWR _36127_/CLK sky130_fd_sc_hd__clkbuf_16
X_16004_ _16057_/A VGND VGND VPWR VPWR _17956_/A sky130_fd_sc_hd__buf_12
XFILLER_109_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32050_ _36019_/CLK _32050_/D VGND VGND VPWR VPWR _32050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31001_ _35724_/Q _29243_/X _31003_/S VGND VGND VPWR VPWR _31002_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17955_ _17700_/X _17953_/X _17954_/X _17703_/X VGND VGND VPWR VPWR _17955_/X sky130_fd_sc_hd__a22o_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16906_ _34533_/Q _32421_/Q _34405_/Q _34341_/Q _16872_/X _16873_/X VGND VGND VPWR
+ VPWR _16906_/X sky130_fd_sc_hd__mux4_1
X_35740_ _35933_/CLK _35740_/D VGND VGND VPWR VPWR _35740_/Q sky130_fd_sc_hd__dfxtp_1
X_32952_ _36089_/CLK _32952_/D VGND VGND VPWR VPWR _32952_/Q sky130_fd_sc_hd__dfxtp_1
X_17886_ _35777_/Q _35137_/Q _34497_/Q _33857_/Q _17846_/X _17847_/X VGND VGND VPWR
+ VPWR _17886_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31903_ _23274_/X _36151_/Q _31919_/S VGND VGND VPWR VPWR _31904_/A sky130_fd_sc_hd__mux2_1
X_19625_ _34545_/Q _32433_/Q _34417_/Q _34353_/Q _19525_/X _19526_/X VGND VGND VPWR
+ VPWR _19625_/X sky130_fd_sc_hd__mux4_1
X_35671_ _35671_/CLK _35671_/D VGND VGND VPWR VPWR _35671_/Q sky130_fd_sc_hd__dfxtp_1
X_16837_ _35043_/Q _34979_/Q _34915_/Q _34851_/Q _16803_/X _16804_/X VGND VGND VPWR
+ VPWR _16837_/X sky130_fd_sc_hd__mux4_1
X_32883_ _35765_/CLK _32883_/D VGND VGND VPWR VPWR _32883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34622_ _36031_/CLK _34622_/D VGND VGND VPWR VPWR _34622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31834_ _31834_/A VGND VGND VPWR VPWR _36118_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19556_ _34799_/Q _34735_/Q _34671_/Q _34607_/Q _19235_/X _19236_/X VGND VGND VPWR
+ VPWR _19556_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_5_22_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_22_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_207_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16768_ _34274_/Q _34210_/Q _34146_/Q _34082_/Q _16736_/X _16737_/X VGND VGND VPWR
+ VPWR _16768_/X sky130_fd_sc_hd__mux4_1
X_18507_ _34258_/Q _34194_/Q _34130_/Q _34066_/Q _18305_/X _18307_/X VGND VGND VPWR
+ VPWR _18507_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34553_ _35771_/CLK _34553_/D VGND VGND VPWR VPWR _34553_/Q sky130_fd_sc_hd__dfxtp_1
X_31765_ _31813_/S VGND VGND VPWR VPWR _31784_/S sky130_fd_sc_hd__buf_4
X_19487_ _35309_/Q _35245_/Q _35181_/Q _32301_/Q _19306_/X _19307_/X VGND VGND VPWR
+ VPWR _19487_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16699_ _34016_/Q _33952_/Q _33888_/Q _32160_/Q _16667_/X _16668_/X VGND VGND VPWR
+ VPWR _16699_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33504_ _34017_/CLK _33504_/D VGND VGND VPWR VPWR _33504_/Q sky130_fd_sc_hd__dfxtp_1
X_30716_ _30716_/A VGND VGND VPWR VPWR _35588_/D sky130_fd_sc_hd__clkbuf_1
X_18438_ _20203_/A VGND VGND VPWR VPWR _18438_/X sky130_fd_sc_hd__buf_6
X_34484_ _35700_/CLK _34484_/D VGND VGND VPWR VPWR _34484_/Q sky130_fd_sc_hd__dfxtp_1
X_31696_ _36053_/Q input62/X _31700_/S VGND VGND VPWR VPWR _31697_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36223_ _36228_/CLK _36223_/D VGND VGND VPWR VPWR _36223_/Q sky130_fd_sc_hd__dfxtp_1
X_33435_ _36194_/CLK _33435_/D VGND VGND VPWR VPWR _33435_/Q sky130_fd_sc_hd__dfxtp_1
X_18369_ _18356_/X _18361_/X _18366_/X _18368_/X VGND VGND VPWR VPWR _18369_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30647_ _30647_/A VGND VGND VPWR VPWR _35555_/D sky130_fd_sc_hd__clkbuf_1
X_20400_ _20208_/X _20398_/X _20399_/X _20211_/X VGND VGND VPWR VPWR _20400_/X sky130_fd_sc_hd__a22o_1
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36154_ _36154_/CLK _36154_/D VGND VGND VPWR VPWR _36154_/Q sky130_fd_sc_hd__dfxtp_1
X_33366_ _36228_/CLK _33366_/D VGND VGND VPWR VPWR _33366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21380_ _32482_/Q _32354_/Q _32034_/Q _36002_/Q _21170_/X _21311_/X VGND VGND VPWR
+ VPWR _21380_/X sky130_fd_sc_hd__mux4_1
X_30578_ _23313_/X _35523_/Q _30590_/S VGND VGND VPWR VPWR _30579_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35105_ _35807_/CLK _35105_/D VGND VGND VPWR VPWR _35105_/Q sky130_fd_sc_hd__dfxtp_1
X_20331_ _20160_/X _20329_/X _20330_/X _20165_/X VGND VGND VPWR VPWR _20331_/X sky130_fd_sc_hd__a22o_1
X_32317_ _35581_/CLK _32317_/D VGND VGND VPWR VPWR _32317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36085_ _36085_/CLK _36085_/D VGND VGND VPWR VPWR _36085_/Q sky130_fd_sc_hd__dfxtp_1
X_33297_ _36232_/CLK _33297_/D VGND VGND VPWR VPWR _33297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_34_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _34017_/CLK sky130_fd_sc_hd__clkbuf_16
X_23050_ input51/X VGND VGND VPWR VPWR _23050_/X sky130_fd_sc_hd__buf_4
XFILLER_179_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35036_ _35036_/CLK _35036_/D VGND VGND VPWR VPWR _35036_/Q sky130_fd_sc_hd__dfxtp_1
X_20262_ _34819_/Q _34755_/Q _34691_/Q _34627_/Q _19941_/X _19942_/X VGND VGND VPWR
+ VPWR _20262_/X sky130_fd_sc_hd__mux4_1
X_32248_ _36152_/CLK _32248_/D VGND VGND VPWR VPWR _32248_/Q sky130_fd_sc_hd__dfxtp_1
X_22001_ _33780_/Q _33716_/Q _33652_/Q _33588_/Q _21796_/X _21797_/X VGND VGND VPWR
+ VPWR _22001_/X sky130_fd_sc_hd__mux4_1
XTAP_6009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20193_ _35329_/Q _35265_/Q _35201_/Q _32321_/Q _20012_/X _20013_/X VGND VGND VPWR
+ VPWR _20193_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32179_ _36063_/CLK _32179_/D VGND VGND VPWR VPWR _32179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23952_ _23047_/X _32516_/Q _23962_/S VGND VGND VPWR VPWR _23953_/A sky130_fd_sc_hd__mux2_1
X_26740_ _33767_/Q _24323_/X _26748_/S VGND VGND VPWR VPWR _26741_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35938_ _35938_/CLK _35938_/D VGND VGND VPWR VPWR _35938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22903_ _22903_/A VGND VGND VPWR VPWR _32021_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26671_ _25168_/X _33735_/Q _26675_/S VGND VGND VPWR VPWR _26672_/A sky130_fd_sc_hd__mux2_1
XTAP_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35869_ _35869_/CLK _35869_/D VGND VGND VPWR VPWR _35869_/Q sky130_fd_sc_hd__dfxtp_1
X_23883_ _22945_/X _32483_/Q _23899_/S VGND VGND VPWR VPWR _23884_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_1014 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_906 _26819_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28410_ _26875_/X _34527_/Q _28414_/S VGND VGND VPWR VPWR _28411_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22834_ _20597_/X _22832_/X _22833_/X _20603_/X VGND VGND VPWR VPWR _22834_/X sky130_fd_sc_hd__a22o_1
X_25622_ _33239_/Q _24273_/X _25622_/S VGND VGND VPWR VPWR _25623_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_917 _26996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29390_ _23093_/X _34960_/Q _29404_/S VGND VGND VPWR VPWR _29391_/A sky130_fd_sc_hd__mux2_1
XANTENNA_928 _28236_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_939 _29092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28341_ _28341_/A VGND VGND VPWR VPWR _34494_/D sky130_fd_sc_hd__clkbuf_1
X_25553_ _25553_/A VGND VGND VPWR VPWR _33207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22765_ _32522_/Q _32394_/Q _32074_/Q _36042_/Q _22582_/X _21607_/A VGND VGND VPWR
+ VPWR _22765_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24504_ _22966_/X _32746_/Q _24506_/S VGND VGND VPWR VPWR _24505_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28272_ _28272_/A VGND VGND VPWR VPWR _34461_/D sky130_fd_sc_hd__clkbuf_1
X_21716_ _21401_/X _21714_/X _21715_/X _21406_/X VGND VGND VPWR VPWR _21716_/X sky130_fd_sc_hd__a22o_1
XFILLER_212_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25484_ _33175_/Q _24273_/X _25484_/S VGND VGND VPWR VPWR _25485_/A sky130_fd_sc_hd__mux2_1
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22696_ _34312_/Q _34248_/Q _34184_/Q _34120_/Q _22395_/X _22396_/X VGND VGND VPWR
+ VPWR _22696_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24435_ _32715_/Q _24434_/X _24441_/S VGND VGND VPWR VPWR _24436_/A sky130_fd_sc_hd__mux2_1
X_27223_ _26919_/X _33965_/Q _27239_/S VGND VGND VPWR VPWR _27224_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21647_ _21647_/A VGND VGND VPWR VPWR _36201_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27154_ _27017_/X _33933_/Q _27154_/S VGND VGND VPWR VPWR _27155_/A sky130_fd_sc_hd__mux2_1
X_24366_ input33/X VGND VGND VPWR VPWR _24366_/X sky130_fd_sc_hd__buf_4
XANTENNA_70 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21578_ _33768_/Q _33704_/Q _33640_/Q _33576_/Q _21443_/X _21444_/X VGND VGND VPWR
+ VPWR _21578_/X sky130_fd_sc_hd__mux4_1
XFILLER_240_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_81 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26105_ _25131_/X _33467_/Q _26113_/S VGND VGND VPWR VPWR _26106_/A sky130_fd_sc_hd__mux2_1
X_23317_ _32223_/Q _23316_/X _23334_/S VGND VGND VPWR VPWR _23318_/A sky130_fd_sc_hd__mux2_1
XANTENNA_92 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20529_ _35852_/Q _32232_/Q _35724_/Q _35660_/Q _18289_/X _18291_/X VGND VGND VPWR
+ VPWR _20529_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27085_ _27154_/S VGND VGND VPWR VPWR _27104_/S sky130_fd_sc_hd__clkbuf_8
X_24297_ _24297_/A VGND VGND VPWR VPWR _32670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_1223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _34142_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_153_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26036_ _25029_/X _33434_/Q _26050_/S VGND VGND VPWR VPWR _26037_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23248_ _32200_/Q _23247_/X _23268_/S VGND VGND VPWR VPWR _23249_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23179_ _23179_/A VGND VGND VPWR VPWR _32172_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1305 _16661_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1316 _32126_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1327 _20295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1338 _19321_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1349 _20660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27987_ _27987_/A VGND VGND VPWR VPWR _34326_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17740_ _17700_/X _17738_/X _17739_/X _17703_/X VGND VGND VPWR VPWR _17740_/X sky130_fd_sc_hd__a22o_1
X_29726_ _29726_/A VGND VGND VPWR VPWR _35119_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26938_ _26937_/X _33843_/Q _26944_/S VGND VGND VPWR VPWR _26939_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_6_12__f_CLK clkbuf_5_6_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_50_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_248_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29657_ _29657_/A VGND VGND VPWR VPWR _35086_/D sky130_fd_sc_hd__clkbuf_1
X_17671_ _35579_/Q _35515_/Q _35451_/Q _35387_/Q _17603_/X _17604_/X VGND VGND VPWR
+ VPWR _17671_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26869_ input7/X VGND VGND VPWR VPWR _26869_/X sky130_fd_sc_hd__buf_4
X_19410_ _19406_/X _19409_/X _19094_/X VGND VGND VPWR VPWR _19418_/C sky130_fd_sc_hd__o21ba_1
XFILLER_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28608_ _26968_/X _34621_/Q _28612_/S VGND VGND VPWR VPWR _28609_/A sky130_fd_sc_hd__mux2_1
X_16622_ _16618_/X _16621_/X _16455_/X VGND VGND VPWR VPWR _16623_/D sky130_fd_sc_hd__o21ba_1
XFILLER_63_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29588_ _35054_/Q _29151_/X _29602_/S VGND VGND VPWR VPWR _29589_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19341_ _19096_/X _19339_/X _19340_/X _19099_/X VGND VGND VPWR VPWR _19341_/X sky130_fd_sc_hd__a22o_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16553_ _34523_/Q _32411_/Q _34395_/Q _34331_/Q _16519_/X _16520_/X VGND VGND VPWR
+ VPWR _16553_/X sky130_fd_sc_hd__mux4_1
X_28539_ _26866_/X _34588_/Q _28549_/S VGND VGND VPWR VPWR _28540_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31550_ _31550_/A VGND VGND VPWR VPWR _35983_/D sky130_fd_sc_hd__clkbuf_1
X_19272_ _34535_/Q _32423_/Q _34407_/Q _34343_/Q _19172_/X _19173_/X VGND VGND VPWR
+ VPWR _19272_/X sky130_fd_sc_hd__mux4_1
X_16484_ _35033_/Q _34969_/Q _34905_/Q _34841_/Q _16450_/X _16451_/X VGND VGND VPWR
+ VPWR _16484_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18223_ _33292_/Q _36172_/Q _33164_/Q _33100_/Q _16028_/X _17157_/A VGND VGND VPWR
+ VPWR _18223_/X sky130_fd_sc_hd__mux4_1
X_30501_ _30501_/A VGND VGND VPWR VPWR _35486_/D sky130_fd_sc_hd__clkbuf_1
X_31481_ _23247_/X _35951_/Q _31493_/S VGND VGND VPWR VPWR _31482_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33220_ _35909_/CLK _33220_/D VGND VGND VPWR VPWR _33220_/Q sky130_fd_sc_hd__dfxtp_1
X_18154_ _18154_/A VGND VGND VPWR VPWR _32009_/D sky130_fd_sc_hd__clkbuf_2
X_30432_ _23297_/X _35454_/Q _30434_/S VGND VGND VPWR VPWR _30433_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17105_ _35755_/Q _35115_/Q _34475_/Q _33835_/Q _16787_/X _16788_/X VGND VGND VPWR
+ VPWR _17105_/X sky130_fd_sc_hd__mux4_1
X_33151_ _36097_/CLK _33151_/D VGND VGND VPWR VPWR _33151_/Q sky130_fd_sc_hd__dfxtp_1
X_18085_ _18081_/X _18084_/X _17853_/X VGND VGND VPWR VPWR _18093_/C sky130_fd_sc_hd__o21ba_1
XFILLER_176_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30363_ _23133_/X _35421_/Q _30371_/S VGND VGND VPWR VPWR _30364_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_16_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _35675_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32102_ _35808_/CLK _32102_/D VGND VGND VPWR VPWR _32102_/Q sky130_fd_sc_hd__dfxtp_1
X_17036_ _33193_/Q _32553_/Q _35945_/Q _35881_/Q _16721_/X _16722_/X VGND VGND VPWR
+ VPWR _17036_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30294_ _35389_/Q _29197_/X _30298_/S VGND VGND VPWR VPWR _30295_/A sky130_fd_sc_hd__mux2_1
X_33082_ _36090_/CLK _33082_/D VGND VGND VPWR VPWR _33082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32033_ _36001_/CLK _32033_/D VGND VGND VPWR VPWR _32033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18987_ _35295_/Q _35231_/Q _35167_/Q _32287_/Q _18953_/X _18954_/X VGND VGND VPWR
+ VPWR _18987_/X sky130_fd_sc_hd__mux4_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _17938_/A VGND VGND VPWR VPWR _32002_/D sky130_fd_sc_hd__clkbuf_2
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33984_ _34305_/CLK _33984_/D VGND VGND VPWR VPWR _33984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35723_ _35787_/CLK _35723_/D VGND VGND VPWR VPWR _35723_/Q sky130_fd_sc_hd__dfxtp_1
X_32935_ _36072_/CLK _32935_/D VGND VGND VPWR VPWR _32935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17869_ _17869_/A _17869_/B _17869_/C _17869_/D VGND VGND VPWR VPWR _17870_/A sky130_fd_sc_hd__or4_4
XFILLER_61_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19608_ _19355_/X _19606_/X _19607_/X _19361_/X VGND VGND VPWR VPWR _19608_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35654_ _35849_/CLK _35654_/D VGND VGND VPWR VPWR _35654_/Q sky130_fd_sc_hd__dfxtp_1
X_20880_ _33236_/Q _36116_/Q _33108_/Q _33044_/Q _20620_/X _20621_/X VGND VGND VPWR
+ VPWR _20880_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32866_ _32994_/CLK _32866_/D VGND VGND VPWR VPWR _32866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34605_ _35304_/CLK _34605_/D VGND VGND VPWR VPWR _34605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31817_ _23077_/X _36110_/Q _31835_/S VGND VGND VPWR VPWR _31818_/A sky130_fd_sc_hd__mux2_1
X_19539_ _19535_/X _19538_/X _19428_/X VGND VGND VPWR VPWR _19563_/A sky130_fd_sc_hd__o21ba_1
X_35585_ _35585_/CLK _35585_/D VGND VGND VPWR VPWR _35585_/Q sky130_fd_sc_hd__dfxtp_1
X_32797_ _34146_/CLK _32797_/D VGND VGND VPWR VPWR _32797_/Q sky130_fd_sc_hd__dfxtp_1
X_22550_ _33027_/Q _32963_/Q _32899_/Q _32835_/Q _22295_/X _22296_/X VGND VGND VPWR
+ VPWR _22550_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34536_ _34922_/CLK _34536_/D VGND VGND VPWR VPWR _34536_/Q sky130_fd_sc_hd__dfxtp_1
X_31748_ _31748_/A VGND VGND VPWR VPWR _36077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21501_ _21246_/X _21499_/X _21500_/X _21249_/X VGND VGND VPWR VPWR _21501_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22481_ _32513_/Q _32385_/Q _32065_/Q _36033_/Q _22229_/X _22370_/X VGND VGND VPWR
+ VPWR _22481_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34467_ _35748_/CLK _34467_/D VGND VGND VPWR VPWR _34467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31679_ _31679_/A VGND VGND VPWR VPWR _36045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36206_ _36211_/CLK _36206_/D VGND VGND VPWR VPWR _36206_/Q sky130_fd_sc_hd__dfxtp_1
X_24220_ _23041_/X _32642_/Q _24234_/S VGND VGND VPWR VPWR _24221_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33418_ _33548_/CLK _33418_/D VGND VGND VPWR VPWR _33418_/Q sky130_fd_sc_hd__dfxtp_1
X_21432_ _21428_/X _21431_/X _21394_/X VGND VGND VPWR VPWR _21440_/C sky130_fd_sc_hd__o21ba_1
X_34398_ _35036_/CLK _34398_/D VGND VGND VPWR VPWR _34398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24151_ _24151_/A VGND VGND VPWR VPWR _32609_/D sky130_fd_sc_hd__clkbuf_1
X_36137_ _36137_/CLK _36137_/D VGND VGND VPWR VPWR _36137_/Q sky130_fd_sc_hd__dfxtp_1
X_33349_ _34050_/CLK _33349_/D VGND VGND VPWR VPWR _33349_/Q sky130_fd_sc_hd__dfxtp_1
X_21363_ _21048_/X _21361_/X _21362_/X _21053_/X VGND VGND VPWR VPWR _21363_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23102_ input56/X VGND VGND VPWR VPWR _23102_/X sky130_fd_sc_hd__buf_6
X_20314_ _20061_/X _20312_/X _20313_/X _20067_/X VGND VGND VPWR VPWR _20314_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24082_ _23038_/X _32577_/Q _24098_/S VGND VGND VPWR VPWR _24083_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36068_ _36069_/CLK _36068_/D VGND VGND VPWR VPWR _36068_/Q sky130_fd_sc_hd__dfxtp_1
X_21294_ _21294_/A VGND VGND VPWR VPWR _36191_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35019_ _35788_/CLK _35019_/D VGND VGND VPWR VPWR _35019_/Q sky130_fd_sc_hd__dfxtp_1
X_23033_ _23033_/A VGND VGND VPWR VPWR _32063_/D sky130_fd_sc_hd__clkbuf_1
X_27910_ _34290_/Q _24357_/X _27916_/S VGND VGND VPWR VPWR _27911_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20245_ _20241_/X _20244_/X _20134_/X VGND VGND VPWR VPWR _20269_/A sky130_fd_sc_hd__o21ba_1
X_28890_ _28890_/A VGND VGND VPWR VPWR _34754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27841_ _34257_/Q _24255_/X _27853_/S VGND VGND VPWR VPWR _27842_/A sky130_fd_sc_hd__mux2_1
XTAP_5105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20176_ _19855_/X _20174_/X _20175_/X _19858_/X VGND VGND VPWR VPWR _20176_/X sky130_fd_sc_hd__a22o_1
XTAP_5116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27772_ _27772_/A VGND VGND VPWR VPWR _34224_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24984_ _24984_/A VGND VGND VPWR VPWR _32971_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29511_ _23336_/X _35018_/Q _29517_/S VGND VGND VPWR VPWR _29512_/A sky130_fd_sc_hd__mux2_1
XTAP_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26723_ _33759_/Q _24298_/X _26727_/S VGND VGND VPWR VPWR _26724_/A sky130_fd_sc_hd__mux2_1
XTAP_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23935_ _23022_/X _32508_/Q _23941_/S VGND VGND VPWR VPWR _23936_/A sky130_fd_sc_hd__mux2_1
XTAP_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29442_ _23228_/X _34985_/Q _29446_/S VGND VGND VPWR VPWR _29443_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26654_ _25143_/X _33727_/Q _26654_/S VGND VGND VPWR VPWR _26655_/A sky130_fd_sc_hd__mux2_1
XANTENNA_703 _22447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23866_ _22920_/X _32475_/Q _23878_/S VGND VGND VPWR VPWR _23867_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_714 _22465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_725 _20703_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_736 _21441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22817_ _20614_/X _22815_/X _22816_/X _20623_/X VGND VGND VPWR VPWR _22817_/X sky130_fd_sc_hd__a22o_1
X_25605_ _25605_/A VGND VGND VPWR VPWR _33230_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29373_ _29373_/A VGND VGND VPWR VPWR _34952_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_747 _22393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_758 _22500_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23797_ _23019_/X _32443_/Q _23805_/S VGND VGND VPWR VPWR _23798_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26585_ _25041_/X _33694_/Q _26591_/S VGND VGND VPWR VPWR _26586_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_769 _22538_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28324_ _34486_/Q _24369_/X _28342_/S VGND VGND VPWR VPWR _28325_/A sky130_fd_sc_hd__mux2_1
X_22748_ _22455_/X _22746_/X _22747_/X _22458_/X VGND VGND VPWR VPWR _22748_/X sky130_fd_sc_hd__a22o_1
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25536_ _25536_/A VGND VGND VPWR VPWR _33199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25467_ _25467_/A VGND VGND VPWR VPWR _33166_/D sky130_fd_sc_hd__clkbuf_1
X_28255_ _28255_/A VGND VGND VPWR VPWR _34453_/D sky130_fd_sc_hd__clkbuf_1
X_22679_ _35847_/Q _32227_/Q _35719_/Q _35655_/Q _20589_/X _20591_/X VGND VGND VPWR
+ VPWR _22679_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24418_ _24418_/A VGND VGND VPWR VPWR _32709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27206_ _26894_/X _33957_/Q _27218_/S VGND VGND VPWR VPWR _27207_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25398_ _25097_/X _33136_/Q _25408_/S VGND VGND VPWR VPWR _25399_/A sky130_fd_sc_hd__mux2_1
X_28186_ _26943_/X _34421_/Q _28186_/S VGND VGND VPWR VPWR _28187_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27137_ _27137_/A VGND VGND VPWR VPWR _33924_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24349_ _32687_/Q _24348_/X _24367_/S VGND VGND VPWR VPWR _24350_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27068_ _27068_/A VGND VGND VPWR VPWR _33891_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26019_ _25004_/X _33426_/Q _26029_/S VGND VGND VPWR VPWR _26020_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18910_ _35741_/Q _35101_/Q _34461_/Q _33821_/Q _18734_/X _18735_/X VGND VGND VPWR
+ VPWR _18910_/X sky130_fd_sc_hd__mux4_1
XTAP_7030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19890_ _34041_/Q _33977_/Q _33913_/Q _32249_/Q _19673_/X _19674_/X VGND VGND VPWR
+ VPWR _19890_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1102 _17368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18841_ _35803_/Q _32178_/Q _35675_/Q _35611_/Q _18554_/X _18555_/X VGND VGND VPWR
+ VPWR _18841_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1113 _28998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1124 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1135 _20155_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1146 _19452_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1157 _22506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18772_ _18768_/X _18771_/X _18730_/X _18731_/X VGND VGND VPWR VPWR _18787_/B sky130_fd_sc_hd__o211a_2
XANTENNA_1168 _22458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15984_ _33742_/Q _33678_/Q _33614_/Q _33550_/Q _15980_/X _15983_/X VGND VGND VPWR
+ VPWR _15984_/X sky130_fd_sc_hd__mux4_1
XTAP_6395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1179 _21125_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17723_ _34301_/Q _34237_/Q _34173_/Q _34109_/Q _17442_/X _17443_/X VGND VGND VPWR
+ VPWR _17723_/X sky130_fd_sc_hd__mux4_1
X_29709_ _29709_/A VGND VGND VPWR VPWR _35111_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30981_ _35714_/Q _29213_/X _30995_/S VGND VGND VPWR VPWR _30982_/A sky130_fd_sc_hd__mux2_1
XTAP_5694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32720_ _36048_/CLK _32720_/D VGND VGND VPWR VPWR _32720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17654_ _17548_/X _17652_/X _17653_/X _17553_/X VGND VGND VPWR VPWR _17654_/X sky130_fd_sc_hd__a22o_1
XTAP_4993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_5_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _34970_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_236_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16605_ _16357_/X _16603_/X _16604_/X _16361_/X VGND VGND VPWR VPWR _16605_/X sky130_fd_sc_hd__a22o_1
XFILLER_223_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32651_ _36171_/CLK _32651_/D VGND VGND VPWR VPWR _32651_/Q sky130_fd_sc_hd__dfxtp_1
X_17585_ _17585_/A VGND VGND VPWR VPWR _31992_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_1_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31602_ _31602_/A VGND VGND VPWR VPWR _36008_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19324_ _19318_/X _19323_/X _19075_/X VGND VGND VPWR VPWR _19346_/A sky130_fd_sc_hd__o21ba_1
X_16536_ _16349_/X _16534_/X _16535_/X _16355_/X VGND VGND VPWR VPWR _16536_/X sky130_fd_sc_hd__a22o_1
X_35370_ _35562_/CLK _35370_/D VGND VGND VPWR VPWR _35370_/Q sky130_fd_sc_hd__dfxtp_1
X_32582_ _35975_/CLK _32582_/D VGND VGND VPWR VPWR _32582_/Q sky130_fd_sc_hd__dfxtp_1
X_34321_ _36204_/CLK _34321_/D VGND VGND VPWR VPWR _34321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31533_ _23330_/X _35976_/Q _31535_/S VGND VGND VPWR VPWR _31534_/A sky130_fd_sc_hd__mux2_1
X_19255_ _19002_/X _19253_/X _19254_/X _19008_/X VGND VGND VPWR VPWR _19255_/X sky130_fd_sc_hd__a22o_1
XFILLER_91_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16467_ _33241_/Q _36121_/Q _33113_/Q _33049_/Q _16352_/X _16353_/X VGND VGND VPWR
+ VPWR _16467_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18206_ _34827_/Q _34763_/Q _34699_/Q _34635_/Q _17994_/X _17995_/X VGND VGND VPWR
+ VPWR _18206_/X sky130_fd_sc_hd__mux4_1
X_34252_ _36048_/CLK _34252_/D VGND VGND VPWR VPWR _34252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31464_ _23220_/X _35943_/Q _31472_/S VGND VGND VPWR VPWR _31465_/A sky130_fd_sc_hd__mux2_1
X_19186_ _19182_/X _19185_/X _19075_/X VGND VGND VPWR VPWR _19210_/A sky130_fd_sc_hd__o21ba_1
XFILLER_145_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16398_ _35799_/Q _32174_/Q _35671_/Q _35607_/Q _16254_/X _16255_/X VGND VGND VPWR
+ VPWR _16398_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33203_ _36141_/CLK _33203_/D VGND VGND VPWR VPWR _33203_/Q sky130_fd_sc_hd__dfxtp_1
X_18137_ _17154_/A _18135_/X _18136_/X _17159_/A VGND VGND VPWR VPWR _18137_/X sky130_fd_sc_hd__a22o_1
X_30415_ _30463_/S VGND VGND VPWR VPWR _30434_/S sky130_fd_sc_hd__buf_6
X_34183_ _34819_/CLK _34183_/D VGND VGND VPWR VPWR _34183_/Q sky130_fd_sc_hd__dfxtp_1
X_31395_ _31395_/A VGND VGND VPWR VPWR _35910_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33134_ _36081_/CLK _33134_/D VGND VGND VPWR VPWR _33134_/Q sky130_fd_sc_hd__dfxtp_1
X_18068_ _33543_/Q _33479_/Q _33415_/Q _33351_/Q _17829_/X _17830_/X VGND VGND VPWR
+ VPWR _18068_/X sky130_fd_sc_hd__mux4_2
XFILLER_176_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30346_ _23108_/X _35413_/Q _30350_/S VGND VGND VPWR VPWR _30347_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1057 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17019_ _33513_/Q _33449_/Q _33385_/Q _33321_/Q _16770_/X _16771_/X VGND VGND VPWR
+ VPWR _17019_/X sky130_fd_sc_hd__mux4_1
X_33065_ _33255_/CLK _33065_/D VGND VGND VPWR VPWR _33065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30277_ _35381_/Q _29172_/X _30277_/S VGND VGND VPWR VPWR _30278_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32016_ _35984_/CLK _32016_/D VGND VGND VPWR VPWR _32016_/Q sky130_fd_sc_hd__dfxtp_1
X_20030_ _20024_/X _20029_/X _19781_/X VGND VGND VPWR VPWR _20052_/A sky130_fd_sc_hd__o21ba_1
XFILLER_217_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_1210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33967_ _36018_/CLK _33967_/D VGND VGND VPWR VPWR _33967_/Q sky130_fd_sc_hd__dfxtp_1
X_21981_ _32499_/Q _32371_/Q _32051_/Q _36019_/Q _21876_/X _21664_/X VGND VGND VPWR
+ VPWR _21981_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23720_ _23720_/A VGND VGND VPWR VPWR _32406_/D sky130_fd_sc_hd__clkbuf_1
X_20932_ _20928_/X _20931_/X _20671_/X VGND VGND VPWR VPWR _20940_/C sky130_fd_sc_hd__o21ba_1
X_32918_ _32983_/CLK _32918_/D VGND VGND VPWR VPWR _32918_/Q sky130_fd_sc_hd__dfxtp_1
X_35706_ _35834_/CLK _35706_/D VGND VGND VPWR VPWR _35706_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33898_ _34282_/CLK _33898_/D VGND VGND VPWR VPWR _33898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23651_ _32375_/Q _23274_/X _23667_/S VGND VGND VPWR VPWR _23652_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32849_ _32978_/CLK _32849_/D VGND VGND VPWR VPWR _32849_/Q sky130_fd_sc_hd__dfxtp_1
X_20863_ _34771_/Q _34707_/Q _34643_/Q _34579_/Q _20829_/X _20830_/X VGND VGND VPWR
+ VPWR _20863_/X sky130_fd_sc_hd__mux4_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35637_ _35828_/CLK _35637_/D VGND VGND VPWR VPWR _35637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22602_ _22598_/X _22601_/X _22467_/X VGND VGND VPWR VPWR _22603_/D sky130_fd_sc_hd__o21ba_1
X_26370_ _26370_/A VGND VGND VPWR VPWR _33592_/D sky130_fd_sc_hd__clkbuf_1
X_23582_ _23582_/A VGND VGND VPWR VPWR _32342_/D sky130_fd_sc_hd__clkbuf_1
X_35568_ _35952_/CLK _35568_/D VGND VGND VPWR VPWR _35568_/Q sky130_fd_sc_hd__dfxtp_1
X_20794_ _33169_/Q _32529_/Q _35921_/Q _35857_/Q _20663_/X _20665_/X VGND VGND VPWR
+ VPWR _20794_/X sky130_fd_sc_hd__mux4_1
X_25321_ _25321_/A VGND VGND VPWR VPWR _33100_/D sky130_fd_sc_hd__clkbuf_1
X_22533_ _34562_/Q _32450_/Q _34434_/Q _34370_/Q _22531_/X _22532_/X VGND VGND VPWR
+ VPWR _22533_/X sky130_fd_sc_hd__mux4_1
X_34519_ _36196_/CLK _34519_/D VGND VGND VPWR VPWR _34519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35499_ _35946_/CLK _35499_/D VGND VGND VPWR VPWR _35499_/Q sky130_fd_sc_hd__dfxtp_1
X_28040_ _28040_/A VGND VGND VPWR VPWR _34351_/D sky130_fd_sc_hd__clkbuf_1
X_25252_ _25252_/A VGND VGND VPWR VPWR _33067_/D sky130_fd_sc_hd__clkbuf_1
X_22464_ _35072_/Q _35008_/Q _34944_/Q _34880_/Q _22462_/X _22463_/X VGND VGND VPWR
+ VPWR _22464_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24203_ _23016_/X _32634_/Q _24213_/S VGND VGND VPWR VPWR _24204_/A sky130_fd_sc_hd__mux2_1
X_21415_ _33507_/Q _33443_/Q _33379_/Q _33315_/Q _21370_/X _21371_/X VGND VGND VPWR
+ VPWR _21415_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25183_ input59/X VGND VGND VPWR VPWR _25183_/X sky130_fd_sc_hd__buf_2
X_22395_ _22395_/A VGND VGND VPWR VPWR _22395_/X sky130_fd_sc_hd__buf_6
XFILLER_120_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24134_ _22914_/X _32601_/Q _24150_/S VGND VGND VPWR VPWR _24135_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21346_ _21302_/X _21344_/X _21345_/X _21308_/X VGND VGND VPWR VPWR _21346_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29991_ _35245_/Q _29148_/X _30007_/S VGND VGND VPWR VPWR _29992_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24065_ _23013_/X _32569_/Q _24077_/S VGND VGND VPWR VPWR _24066_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28942_ _34779_/Q _24286_/X _28954_/S VGND VGND VPWR VPWR _28943_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21277_ _20957_/X _21275_/X _21276_/X _20961_/X VGND VGND VPWR VPWR _21277_/X sky130_fd_sc_hd__a22o_1
XFILLER_46_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23016_ input39/X VGND VGND VPWR VPWR _23016_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_81_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20228_ _34818_/Q _34754_/Q _34690_/Q _34626_/Q _19941_/X _19942_/X VGND VGND VPWR
+ VPWR _20228_/X sky130_fd_sc_hd__mux4_1
X_28873_ _28873_/A VGND VGND VPWR VPWR _34746_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27824_ _27824_/A VGND VGND VPWR VPWR _34249_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20159_ _20155_/X _20156_/X _20157_/X _20158_/X VGND VGND VPWR VPWR _20159_/X sky130_fd_sc_hd__a22o_1
XTAP_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27755_ _27755_/A VGND VGND VPWR VPWR _34216_/D sky130_fd_sc_hd__clkbuf_1
X_24967_ _23044_/X _32963_/Q _24979_/S VGND VGND VPWR VPWR _24968_/A sky130_fd_sc_hd__mux2_1
XTAP_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26706_ _33751_/Q _24273_/X _26706_/S VGND VGND VPWR VPWR _26707_/A sky130_fd_sc_hd__mux2_1
XTAP_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23918_ _22997_/X _32500_/Q _23920_/S VGND VGND VPWR VPWR _23919_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27686_ _34184_/Q _24425_/X _27688_/S VGND VGND VPWR VPWR _27687_/A sky130_fd_sc_hd__mux2_1
XANTENNA_500 _32009_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24898_ _22941_/X _32930_/Q _24916_/S VGND VGND VPWR VPWR _24899_/A sky130_fd_sc_hd__mux2_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_511 _17938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_522 _18004_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29425_ _23145_/X _34977_/Q _29425_/S VGND VGND VPWR VPWR _29426_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26637_ _26637_/A VGND VGND VPWR VPWR _33718_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_533 _20206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23849_ _22895_/X _32467_/Q _23857_/S VGND VGND VPWR VPWR _23850_/A sky130_fd_sc_hd__mux2_1
XTAP_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_544 _20134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_555 _20295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_566 _20147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29356_ _23303_/X _34944_/Q _29374_/S VGND VGND VPWR VPWR _29357_/A sky130_fd_sc_hd__mux2_1
XANTENNA_577 _20153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17370_ _34291_/Q _34227_/Q _34163_/Q _34099_/Q _17089_/X _17090_/X VGND VGND VPWR
+ VPWR _17370_/X sky130_fd_sc_hd__mux4_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26568_ _25016_/X _33686_/Q _26570_/S VGND VGND VPWR VPWR _26569_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_588 _19454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_599 _20167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16321_ _16014_/X _16319_/X _16320_/X _16023_/X VGND VGND VPWR VPWR _16321_/X sky130_fd_sc_hd__a22o_1
X_28307_ _34478_/Q _24345_/X _28321_/S VGND VGND VPWR VPWR _28308_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25519_ _25519_/A VGND VGND VPWR VPWR _33191_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29287_ _29287_/A VGND VGND VPWR VPWR _34911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26499_ _26547_/S VGND VGND VPWR VPWR _26518_/S sky130_fd_sc_hd__buf_4
XFILLER_207_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19040_ _33505_/Q _33441_/Q _33377_/Q _33313_/Q _18717_/X _18718_/X VGND VGND VPWR
+ VPWR _19040_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28238_ _31275_/B _30870_/B VGND VGND VPWR VPWR _28371_/S sky130_fd_sc_hd__nor2_8
XFILLER_186_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16252_ _16026_/X _16250_/X _16251_/X _16037_/X VGND VGND VPWR VPWR _16252_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16183_ _16014_/X _16181_/X _16182_/X _16023_/X VGND VGND VPWR VPWR _16183_/X sky130_fd_sc_hd__a22o_1
X_28169_ _28169_/A VGND VGND VPWR VPWR _34412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30200_ _35344_/Q _29058_/X _30214_/S VGND VGND VPWR VPWR _30201_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput209 _36179_/Q VGND VGND VPWR VPWR D2[5] sky130_fd_sc_hd__buf_2
X_31180_ _31180_/A VGND VGND VPWR VPWR _35808_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19942_ _20295_/A VGND VGND VPWR VPWR _19942_/X sky130_fd_sc_hd__buf_6
X_30131_ _30131_/A VGND VGND VPWR VPWR _35311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30062_ _30062_/A VGND VGND VPWR VPWR _35278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19873_ _19652_/X _19871_/X _19872_/X _19655_/X VGND VGND VPWR VPWR _19873_/X sky130_fd_sc_hd__a22o_1
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_919 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18824_ _18818_/X _18823_/X _18755_/X VGND VGND VPWR VPWR _18825_/D sky130_fd_sc_hd__o21ba_1
XTAP_6170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34870_ _34870_/CLK _34870_/D VGND VGND VPWR VPWR _34870_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33821_ _35933_/CLK _33821_/D VGND VGND VPWR VPWR _33821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18755_ _20167_/A VGND VGND VPWR VPWR _18755_/X sky130_fd_sc_hd__buf_2
XFILLER_209_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17706_ _35580_/Q _35516_/Q _35452_/Q _35388_/Q _17603_/X _17604_/X VGND VGND VPWR
+ VPWR _17706_/X sky130_fd_sc_hd__mux4_1
X_33752_ _35671_/CLK _33752_/D VGND VGND VPWR VPWR _33752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18686_ _18436_/X _18682_/X _18685_/X _18441_/X VGND VGND VPWR VPWR _18686_/X sky130_fd_sc_hd__a22o_1
X_30964_ _35706_/Q _29188_/X _30974_/S VGND VGND VPWR VPWR _30965_/A sky130_fd_sc_hd__mux2_1
XTAP_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32703_ _36097_/CLK _32703_/D VGND VGND VPWR VPWR _32703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17637_ _35578_/Q _35514_/Q _35450_/Q _35386_/Q _17603_/X _17604_/X VGND VGND VPWR
+ VPWR _17637_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33683_ _34259_/CLK _33683_/D VGND VGND VPWR VPWR _33683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30895_ _35673_/Q _29086_/X _30911_/S VGND VGND VPWR VPWR _30896_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35422_ _35808_/CLK _35422_/D VGND VGND VPWR VPWR _35422_/Q sky130_fd_sc_hd__dfxtp_1
X_32634_ _33083_/CLK _32634_/D VGND VGND VPWR VPWR _32634_/Q sky130_fd_sc_hd__dfxtp_1
X_17568_ _35832_/Q _32210_/Q _35704_/Q _35640_/Q _17313_/X _17314_/X VGND VGND VPWR
+ VPWR _17568_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19307_ _19307_/A VGND VGND VPWR VPWR _19307_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_210_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16519_ _17712_/A VGND VGND VPWR VPWR _16519_/X sky130_fd_sc_hd__buf_6
X_35353_ _35801_/CLK _35353_/D VGND VGND VPWR VPWR _35353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32565_ _35958_/CLK _32565_/D VGND VGND VPWR VPWR _32565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17499_ _17352_/X _17497_/X _17498_/X _17355_/X VGND VGND VPWR VPWR _17499_/X sky130_fd_sc_hd__a22o_1
XFILLER_225_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34304_ _34305_/CLK _34304_/D VGND VGND VPWR VPWR _34304_/Q sky130_fd_sc_hd__dfxtp_1
X_31516_ _31543_/S VGND VGND VPWR VPWR _31535_/S sky130_fd_sc_hd__buf_4
X_19238_ _35302_/Q _35238_/Q _35174_/Q _32294_/Q _18953_/X _18954_/X VGND VGND VPWR
+ VPWR _19238_/X sky130_fd_sc_hd__mux4_1
X_35284_ _35284_/CLK _35284_/D VGND VGND VPWR VPWR _35284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32496_ _36078_/CLK _32496_/D VGND VGND VPWR VPWR _32496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34235_ _34298_/CLK _34235_/D VGND VGND VPWR VPWR _34235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31447_ _23139_/X _35935_/Q _31451_/S VGND VGND VPWR VPWR _31448_/A sky130_fd_sc_hd__mux2_1
X_19169_ _34788_/Q _34724_/Q _34660_/Q _34596_/Q _18882_/X _18883_/X VGND VGND VPWR
+ VPWR _19169_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21200_ _32733_/Q _32669_/Q _32605_/Q _36061_/Q _21166_/X _20950_/X VGND VGND VPWR
+ VPWR _21200_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22180_ _34552_/Q _32440_/Q _34424_/Q _34360_/Q _22178_/X _22179_/X VGND VGND VPWR
+ VPWR _22180_/X sky130_fd_sc_hd__mux4_1
X_34166_ _34229_/CLK _34166_/D VGND VGND VPWR VPWR _34166_/Q sky130_fd_sc_hd__dfxtp_1
X_31378_ _31378_/A VGND VGND VPWR VPWR _35902_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21131_ _34011_/Q _33947_/Q _33883_/Q _32155_/Q _20914_/X _20915_/X VGND VGND VPWR
+ VPWR _21131_/X sky130_fd_sc_hd__mux4_1
X_33117_ _33244_/CLK _33117_/D VGND VGND VPWR VPWR _33117_/Q sky130_fd_sc_hd__dfxtp_1
X_30329_ _30329_/A _30329_/B _29049_/B VGND VGND VPWR VPWR _30735_/A sky130_fd_sc_hd__nor3b_4
XFILLER_160_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34097_ _34291_/CLK _34097_/D VGND VGND VPWR VPWR _34097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21062_ _33497_/Q _33433_/Q _33369_/Q _33305_/Q _21017_/X _21018_/X VGND VGND VPWR
+ VPWR _21062_/X sky130_fd_sc_hd__mux4_1
X_33048_ _36123_/CLK _33048_/D VGND VGND VPWR VPWR _33048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20013_ _20013_/A VGND VGND VPWR VPWR _20013_/X sky130_fd_sc_hd__buf_6
XFILLER_119_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25870_ _25183_/X _33356_/Q _25872_/S VGND VGND VPWR VPWR _25871_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24821_ _23028_/X _32894_/Q _24823_/S VGND VGND VPWR VPWR _24822_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34999_ _35257_/CLK _34999_/D VGND VGND VPWR VPWR _34999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27540_ _27540_/A VGND VGND VPWR VPWR _34115_/D sky130_fd_sc_hd__clkbuf_1
X_21964_ _35058_/Q _34994_/Q _34930_/Q _34866_/Q _21756_/X _21757_/X VGND VGND VPWR
+ VPWR _21964_/X sky130_fd_sc_hd__mux4_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24752_ _22926_/X _32861_/Q _24760_/S VGND VGND VPWR VPWR _24753_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23703_ _22875_/X _32398_/Q _23721_/S VGND VGND VPWR VPWR _23704_/A sky130_fd_sc_hd__mux2_1
X_20915_ _22447_/A VGND VGND VPWR VPWR _20915_/X sky130_fd_sc_hd__clkbuf_8
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24683_ _24683_/A VGND VGND VPWR VPWR _32829_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27471_ _27471_/A VGND VGND VPWR VPWR _34082_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21895_ _21754_/X _21893_/X _21894_/X _21759_/X VGND VGND VPWR VPWR _21895_/X sky130_fd_sc_hd__a22o_1
XFILLER_243_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29210_ input47/X VGND VGND VPWR VPWR _29210_/X sky130_fd_sc_hd__buf_4
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26422_ _25001_/X _33617_/Q _26434_/S VGND VGND VPWR VPWR _26423_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23634_ _32367_/Q _23247_/X _23646_/S VGND VGND VPWR VPWR _23635_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20846_ _20842_/X _20845_/X _20611_/X VGND VGND VPWR VPWR _20870_/A sky130_fd_sc_hd__o21ba_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29141_ input22/X VGND VGND VPWR VPWR _29141_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_35_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23565_ _32334_/Q _23077_/X _23583_/S VGND VGND VPWR VPWR _23566_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26353_ _26353_/A VGND VGND VPWR VPWR _33584_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20777_ _33489_/Q _33425_/Q _33361_/Q _33297_/Q _20598_/X _20599_/X VGND VGND VPWR
+ VPWR _20777_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25304_ _25159_/X _33092_/Q _25314_/S VGND VGND VPWR VPWR _25305_/A sky130_fd_sc_hd__mux2_1
X_22516_ _22361_/X _22514_/X _22515_/X _22367_/X VGND VGND VPWR VPWR _22516_/X sky130_fd_sc_hd__a22o_1
X_26284_ _26284_/A VGND VGND VPWR VPWR _33551_/D sky130_fd_sc_hd__clkbuf_1
X_29072_ _29072_/A VGND VGND VPWR VPWR _34836_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23496_ _23496_/A VGND VGND VPWR VPWR _32302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28023_ _28023_/A VGND VGND VPWR VPWR _34343_/D sky130_fd_sc_hd__clkbuf_1
X_22447_ _22447_/A VGND VGND VPWR VPWR _22447_/X sky130_fd_sc_hd__clkbuf_4
X_25235_ _25057_/X _33059_/Q _25251_/S VGND VGND VPWR VPWR _25236_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25166_ _25165_/X _33030_/Q _25175_/S VGND VGND VPWR VPWR _25167_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22378_ _22300_/X _22376_/X _22377_/X _22303_/X VGND VGND VPWR VPWR _22378_/X sky130_fd_sc_hd__a22o_1
XFILLER_159_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24117_ _22889_/X _32593_/Q _24129_/S VGND VGND VPWR VPWR _24118_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21329_ _34528_/Q _32416_/Q _34400_/Q _34336_/Q _21119_/X _21120_/X VGND VGND VPWR
+ VPWR _21329_/X sky130_fd_sc_hd__mux4_1
X_25097_ input28/X VGND VGND VPWR VPWR _25097_/X sky130_fd_sc_hd__buf_2
X_29974_ _35237_/Q _29123_/X _29986_/S VGND VGND VPWR VPWR _29975_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28925_ _34771_/Q _24261_/X _28933_/S VGND VGND VPWR VPWR _28926_/A sky130_fd_sc_hd__mux2_1
X_24048_ _22988_/X _32561_/Q _24056_/S VGND VGND VPWR VPWR _24049_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16870_ _35300_/Q _35236_/Q _35172_/Q _32292_/Q _16653_/X _16654_/X VGND VGND VPWR
+ VPWR _16870_/X sky130_fd_sc_hd__mux4_1
X_28856_ _28856_/A VGND VGND VPWR VPWR _34738_/D sky130_fd_sc_hd__clkbuf_1
X_27807_ _34241_/Q _24404_/X _27823_/S VGND VGND VPWR VPWR _27808_/A sky130_fd_sc_hd__mux2_1
XTAP_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28787_ _28787_/A VGND VGND VPWR VPWR _34705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25999_ _25174_/X _33417_/Q _25999_/S VGND VGND VPWR VPWR _26000_/A sky130_fd_sc_hd__mux2_1
XTAP_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18540_ _33747_/Q _33683_/Q _33619_/Q _33555_/Q _18437_/X _18438_/X VGND VGND VPWR
+ VPWR _18540_/X sky130_fd_sc_hd__mux4_1
XFILLER_218_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27738_ _27738_/A VGND VGND VPWR VPWR _34208_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18471_ _18465_/X _18470_/X _18400_/X VGND VGND VPWR VPWR _18472_/D sky130_fd_sc_hd__o21ba_1
XTAP_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27669_ _27696_/S VGND VGND VPWR VPWR _27688_/S sky130_fd_sc_hd__buf_4
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_330 _32141_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_341 _36205_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_352 _36206_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29408_ _29408_/A VGND VGND VPWR VPWR _34968_/D sky130_fd_sc_hd__clkbuf_1
X_17422_ _17415_/X _17421_/X _17136_/X _17137_/X VGND VGND VPWR VPWR _17439_/B sky130_fd_sc_hd__o211a_1
XANTENNA_363 _36207_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_374 _36208_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30680_ _30680_/A VGND VGND VPWR VPWR _35571_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_385 _36209_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_396 _36210_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29339_ _23277_/X _34936_/Q _29353_/S VGND VGND VPWR VPWR _29340_/A sky130_fd_sc_hd__mux2_1
X_17353_ _35570_/Q _35506_/Q _35442_/Q _35378_/Q _17250_/X _17251_/X VGND VGND VPWR
+ VPWR _17353_/X sky130_fd_sc_hd__mux4_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _34516_/Q _32404_/Q _34388_/Q _34324_/Q _16166_/X _16167_/X VGND VGND VPWR
+ VPWR _16304_/X sky130_fd_sc_hd__mux4_1
X_32350_ _36125_/CLK _32350_/D VGND VGND VPWR VPWR _32350_/Q sky130_fd_sc_hd__dfxtp_1
X_17284_ _35568_/Q _35504_/Q _35440_/Q _35376_/Q _17250_/X _17251_/X VGND VGND VPWR
+ VPWR _17284_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19023_ _33184_/Q _32544_/Q _35936_/Q _35872_/Q _19021_/X _19022_/X VGND VGND VPWR
+ VPWR _19023_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31301_ _31301_/A VGND VGND VPWR VPWR _35865_/D sky130_fd_sc_hd__clkbuf_1
X_16235_ _35026_/Q _34962_/Q _34898_/Q _34834_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _16235_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32281_ _36201_/CLK _32281_/D VGND VGND VPWR VPWR _32281_/Q sky130_fd_sc_hd__dfxtp_1
X_34020_ _34149_/CLK _34020_/D VGND VGND VPWR VPWR _34020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31232_ _35833_/Q input38/X _31244_/S VGND VGND VPWR VPWR _31233_/A sky130_fd_sc_hd__mux2_1
X_16166_ _17712_/A VGND VGND VPWR VPWR _16166_/X sky130_fd_sc_hd__buf_6
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1013 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31163_ _35800_/Q input2/X _31181_/S VGND VGND VPWR VPWR _31164_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16097_ _17159_/A VGND VGND VPWR VPWR _16097_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_142_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30114_ _30114_/A VGND VGND VPWR VPWR _35303_/D sky130_fd_sc_hd__clkbuf_1
X_19925_ _20278_/A VGND VGND VPWR VPWR _19925_/X sky130_fd_sc_hd__buf_6
X_35971_ _35971_/CLK _35971_/D VGND VGND VPWR VPWR _35971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31094_ _31094_/A VGND VGND VPWR VPWR _35767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_296_CLK clkbuf_6_51__f_CLK/X VGND VGND VPWR VPWR _35711_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30045_ _35271_/Q _29228_/X _30049_/S VGND VGND VPWR VPWR _30046_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19856_ _33528_/Q _33464_/Q _33400_/Q _33336_/Q _19776_/X _19777_/X VGND VGND VPWR
+ VPWR _19856_/X sky130_fd_sc_hd__mux4_1
X_34922_ _34922_/CLK _34922_/D VGND VGND VPWR VPWR _34922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18807_ _18657_/X _18805_/X _18806_/X _18661_/X VGND VGND VPWR VPWR _18807_/X sky130_fd_sc_hd__a22o_1
XFILLER_228_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34853_ _35299_/CLK _34853_/D VGND VGND VPWR VPWR _34853_/Q sky130_fd_sc_hd__dfxtp_1
X_19787_ _33014_/Q _32950_/Q _32886_/Q _32822_/Q _19642_/X _19643_/X VGND VGND VPWR
+ VPWR _19787_/X sky130_fd_sc_hd__mux4_1
X_16999_ _17860_/A VGND VGND VPWR VPWR _16999_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_205_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33804_ _36048_/CLK _33804_/D VGND VGND VPWR VPWR _33804_/Q sky130_fd_sc_hd__dfxtp_1
X_18738_ _35544_/Q _35480_/Q _35416_/Q _35352_/Q _18491_/X _18492_/X VGND VGND VPWR
+ VPWR _18738_/X sky130_fd_sc_hd__mux4_1
X_34784_ _35098_/CLK _34784_/D VGND VGND VPWR VPWR _34784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31996_ _34205_/CLK _31996_/D VGND VGND VPWR VPWR _31996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33735_ _34819_/CLK _33735_/D VGND VGND VPWR VPWR _33735_/Q sky130_fd_sc_hd__dfxtp_1
X_18669_ _20232_/A VGND VGND VPWR VPWR _18669_/X sky130_fd_sc_hd__buf_4
X_30947_ _35698_/Q _29163_/X _30953_/S VGND VGND VPWR VPWR _30948_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_1126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20700_ _22467_/A VGND VGND VPWR VPWR _20700_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_240_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33666_ _33795_/CLK _33666_/D VGND VGND VPWR VPWR _33666_/Q sky130_fd_sc_hd__dfxtp_1
X_21680_ _35306_/Q _35242_/Q _35178_/Q _32298_/Q _21606_/X _21607_/X VGND VGND VPWR
+ VPWR _21680_/X sky130_fd_sc_hd__mux4_1
X_30878_ _35665_/Q _29061_/X _30890_/S VGND VGND VPWR VPWR _30879_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35405_ _35792_/CLK _35405_/D VGND VGND VPWR VPWR _35405_/Q sky130_fd_sc_hd__dfxtp_1
X_20631_ _32462_/Q _32334_/Q _32014_/Q _35982_/Q _20628_/X _22463_/A VGND VGND VPWR
+ VPWR _20631_/X sky130_fd_sc_hd__mux4_1
X_32617_ _36137_/CLK _32617_/D VGND VGND VPWR VPWR _32617_/Q sky130_fd_sc_hd__dfxtp_1
X_33597_ _33723_/CLK _33597_/D VGND VGND VPWR VPWR _33597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_220_CLK clkbuf_6_55__f_CLK/X VGND VGND VPWR VPWR _35332_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_225_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35336_ _35337_/CLK _35336_/D VGND VGND VPWR VPWR _35336_/Q sky130_fd_sc_hd__dfxtp_1
X_23350_ _32235_/Q _23234_/X _23350_/S VGND VGND VPWR VPWR _23351_/A sky130_fd_sc_hd__mux2_1
X_20562_ _35597_/Q _35533_/Q _35469_/Q _35405_/Q _18305_/X _18307_/X VGND VGND VPWR
+ VPWR _20562_/X sky130_fd_sc_hd__mux4_1
X_32548_ _35876_/CLK _32548_/D VGND VGND VPWR VPWR _32548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22301_ _35836_/Q _32214_/Q _35708_/Q _35644_/Q _22266_/X _22267_/X VGND VGND VPWR
+ VPWR _22301_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35267_ _35331_/CLK _35267_/D VGND VGND VPWR VPWR _35267_/Q sky130_fd_sc_hd__dfxtp_1
X_23281_ _32211_/Q _23280_/X _23301_/S VGND VGND VPWR VPWR _23282_/A sky130_fd_sc_hd__mux2_1
X_20493_ _33291_/Q _36171_/Q _33163_/Q _33099_/Q _18328_/X _19457_/A VGND VGND VPWR
+ VPWR _20493_/X sky130_fd_sc_hd__mux4_1
X_32479_ _36129_/CLK _32479_/D VGND VGND VPWR VPWR _32479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25020_ _25019_/X _32983_/Q _25020_/S VGND VGND VPWR VPWR _25021_/A sky130_fd_sc_hd__mux2_1
X_22232_ _22016_/X _22230_/X _22231_/X _22020_/X VGND VGND VPWR VPWR _22232_/X sky130_fd_sc_hd__a22o_1
X_34218_ _34281_/CLK _34218_/D VGND VGND VPWR VPWR _34218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35198_ _35583_/CLK _35198_/D VGND VGND VPWR VPWR _35198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22163_ _22008_/X _22161_/X _22162_/X _22014_/X VGND VGND VPWR VPWR _22163_/X sky130_fd_sc_hd__a22o_1
X_34149_ _34149_/CLK _34149_/D VGND VGND VPWR VPWR _34149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21114_ _20893_/X _21112_/X _21113_/X _20896_/X VGND VGND VPWR VPWR _21114_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26971_ input43/X VGND VGND VPWR VPWR _26971_/X sky130_fd_sc_hd__clkbuf_4
X_22094_ _22447_/A VGND VGND VPWR VPWR _22094_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_287_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _36029_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_115_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28710_ _26919_/X _34669_/Q _28726_/S VGND VGND VPWR VPWR _28711_/A sky130_fd_sc_hd__mux2_1
X_25922_ _25060_/X _33380_/Q _25936_/S VGND VGND VPWR VPWR _25923_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21045_ _35288_/Q _35224_/Q _35160_/Q _32280_/Q _20900_/X _20901_/X VGND VGND VPWR
+ VPWR _21045_/X sky130_fd_sc_hd__mux4_1
X_29690_ _29690_/A VGND VGND VPWR VPWR _35102_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28641_ _27017_/X _34637_/Q _28641_/S VGND VGND VPWR VPWR _28642_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25853_ _25853_/A VGND VGND VPWR VPWR _33347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24804_ _24852_/S VGND VGND VPWR VPWR _24823_/S sky130_fd_sc_hd__buf_4
X_28572_ _28641_/S VGND VGND VPWR VPWR _28591_/S sky130_fd_sc_hd__buf_4
X_25784_ _25784_/A VGND VGND VPWR VPWR _33314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22996_ _22996_/A VGND VGND VPWR VPWR _32051_/D sky130_fd_sc_hd__clkbuf_1
X_27523_ _27523_/A VGND VGND VPWR VPWR _34107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24735_ _22901_/X _32853_/Q _24739_/S VGND VGND VPWR VPWR _24736_/A sky130_fd_sc_hd__mux2_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21947_ _22455_/A VGND VGND VPWR VPWR _21947_/X sky130_fd_sc_hd__buf_4
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27454_ _27454_/A VGND VGND VPWR VPWR _34074_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21878_ _33008_/Q _32944_/Q _32880_/Q _32816_/Q _21589_/X _21590_/X VGND VGND VPWR
+ VPWR _21878_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24666_ _24666_/A VGND VGND VPWR VPWR _32821_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26405_ _26405_/A VGND VGND VPWR VPWR _33609_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20829_ _22594_/A VGND VGND VPWR VPWR _20829_/X sky130_fd_sc_hd__buf_6
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23617_ _32359_/Q _23220_/X _23625_/S VGND VGND VPWR VPWR _23618_/A sky130_fd_sc_hd__mux2_1
X_27385_ _34042_/Q _24382_/X _27395_/S VGND VGND VPWR VPWR _27386_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24597_ _24597_/A VGND VGND VPWR VPWR _32788_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_211_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _35784_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_243_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29124_ _34853_/Q _29123_/X _29142_/S VGND VGND VPWR VPWR _29125_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26336_ _26336_/A VGND VGND VPWR VPWR _33576_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23548_ _23548_/A VGND VGND VPWR VPWR _32327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29055_ input12/X VGND VGND VPWR VPWR _29055_/X sky130_fd_sc_hd__buf_2
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26267_ _25171_/X _33544_/Q _26269_/S VGND VGND VPWR VPWR _26268_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23479_ _23479_/A VGND VGND VPWR VPWR _32294_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16020_ _17902_/A VGND VGND VPWR VPWR _16020_/X sky130_fd_sc_hd__buf_4
X_28006_ _28006_/A VGND VGND VPWR VPWR _34335_/D sky130_fd_sc_hd__clkbuf_1
X_25218_ _25032_/X _33051_/Q _25230_/S VGND VGND VPWR VPWR _25219_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26198_ _25069_/X _33511_/Q _26206_/S VGND VGND VPWR VPWR _26199_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25149_ _25149_/A VGND VGND VPWR VPWR _33024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17971_ _33796_/Q _33732_/Q _33668_/Q _33604_/Q _17902_/X _17903_/X VGND VGND VPWR
+ VPWR _17971_/X sky130_fd_sc_hd__mux4_1
X_29957_ _35229_/Q _29098_/X _29965_/S VGND VGND VPWR VPWR _29958_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_278_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _34299_/CLK sky130_fd_sc_hd__clkbuf_16
X_19710_ _32756_/Q _32692_/Q _32628_/Q _36084_/Q _19572_/X _19709_/X VGND VGND VPWR
+ VPWR _19710_/X sky130_fd_sc_hd__mux4_1
X_28908_ _28908_/A VGND VGND VPWR VPWR _34763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16922_ _16702_/X _16920_/X _16921_/X _16708_/X VGND VGND VPWR VPWR _16922_/X sky130_fd_sc_hd__a22o_1
XFILLER_137_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29888_ _29888_/A VGND VGND VPWR VPWR _35196_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19641_ _32498_/Q _32370_/Q _32050_/Q _36018_/Q _19576_/X _19364_/X VGND VGND VPWR
+ VPWR _19641_/X sky130_fd_sc_hd__mux4_1
X_28839_ _28839_/A VGND VGND VPWR VPWR _34730_/D sky130_fd_sc_hd__clkbuf_1
X_16853_ _16849_/X _16850_/X _16851_/X _16852_/X VGND VGND VPWR VPWR _16853_/X sky130_fd_sc_hd__a22o_1
XFILLER_215_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31850_ _23136_/X _36126_/Q _31856_/S VGND VGND VPWR VPWR _31851_/A sky130_fd_sc_hd__mux2_1
X_19572_ _20278_/A VGND VGND VPWR VPWR _19572_/X sky130_fd_sc_hd__buf_6
X_16784_ _17843_/A VGND VGND VPWR VPWR _16784_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_92_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18523_ _35730_/Q _35090_/Q _34450_/Q _33810_/Q _18349_/X _18351_/X VGND VGND VPWR
+ VPWR _18523_/X sky130_fd_sc_hd__mux4_1
X_30801_ _30801_/A VGND VGND VPWR VPWR _35628_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31781_ _31781_/A VGND VGND VPWR VPWR _36093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33520_ _33520_/CLK _33520_/D VGND VGND VPWR VPWR _33520_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_450_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _36004_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30732_ _30732_/A VGND VGND VPWR VPWR _35596_/D sky130_fd_sc_hd__clkbuf_1
X_18454_ _18326_/X _18452_/X _18453_/X _18337_/X VGND VGND VPWR VPWR _18454_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_160 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_171 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _34036_/Q _33972_/Q _33908_/Q _32244_/Q _17373_/X _17374_/X VGND VGND VPWR
+ VPWR _17405_/X sky130_fd_sc_hd__mux4_1
X_33451_ _34870_/CLK _33451_/D VGND VGND VPWR VPWR _33451_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_193 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18385_ _18374_/X _18377_/X _18382_/X _18384_/X VGND VGND VPWR VPWR _18385_/X sky130_fd_sc_hd__a22o_1
X_30663_ _30663_/A VGND VGND VPWR VPWR _35563_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_202_CLK clkbuf_6_54__f_CLK/X VGND VGND VPWR VPWR _35971_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32402_ _35026_/CLK _32402_/D VGND VGND VPWR VPWR _32402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36170_ _36170_/CLK _36170_/D VGND VGND VPWR VPWR _36170_/Q sky130_fd_sc_hd__dfxtp_1
X_17336_ _17202_/X _17334_/X _17335_/X _17205_/X VGND VGND VPWR VPWR _17336_/X sky130_fd_sc_hd__a22o_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33382_ _33702_/CLK _33382_/D VGND VGND VPWR VPWR _33382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30594_ _23339_/X _35531_/Q _30598_/S VGND VGND VPWR VPWR _30595_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35121_ _35953_/CLK _35121_/D VGND VGND VPWR VPWR _35121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32333_ _35277_/CLK _32333_/D VGND VGND VPWR VPWR _32333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17267_ _17195_/X _17265_/X _17266_/X _17200_/X VGND VGND VPWR VPWR _17267_/X sky130_fd_sc_hd__a22o_1
XFILLER_220_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19006_ _20203_/A VGND VGND VPWR VPWR _19006_/X sky130_fd_sc_hd__clkbuf_4
X_16218_ _32466_/Q _32338_/Q _32018_/Q _35986_/Q _16217_/X _17863_/A VGND VGND VPWR
+ VPWR _16218_/X sky130_fd_sc_hd__mux4_1
X_35052_ _35052_/CLK _35052_/D VGND VGND VPWR VPWR _35052_/Q sky130_fd_sc_hd__dfxtp_1
X_32264_ _34816_/CLK _32264_/D VGND VGND VPWR VPWR _32264_/Q sky130_fd_sc_hd__dfxtp_1
X_17198_ _33774_/Q _33710_/Q _33646_/Q _33582_/Q _17196_/X _17197_/X VGND VGND VPWR
+ VPWR _17198_/X sky130_fd_sc_hd__mux4_1
X_34003_ _36232_/CLK _34003_/D VGND VGND VPWR VPWR _34003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31215_ _35825_/Q input29/X _31223_/S VGND VGND VPWR VPWR _31216_/A sky130_fd_sc_hd__mux2_1
X_16149_ _32720_/Q _32656_/Q _32592_/Q _36048_/Q _17862_/A _17713_/A VGND VGND VPWR
+ VPWR _16149_/X sky130_fd_sc_hd__mux4_1
X_32195_ _35818_/CLK _32195_/D VGND VGND VPWR VPWR _32195_/Q sky130_fd_sc_hd__dfxtp_1
X_31146_ _35792_/Q input23/X _31160_/S VGND VGND VPWR VPWR _31147_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_269_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _33729_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19908_ _19902_/X _19907_/X _19800_/X VGND VGND VPWR VPWR _19916_/C sky130_fd_sc_hd__o21ba_1
X_31077_ _31077_/A VGND VGND VPWR VPWR _35759_/D sky130_fd_sc_hd__clkbuf_1
X_35954_ _35954_/CLK _35954_/D VGND VGND VPWR VPWR _35954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30028_ _35263_/Q _29203_/X _30028_/S VGND VGND VPWR VPWR _30029_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_1158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34905_ _35293_/CLK _34905_/D VGND VGND VPWR VPWR _34905_/Q sky130_fd_sc_hd__dfxtp_1
X_19839_ _34807_/Q _34743_/Q _34679_/Q _34615_/Q _19588_/X _19589_/X VGND VGND VPWR
+ VPWR _19839_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35885_ _35885_/CLK _35885_/D VGND VGND VPWR VPWR _35885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22850_ _20626_/X _22848_/X _22849_/X _20637_/X VGND VGND VPWR VPWR _22850_/X sky130_fd_sc_hd__a22o_1
X_34836_ _35031_/CLK _34836_/D VGND VGND VPWR VPWR _34836_/Q sky130_fd_sc_hd__dfxtp_1
X_21801_ _21795_/X _21798_/X _21799_/X _21800_/X VGND VGND VPWR VPWR _21801_/X sky130_fd_sc_hd__a22o_1
X_22781_ _20656_/X _22779_/X _22780_/X _20668_/X VGND VGND VPWR VPWR _22781_/X sky130_fd_sc_hd__a22o_1
X_34767_ _35279_/CLK _34767_/D VGND VGND VPWR VPWR _34767_/Q sky130_fd_sc_hd__dfxtp_1
X_31979_ _35293_/CLK _31979_/D VGND VGND VPWR VPWR _31979_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_441_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _36072_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_225_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24520_ _24520_/A VGND VGND VPWR VPWR _32753_/D sky130_fd_sc_hd__clkbuf_1
X_21732_ _21655_/X _21730_/X _21731_/X _21661_/X VGND VGND VPWR VPWR _21732_/X sky130_fd_sc_hd__a22o_1
X_33718_ _34039_/CLK _33718_/D VGND VGND VPWR VPWR _33718_/Q sky130_fd_sc_hd__dfxtp_1
X_34698_ _35338_/CLK _34698_/D VGND VGND VPWR VPWR _34698_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24451_ _24451_/A VGND VGND VPWR VPWR _32720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21663_ _22508_/A VGND VGND VPWR VPWR _21663_/X sky130_fd_sc_hd__buf_4
XFILLER_178_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33649_ _33779_/CLK _33649_/D VGND VGND VPWR VPWR _33649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23402_ _23402_/A VGND VGND VPWR VPWR _32259_/D sky130_fd_sc_hd__clkbuf_1
X_20614_ _22501_/A VGND VGND VPWR VPWR _20614_/X sky130_fd_sc_hd__buf_2
X_27170_ _26841_/X _33940_/Q _27176_/S VGND VGND VPWR VPWR _27171_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24382_ input39/X VGND VGND VPWR VPWR _24382_/X sky130_fd_sc_hd__clkbuf_4
X_21594_ _22455_/A VGND VGND VPWR VPWR _21594_/X sky130_fd_sc_hd__buf_4
XFILLER_32_1118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26121_ _26121_/A VGND VGND VPWR VPWR _33474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23333_ input55/X VGND VGND VPWR VPWR _23333_/X sky130_fd_sc_hd__buf_4
X_20545_ _33805_/Q _33741_/Q _33677_/Q _33613_/Q _18320_/X _18321_/X VGND VGND VPWR
+ VPWR _20545_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35319_ _35319_/CLK _35319_/D VGND VGND VPWR VPWR _35319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26052_ _26142_/S VGND VGND VPWR VPWR _26071_/S sky130_fd_sc_hd__buf_4
X_23264_ input32/X VGND VGND VPWR VPWR _23264_/X sky130_fd_sc_hd__clkbuf_4
X_20476_ _34826_/Q _34762_/Q _34698_/Q _34634_/Q _20294_/X _20295_/X VGND VGND VPWR
+ VPWR _20476_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25003_ _25003_/A VGND VGND VPWR VPWR _32977_/D sky130_fd_sc_hd__clkbuf_1
X_22215_ _22211_/X _22214_/X _22114_/X VGND VGND VPWR VPWR _22216_/D sky130_fd_sc_hd__o21ba_1
XFILLER_10_1449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23195_ _32180_/Q _23133_/X _23206_/S VGND VGND VPWR VPWR _23196_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29811_ _29922_/S VGND VGND VPWR VPWR _29830_/S sky130_fd_sc_hd__buf_4
XTAP_6703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22146_ _22146_/A _22146_/B _22146_/C _22146_/D VGND VGND VPWR VPWR _22147_/A sky130_fd_sc_hd__or4_4
XFILLER_105_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29742_ _35127_/Q _29179_/X _29758_/S VGND VGND VPWR VPWR _29743_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22077_ _22430_/A VGND VGND VPWR VPWR _22077_/X sky130_fd_sc_hd__clkbuf_4
X_26954_ _26953_/X _33848_/Q _26975_/S VGND VGND VPWR VPWR _26955_/A sky130_fd_sc_hd__mux2_1
XTAP_6769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21028_ _32984_/Q _32920_/Q _32856_/Q _32792_/Q _20883_/X _20884_/X VGND VGND VPWR
+ VPWR _21028_/X sky130_fd_sc_hd__mux4_1
X_25905_ _25035_/X _33372_/Q _25915_/S VGND VGND VPWR VPWR _25906_/A sky130_fd_sc_hd__mux2_1
X_29673_ _29673_/A VGND VGND VPWR VPWR _35094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26885_ _27018_/S VGND VGND VPWR VPWR _26913_/S sky130_fd_sc_hd__buf_4
XFILLER_142_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28624_ _28624_/A VGND VGND VPWR VPWR _34628_/D sky130_fd_sc_hd__clkbuf_1
X_25836_ _25836_/A VGND VGND VPWR VPWR _33339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28555_ _28555_/A VGND VGND VPWR VPWR _34595_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25767_ _25767_/A VGND VGND VPWR VPWR _33306_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22979_ input26/X VGND VGND VPWR VPWR _22979_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_432_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _34154_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27506_ _27506_/A VGND VGND VPWR VPWR _34099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24718_ _31545_/A _27561_/B VGND VGND VPWR VPWR _31410_/B sky130_fd_sc_hd__nor2_8
XFILLER_128_1113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28486_ _26987_/X _34563_/Q _28498_/S VGND VGND VPWR VPWR _28487_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25698_ _33275_/Q _24385_/X _25706_/S VGND VGND VPWR VPWR _25699_/A sky130_fd_sc_hd__mux2_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27437_ _27437_/A VGND VGND VPWR VPWR _34066_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24649_ _22976_/X _32813_/Q _24665_/S VGND VGND VPWR VPWR _24650_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18170_ _35786_/Q _35146_/Q _34506_/Q _33866_/Q _16108_/X _16109_/X VGND VGND VPWR
+ VPWR _18170_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_1351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27368_ _34034_/Q _24357_/X _27374_/S VGND VGND VPWR VPWR _27369_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29107_ input10/X VGND VGND VPWR VPWR _29107_/X sky130_fd_sc_hd__clkbuf_4
X_17121_ _34284_/Q _34220_/Q _34156_/Q _34092_/Q _17089_/X _17090_/X VGND VGND VPWR
+ VPWR _17121_/X sky130_fd_sc_hd__mux4_1
X_26319_ _26319_/A VGND VGND VPWR VPWR _33568_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27299_ _34001_/Q _24255_/X _27311_/S VGND VGND VPWR VPWR _27300_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_35__f_CLK clkbuf_5_17_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_35__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_141_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29038_ _34825_/Q _24428_/X _29038_/S VGND VGND VPWR VPWR _29039_/A sky130_fd_sc_hd__mux2_1
X_17052_ _34026_/Q _33962_/Q _33898_/Q _32234_/Q _17020_/X _17021_/X VGND VGND VPWR
+ VPWR _17052_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16003_ _17911_/A VGND VGND VPWR VPWR _16003_/X sky130_fd_sc_hd__buf_4
XFILLER_174_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31000_ _31000_/A VGND VGND VPWR VPWR _35723_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_946 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17954_ _35779_/Q _35139_/Q _34499_/Q _33859_/Q _17846_/X _17847_/X VGND VGND VPWR
+ VPWR _17954_/X sky130_fd_sc_hd__mux4_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16905_ _16796_/X _16903_/X _16904_/X _16799_/X VGND VGND VPWR VPWR _16905_/X sky130_fd_sc_hd__a22o_1
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32951_ _36024_/CLK _32951_/D VGND VGND VPWR VPWR _32951_/Q sky130_fd_sc_hd__dfxtp_1
X_17885_ _35841_/Q _32220_/Q _35713_/Q _35649_/Q _17666_/X _17667_/X VGND VGND VPWR
+ VPWR _17885_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31902_ _31902_/A VGND VGND VPWR VPWR _36150_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16836_ _34531_/Q _32419_/Q _34403_/Q _34339_/Q _16519_/X _16520_/X VGND VGND VPWR
+ VPWR _16836_/X sky130_fd_sc_hd__mux4_1
X_19624_ _19449_/X _19622_/X _19623_/X _19452_/X VGND VGND VPWR VPWR _19624_/X sky130_fd_sc_hd__a22o_1
X_35670_ _35799_/CLK _35670_/D VGND VGND VPWR VPWR _35670_/Q sky130_fd_sc_hd__dfxtp_1
X_32882_ _35765_/CLK _32882_/D VGND VGND VPWR VPWR _32882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34621_ _36028_/CLK _34621_/D VGND VGND VPWR VPWR _34621_/Q sky130_fd_sc_hd__dfxtp_1
X_31833_ _23111_/X _36118_/Q _31835_/S VGND VGND VPWR VPWR _31834_/A sky130_fd_sc_hd__mux2_1
X_19555_ _19549_/X _19554_/X _19447_/X VGND VGND VPWR VPWR _19563_/C sky130_fd_sc_hd__o21ba_1
XFILLER_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16767_ _33762_/Q _33698_/Q _33634_/Q _33570_/Q _16490_/X _16491_/X VGND VGND VPWR
+ VPWR _16767_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18506_ _33746_/Q _33682_/Q _33618_/Q _33554_/Q _18437_/X _18438_/X VGND VGND VPWR
+ VPWR _18506_/X sky130_fd_sc_hd__mux4_1
XFILLER_206_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_423_CLK clkbuf_6_36__f_CLK/X VGND VGND VPWR VPWR _35187_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_222_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34552_ _35319_/CLK _34552_/D VGND VGND VPWR VPWR _34552_/Q sky130_fd_sc_hd__dfxtp_1
X_19486_ _34797_/Q _34733_/Q _34669_/Q _34605_/Q _19235_/X _19236_/X VGND VGND VPWR
+ VPWR _19486_/X sky130_fd_sc_hd__mux4_1
X_31764_ _31764_/A VGND VGND VPWR VPWR _36085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16698_ _33504_/Q _33440_/Q _33376_/Q _33312_/Q _16417_/X _16418_/X VGND VGND VPWR
+ VPWR _16698_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30715_ _35588_/Q _29219_/X _30725_/S VGND VGND VPWR VPWR _30716_/A sky130_fd_sc_hd__mux2_1
X_18437_ _20202_/A VGND VGND VPWR VPWR _18437_/X sky130_fd_sc_hd__buf_6
XFILLER_146_1246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33503_ _34017_/CLK _33503_/D VGND VGND VPWR VPWR _33503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34483_ _35828_/CLK _34483_/D VGND VGND VPWR VPWR _34483_/Q sky130_fd_sc_hd__dfxtp_1
X_31695_ _31695_/A VGND VGND VPWR VPWR _36052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36222_ _36228_/CLK _36222_/D VGND VGND VPWR VPWR _36222_/Q sky130_fd_sc_hd__dfxtp_1
X_33434_ _33946_/CLK _33434_/D VGND VGND VPWR VPWR _33434_/Q sky130_fd_sc_hd__dfxtp_1
X_18368_ _20165_/A VGND VGND VPWR VPWR _18368_/X sky130_fd_sc_hd__buf_4
X_30646_ _35555_/Q _29117_/X _30662_/S VGND VGND VPWR VPWR _30647_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36153_ _36154_/CLK _36153_/D VGND VGND VPWR VPWR _36153_/Q sky130_fd_sc_hd__dfxtp_1
X_17319_ _33201_/Q _32561_/Q _35953_/Q _35889_/Q _17074_/X _17075_/X VGND VGND VPWR
+ VPWR _17319_/X sky130_fd_sc_hd__mux4_1
X_33365_ _34001_/CLK _33365_/D VGND VGND VPWR VPWR _33365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18299_ _20096_/A VGND VGND VPWR VPWR _18299_/X sky130_fd_sc_hd__clkbuf_4
X_30577_ _30577_/A VGND VGND VPWR VPWR _35522_/D sky130_fd_sc_hd__clkbuf_1
X_20330_ _35077_/Q _35013_/Q _34949_/Q _34885_/Q _20162_/X _20163_/X VGND VGND VPWR
+ VPWR _20330_/X sky130_fd_sc_hd__mux4_1
X_32316_ _35583_/CLK _32316_/D VGND VGND VPWR VPWR _32316_/Q sky130_fd_sc_hd__dfxtp_1
X_35104_ _35745_/CLK _35104_/D VGND VGND VPWR VPWR _35104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36084_ _36149_/CLK _36084_/D VGND VGND VPWR VPWR _36084_/Q sky130_fd_sc_hd__dfxtp_1
X_33296_ _33940_/CLK _33296_/D VGND VGND VPWR VPWR _33296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35035_ _35166_/CLK _35035_/D VGND VGND VPWR VPWR _35035_/Q sky130_fd_sc_hd__dfxtp_1
X_20261_ _20255_/X _20260_/X _20153_/X VGND VGND VPWR VPWR _20269_/C sky130_fd_sc_hd__o21ba_1
X_32247_ _36152_/CLK _32247_/D VGND VGND VPWR VPWR _32247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22000_ _22000_/A VGND VGND VPWR VPWR _36211_/D sky130_fd_sc_hd__buf_6
X_20192_ _34817_/Q _34753_/Q _34689_/Q _34625_/Q _19941_/X _19942_/X VGND VGND VPWR
+ VPWR _20192_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32178_ _35803_/CLK _32178_/D VGND VGND VPWR VPWR _32178_/Q sky130_fd_sc_hd__dfxtp_1
X_31129_ _31129_/A VGND VGND VPWR VPWR _35784_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23951_ _23951_/A VGND VGND VPWR VPWR _32515_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35937_ _35937_/CLK _35937_/D VGND VGND VPWR VPWR _35937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22902_ _22901_/X _32021_/Q _22908_/S VGND VGND VPWR VPWR _22903_/A sky130_fd_sc_hd__mux2_1
X_26670_ _26670_/A VGND VGND VPWR VPWR _33734_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35868_ _35932_/CLK _35868_/D VGND VGND VPWR VPWR _35868_/Q sky130_fd_sc_hd__dfxtp_1
X_23882_ _23882_/A VGND VGND VPWR VPWR _32482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25621_ _25621_/A VGND VGND VPWR VPWR _33238_/D sky130_fd_sc_hd__clkbuf_1
X_34819_ _34819_/CLK _34819_/D VGND VGND VPWR VPWR _34819_/Q sky130_fd_sc_hd__dfxtp_1
X_22833_ _33228_/Q _32588_/Q _35980_/Q _35916_/Q _20675_/X _20676_/X VGND VGND VPWR
+ VPWR _22833_/X sky130_fd_sc_hd__mux4_1
XFILLER_186_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_907 _26769_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_918 _26996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35799_ _35799_/CLK _35799_/D VGND VGND VPWR VPWR _35799_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_929 _28776_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_414_CLK clkbuf_6_33__f_CLK/X VGND VGND VPWR VPWR _35304_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_77_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28340_ _34494_/Q _24394_/X _28342_/S VGND VGND VPWR VPWR _28341_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25552_ _33207_/Q _24373_/X _25568_/S VGND VGND VPWR VPWR _25553_/A sky130_fd_sc_hd__mux2_1
X_22764_ _21749_/A _22762_/X _22763_/X _21752_/A VGND VGND VPWR VPWR _22764_/X sky130_fd_sc_hd__a22o_1
XFILLER_225_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24503_ _24503_/A VGND VGND VPWR VPWR _32745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28271_ _34461_/Q _24292_/X _28279_/S VGND VGND VPWR VPWR _28272_/A sky130_fd_sc_hd__mux2_1
X_21715_ _35051_/Q _34987_/Q _34923_/Q _34859_/Q _21403_/X _21404_/X VGND VGND VPWR
+ VPWR _21715_/X sky130_fd_sc_hd__mux4_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22695_ _33800_/Q _33736_/Q _33672_/Q _33608_/Q _22502_/X _22503_/X VGND VGND VPWR
+ VPWR _22695_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25483_ _25483_/A VGND VGND VPWR VPWR _33174_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27222_ _27222_/A VGND VGND VPWR VPWR _33964_/D sky130_fd_sc_hd__clkbuf_1
X_24434_ input58/X VGND VGND VPWR VPWR _24434_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21646_ _21646_/A _21646_/B _21646_/C _21646_/D VGND VGND VPWR VPWR _21647_/A sky130_fd_sc_hd__or4_4
XFILLER_166_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27153_ _27153_/A VGND VGND VPWR VPWR _33932_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21577_ _21577_/A VGND VGND VPWR VPWR _36199_/D sky130_fd_sc_hd__clkbuf_1
X_24365_ _24365_/A VGND VGND VPWR VPWR _32692_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_60 _32126_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26104_ _26104_/A VGND VGND VPWR VPWR _33466_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_82 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23316_ input50/X VGND VGND VPWR VPWR _23316_/X sky130_fd_sc_hd__buf_4
X_20528_ _20524_/X _20527_/X _20142_/A _20143_/A VGND VGND VPWR VPWR _20543_/B sky130_fd_sc_hd__o211a_1
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_93 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24296_ _32670_/Q _24295_/X _24305_/S VGND VGND VPWR VPWR _24297_/A sky130_fd_sc_hd__mux2_1
X_27084_ _27084_/A VGND VGND VPWR VPWR _33899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26035_ _26035_/A VGND VGND VPWR VPWR _33433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20459_ _34058_/Q _33994_/Q _33930_/Q _32266_/Q _18358_/X _18360_/X VGND VGND VPWR
+ VPWR _20459_/X sky130_fd_sc_hd__mux4_1
X_23247_ input27/X VGND VGND VPWR VPWR _23247_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23178_ _32172_/Q _23108_/X _23182_/S VGND VGND VPWR VPWR _23179_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1306 _16811_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22129_ _33015_/Q _32951_/Q _32887_/Q _32823_/Q _21942_/X _21943_/X VGND VGND VPWR
+ VPWR _22129_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1317 input29/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1328 _20158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1339 _20170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27986_ _26847_/X _34326_/Q _27988_/S VGND VGND VPWR VPWR _27987_/A sky130_fd_sc_hd__mux2_1
XTAP_5821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29725_ _35119_/Q _29154_/X _29737_/S VGND VGND VPWR VPWR _29726_/A sky130_fd_sc_hd__mux2_1
XTAP_6588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26937_ input31/X VGND VGND VPWR VPWR _26937_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29656_ _35086_/Q _29048_/X _29674_/S VGND VGND VPWR VPWR _29657_/A sky130_fd_sc_hd__mux2_1
X_17670_ _17347_/X _17668_/X _17669_/X _17350_/X VGND VGND VPWR VPWR _17670_/X sky130_fd_sc_hd__a22o_1
XFILLER_48_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26868_ _26868_/A VGND VGND VPWR VPWR _33820_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28607_ _28607_/A VGND VGND VPWR VPWR _34620_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16621_ _16448_/X _16619_/X _16620_/X _16453_/X VGND VGND VPWR VPWR _16621_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25819_ _25819_/A VGND VGND VPWR VPWR _33331_/D sky130_fd_sc_hd__clkbuf_1
X_29587_ _29587_/A VGND VGND VPWR VPWR _35053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26799_ _33795_/Q _24410_/X _26811_/S VGND VGND VPWR VPWR _26800_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_405_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _35944_/CLK sky130_fd_sc_hd__clkbuf_16
X_19340_ _35305_/Q _35241_/Q _35177_/Q _32297_/Q _19306_/X _19307_/X VGND VGND VPWR
+ VPWR _19340_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16552_ _16443_/X _16550_/X _16551_/X _16446_/X VGND VGND VPWR VPWR _16552_/X sky130_fd_sc_hd__a22o_1
X_28538_ _28538_/A VGND VGND VPWR VPWR _34587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19271_ _19096_/X _19269_/X _19270_/X _19099_/X VGND VGND VPWR VPWR _19271_/X sky130_fd_sc_hd__a22o_1
X_28469_ _26962_/X _34555_/Q _28477_/S VGND VGND VPWR VPWR _28470_/A sky130_fd_sc_hd__mux2_1
X_16483_ _34521_/Q _32409_/Q _34393_/Q _34329_/Q _16166_/X _16167_/X VGND VGND VPWR
+ VPWR _16483_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18222_ _32780_/Q _32716_/Q _32652_/Q _36108_/Q _17978_/X _16873_/A VGND VGND VPWR
+ VPWR _18222_/X sky130_fd_sc_hd__mux4_1
X_30500_ _23136_/X _35486_/Q _30506_/S VGND VGND VPWR VPWR _30501_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31480_ _31480_/A VGND VGND VPWR VPWR _35950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18153_ _18153_/A _18153_/B _18153_/C _18153_/D VGND VGND VPWR VPWR _18154_/A sky130_fd_sc_hd__or4_4
X_30431_ _30431_/A VGND VGND VPWR VPWR _35453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17104_ _35819_/Q _32196_/Q _35691_/Q _35627_/Q _16960_/X _16961_/X VGND VGND VPWR
+ VPWR _17104_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33150_ _34046_/CLK _33150_/D VGND VGND VPWR VPWR _33150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18084_ _15997_/X _18082_/X _18083_/X _16003_/X VGND VGND VPWR VPWR _18084_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30362_ _30362_/A VGND VGND VPWR VPWR _35420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32101_ _35552_/CLK _32101_/D VGND VGND VPWR VPWR _32101_/Q sky130_fd_sc_hd__dfxtp_1
X_17035_ _35561_/Q _35497_/Q _35433_/Q _35369_/Q _16897_/X _16898_/X VGND VGND VPWR
+ VPWR _17035_/X sky130_fd_sc_hd__mux4_1
XFILLER_171_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33081_ _36090_/CLK _33081_/D VGND VGND VPWR VPWR _33081_/Q sky130_fd_sc_hd__dfxtp_1
X_30293_ _30293_/A VGND VGND VPWR VPWR _35388_/D sky130_fd_sc_hd__clkbuf_1
X_32032_ _36001_/CLK _32032_/D VGND VGND VPWR VPWR _32032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _34783_/Q _34719_/Q _34655_/Q _34591_/Q _18882_/X _18883_/X VGND VGND VPWR
+ VPWR _18986_/X sky130_fd_sc_hd__mux4_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17937_ _17937_/A _17937_/B _17937_/C _17937_/D VGND VGND VPWR VPWR _17938_/A sky130_fd_sc_hd__or4_4
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33983_ _36161_/CLK _33983_/D VGND VGND VPWR VPWR _33983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35722_ _35852_/CLK _35722_/D VGND VGND VPWR VPWR _35722_/Q sky130_fd_sc_hd__dfxtp_1
X_17868_ _17859_/X _17866_/X _17867_/X VGND VGND VPWR VPWR _17869_/D sky130_fd_sc_hd__o21ba_1
XFILLER_22_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32934_ _36007_/CLK _32934_/D VGND VGND VPWR VPWR _32934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19607_ _33265_/Q _36145_/Q _33137_/Q _33073_/Q _19358_/X _19359_/X VGND VGND VPWR
+ VPWR _19607_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_896 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35653_ _35845_/CLK _35653_/D VGND VGND VPWR VPWR _35653_/Q sky130_fd_sc_hd__dfxtp_1
X_16819_ _32739_/Q _32675_/Q _32611_/Q _36067_/Q _16566_/X _16703_/X VGND VGND VPWR
+ VPWR _16819_/X sky130_fd_sc_hd__mux4_1
XFILLER_214_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17799_ _33535_/Q _33471_/Q _33407_/Q _33343_/Q _17476_/X _17477_/X VGND VGND VPWR
+ VPWR _17799_/X sky130_fd_sc_hd__mux4_1
X_32865_ _35481_/CLK _32865_/D VGND VGND VPWR VPWR _32865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34604_ _35242_/CLK _34604_/D VGND VGND VPWR VPWR _34604_/Q sky130_fd_sc_hd__dfxtp_1
X_31816_ _31948_/S VGND VGND VPWR VPWR _31835_/S sky130_fd_sc_hd__buf_4
X_19538_ _19502_/X _19536_/X _19537_/X _19505_/X VGND VGND VPWR VPWR _19538_/X sky130_fd_sc_hd__a22o_1
X_35584_ _35909_/CLK _35584_/D VGND VGND VPWR VPWR _35584_/Q sky130_fd_sc_hd__dfxtp_1
X_32796_ _32860_/CLK _32796_/D VGND VGND VPWR VPWR _32796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31747_ _36077_/Q input25/X _31763_/S VGND VGND VPWR VPWR _31748_/A sky130_fd_sc_hd__mux2_1
X_34535_ _35943_/CLK _34535_/D VGND VGND VPWR VPWR _34535_/Q sky130_fd_sc_hd__dfxtp_1
X_19469_ _34029_/Q _33965_/Q _33901_/Q _32237_/Q _19320_/X _19321_/X VGND VGND VPWR
+ VPWR _19469_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21500_ _33189_/Q _32549_/Q _35941_/Q _35877_/Q _21321_/X _21322_/X VGND VGND VPWR
+ VPWR _21500_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22480_ _22361_/X _22478_/X _22479_/X _22367_/X VGND VGND VPWR VPWR _22480_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31678_ _36045_/Q input60/X _31678_/S VGND VGND VPWR VPWR _31679_/A sky130_fd_sc_hd__mux2_1
X_34466_ _35876_/CLK _34466_/D VGND VGND VPWR VPWR _34466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36205_ _36211_/CLK _36205_/D VGND VGND VPWR VPWR _36205_/Q sky130_fd_sc_hd__dfxtp_1
X_21431_ _21246_/X _21429_/X _21430_/X _21249_/X VGND VGND VPWR VPWR _21431_/X sky130_fd_sc_hd__a22o_1
X_33417_ _33545_/CLK _33417_/D VGND VGND VPWR VPWR _33417_/Q sky130_fd_sc_hd__dfxtp_1
X_30629_ _35547_/Q _29092_/X _30641_/S VGND VGND VPWR VPWR _30630_/A sky130_fd_sc_hd__mux2_1
X_34397_ _35036_/CLK _34397_/D VGND VGND VPWR VPWR _34397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24150_ _22938_/X _32609_/Q _24150_/S VGND VGND VPWR VPWR _24151_/A sky130_fd_sc_hd__mux2_1
X_33348_ _33545_/CLK _33348_/D VGND VGND VPWR VPWR _33348_/Q sky130_fd_sc_hd__dfxtp_1
X_21362_ _35041_/Q _34977_/Q _34913_/Q _34849_/Q _21050_/X _21051_/X VGND VGND VPWR
+ VPWR _21362_/X sky130_fd_sc_hd__mux4_1
X_36136_ _36136_/CLK _36136_/D VGND VGND VPWR VPWR _36136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23101_ _23101_/A VGND VGND VPWR VPWR _32146_/D sky130_fd_sc_hd__clkbuf_1
X_20313_ _33285_/Q _36165_/Q _33157_/Q _33093_/Q _20064_/X _20065_/X VGND VGND VPWR
+ VPWR _20313_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24081_ _24081_/A VGND VGND VPWR VPWR _32576_/D sky130_fd_sc_hd__clkbuf_1
Xinput80 R3[3] VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__clkbuf_4
X_33279_ _36097_/CLK _33279_/D VGND VGND VPWR VPWR _33279_/Q sky130_fd_sc_hd__dfxtp_1
X_36067_ _36067_/CLK _36067_/D VGND VGND VPWR VPWR _36067_/Q sky130_fd_sc_hd__dfxtp_1
X_21293_ _21293_/A _21293_/B _21293_/C _21293_/D VGND VGND VPWR VPWR _21294_/A sky130_fd_sc_hd__or4_2
XFILLER_174_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23032_ _23031_/X _32063_/Q _23032_/S VGND VGND VPWR VPWR _23033_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35018_ _35788_/CLK _35018_/D VGND VGND VPWR VPWR _35018_/Q sky130_fd_sc_hd__dfxtp_1
X_20244_ _20208_/X _20242_/X _20243_/X _20211_/X VGND VGND VPWR VPWR _20244_/X sky130_fd_sc_hd__a22o_1
XFILLER_122_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27840_ _27840_/A VGND VGND VPWR VPWR _34256_/D sky130_fd_sc_hd__clkbuf_1
X_20175_ _34049_/Q _33985_/Q _33921_/Q _32257_/Q _20026_/X _20027_/X VGND VGND VPWR
+ VPWR _20175_/X sky130_fd_sc_hd__mux4_1
XTAP_5106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27771_ _34224_/Q _24351_/X _27781_/S VGND VGND VPWR VPWR _27772_/A sky130_fd_sc_hd__mux2_1
X_24983_ _23068_/X _32971_/Q _24987_/S VGND VGND VPWR VPWR _24984_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29510_ _29510_/A VGND VGND VPWR VPWR _35017_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26722_ _26722_/A VGND VGND VPWR VPWR _33758_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23934_ _23934_/A VGND VGND VPWR VPWR _32507_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29441_ _29441_/A VGND VGND VPWR VPWR _34984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26653_ _26653_/A VGND VGND VPWR VPWR _33726_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23865_ _23865_/A VGND VGND VPWR VPWR _32474_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_704 _22532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_715 _22465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_726 _20804_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25604_ _33230_/Q _24244_/X _25622_/S VGND VGND VPWR VPWR _25605_/A sky130_fd_sc_hd__mux2_1
X_29372_ _23330_/X _34952_/Q _29374_/S VGND VGND VPWR VPWR _29373_/A sky130_fd_sc_hd__mux2_1
X_22816_ _34316_/Q _34252_/Q _34188_/Q _34124_/Q _20645_/X _20646_/X VGND VGND VPWR
+ VPWR _22816_/X sky130_fd_sc_hd__mux4_1
XANTENNA_737 _21479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_748 _22393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26584_ _26584_/A VGND VGND VPWR VPWR _33693_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23796_ _23796_/A VGND VGND VPWR VPWR _32442_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_759 _22500_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28323_ _28371_/S VGND VGND VPWR VPWR _28342_/S sky130_fd_sc_hd__buf_4
XFILLER_41_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25535_ _33199_/Q _24348_/X _25547_/S VGND VGND VPWR VPWR _25536_/A sky130_fd_sc_hd__mux2_1
X_22747_ _35337_/Q _35273_/Q _35209_/Q _32329_/Q _20688_/X _20690_/X VGND VGND VPWR
+ VPWR _22747_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28254_ _34453_/Q _24267_/X _28258_/S VGND VGND VPWR VPWR _28255_/A sky130_fd_sc_hd__mux2_1
X_25466_ _33166_/Q _24244_/X _25484_/S VGND VGND VPWR VPWR _25467_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22678_ _22674_/X _22677_/X _22442_/X _22443_/X VGND VGND VPWR VPWR _22693_/B sky130_fd_sc_hd__o211a_2
XFILLER_186_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27205_ _27205_/A VGND VGND VPWR VPWR _33956_/D sky130_fd_sc_hd__clkbuf_1
X_24417_ _32709_/Q _24416_/X _24429_/S VGND VGND VPWR VPWR _24418_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28185_ _28185_/A VGND VGND VPWR VPWR _34420_/D sky130_fd_sc_hd__clkbuf_1
X_21629_ _33001_/Q _32937_/Q _32873_/Q _32809_/Q _21589_/X _21590_/X VGND VGND VPWR
+ VPWR _21629_/X sky130_fd_sc_hd__mux4_1
X_25397_ _25397_/A VGND VGND VPWR VPWR _33135_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27136_ _26990_/X _33924_/Q _27146_/S VGND VGND VPWR VPWR _27137_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24348_ input27/X VGND VGND VPWR VPWR _24348_/X sky130_fd_sc_hd__buf_6
XFILLER_181_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27067_ _26888_/X _33891_/Q _27083_/S VGND VGND VPWR VPWR _27068_/A sky130_fd_sc_hd__mux2_1
X_24279_ _24279_/A VGND VGND VPWR VPWR _32664_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_21_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_21_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_26018_ _26018_/A VGND VGND VPWR VPWR _33425_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1103 _17400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1114 _24441_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18840_ _18836_/X _18839_/X _18730_/X _18731_/X VGND VGND VPWR VPWR _18857_/B sky130_fd_sc_hd__o211a_2
XTAP_7075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1125 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1136 _20203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1147 _19459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1158 _22506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18771_ _18657_/X _18769_/X _18770_/X _18661_/X VGND VGND VPWR VPWR _18771_/X sky130_fd_sc_hd__a22o_1
XANTENNA_1169 _22458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15983_ _17903_/A VGND VGND VPWR VPWR _15983_/X sky130_fd_sc_hd__buf_6
XTAP_5640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27969_ _28101_/S VGND VGND VPWR VPWR _27988_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17722_ _33789_/Q _33725_/Q _33661_/Q _33597_/Q _17549_/X _17550_/X VGND VGND VPWR
+ VPWR _17722_/X sky130_fd_sc_hd__mux4_1
XTAP_5673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29708_ _35111_/Q _29129_/X _29716_/S VGND VGND VPWR VPWR _29709_/A sky130_fd_sc_hd__mux2_1
XFILLER_209_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30980_ _30980_/A VGND VGND VPWR VPWR _35713_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ _34299_/Q _34235_/Q _34171_/Q _34107_/Q _17442_/X _17443_/X VGND VGND VPWR
+ VPWR _17653_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29639_ _29639_/A VGND VGND VPWR VPWR _35078_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16604_ _32989_/Q _32925_/Q _32861_/Q _32797_/Q _16283_/X _16284_/X VGND VGND VPWR
+ VPWR _16604_/X sky130_fd_sc_hd__mux4_1
X_32650_ _36170_/CLK _32650_/D VGND VGND VPWR VPWR _32650_/Q sky130_fd_sc_hd__dfxtp_1
X_17584_ _17584_/A _17584_/B _17584_/C _17584_/D VGND VGND VPWR VPWR _17585_/A sky130_fd_sc_hd__or4_1
XFILLER_95_1262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31601_ _36008_/Q input19/X _31607_/S VGND VGND VPWR VPWR _31602_/A sky130_fd_sc_hd__mux2_1
X_19323_ _19149_/X _19319_/X _19322_/X _19152_/X VGND VGND VPWR VPWR _19323_/X sky130_fd_sc_hd__a22o_1
X_16535_ _33243_/Q _36123_/Q _33115_/Q _33051_/Q _16352_/X _16353_/X VGND VGND VPWR
+ VPWR _16535_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32581_ _35909_/CLK _32581_/D VGND VGND VPWR VPWR _32581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31532_ _31532_/A VGND VGND VPWR VPWR _35975_/D sky130_fd_sc_hd__clkbuf_1
X_34320_ _35281_/CLK _34320_/D VGND VGND VPWR VPWR _34320_/Q sky130_fd_sc_hd__dfxtp_1
X_19254_ _33255_/Q _36135_/Q _33127_/Q _33063_/Q _19005_/X _19006_/X VGND VGND VPWR
+ VPWR _19254_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16466_ _32729_/Q _32665_/Q _32601_/Q _36057_/Q _16213_/X _16350_/X VGND VGND VPWR
+ VPWR _16466_/X sky130_fd_sc_hd__mux4_1
XFILLER_231_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18205_ _18201_/X _18204_/X _17853_/A VGND VGND VPWR VPWR _18213_/C sky130_fd_sc_hd__o21ba_1
X_34251_ _34251_/CLK _34251_/D VGND VGND VPWR VPWR _34251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31463_ _31463_/A VGND VGND VPWR VPWR _35942_/D sky130_fd_sc_hd__clkbuf_1
X_19185_ _19149_/X _19183_/X _19184_/X _19152_/X VGND VGND VPWR VPWR _19185_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16397_ _16393_/X _16396_/X _16040_/X _16042_/X VGND VGND VPWR VPWR _16412_/B sky130_fd_sc_hd__o211a_1
X_33202_ _36141_/CLK _33202_/D VGND VGND VPWR VPWR _33202_/Q sky130_fd_sc_hd__dfxtp_1
X_18136_ _33033_/Q _32969_/Q _32905_/Q _32841_/Q _15980_/X _15983_/X VGND VGND VPWR
+ VPWR _18136_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30414_ _30414_/A VGND VGND VPWR VPWR _35445_/D sky130_fd_sc_hd__clkbuf_1
X_34182_ _34312_/CLK _34182_/D VGND VGND VPWR VPWR _34182_/Q sky130_fd_sc_hd__dfxtp_1
X_31394_ _35910_/Q input52/X _31400_/S VGND VGND VPWR VPWR _31395_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33133_ _35889_/CLK _33133_/D VGND VGND VPWR VPWR _33133_/Q sky130_fd_sc_hd__dfxtp_1
X_18067_ _17901_/X _18065_/X _18066_/X _17906_/X VGND VGND VPWR VPWR _18067_/X sky130_fd_sc_hd__a22o_1
X_30345_ _30345_/A VGND VGND VPWR VPWR _35412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17018_ _16842_/X _17016_/X _17017_/X _16847_/X VGND VGND VPWR VPWR _17018_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33064_ _34153_/CLK _33064_/D VGND VGND VPWR VPWR _33064_/Q sky130_fd_sc_hd__dfxtp_1
X_30276_ _30276_/A VGND VGND VPWR VPWR _35380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32015_ _36041_/CLK _32015_/D VGND VGND VPWR VPWR _32015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18969_ _34015_/Q _33951_/Q _33887_/Q _32159_/Q _18967_/X _18968_/X VGND VGND VPWR
+ VPWR _18969_/X sky130_fd_sc_hd__mux4_1
XFILLER_230_1222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21980_ _21655_/X _21978_/X _21979_/X _21661_/X VGND VGND VPWR VPWR _21980_/X sky130_fd_sc_hd__a22o_1
X_33966_ _34222_/CLK _33966_/D VGND VGND VPWR VPWR _33966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35705_ _35766_/CLK _35705_/D VGND VGND VPWR VPWR _35705_/Q sky130_fd_sc_hd__dfxtp_1
X_20931_ _20893_/X _20929_/X _20930_/X _20896_/X VGND VGND VPWR VPWR _20931_/X sky130_fd_sc_hd__a22o_1
X_32917_ _32983_/CLK _32917_/D VGND VGND VPWR VPWR _32917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33897_ _36136_/CLK _33897_/D VGND VGND VPWR VPWR _33897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20862_ _20858_/X _20861_/X _20671_/X VGND VGND VPWR VPWR _20870_/C sky130_fd_sc_hd__o21ba_1
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35636_ _35700_/CLK _35636_/D VGND VGND VPWR VPWR _35636_/Q sky130_fd_sc_hd__dfxtp_1
X_23650_ _23650_/A VGND VGND VPWR VPWR _32374_/D sky130_fd_sc_hd__clkbuf_1
X_32848_ _36049_/CLK _32848_/D VGND VGND VPWR VPWR _32848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22601_ _22460_/X _22599_/X _22600_/X _22465_/X VGND VGND VPWR VPWR _22601_/X sky130_fd_sc_hd__a22o_1
XFILLER_165_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_861 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20793_ _35537_/Q _35473_/Q _35409_/Q _35345_/Q _20791_/X _20792_/X VGND VGND VPWR
+ VPWR _20793_/X sky130_fd_sc_hd__mux4_1
X_23581_ _32342_/Q _23111_/X _23583_/S VGND VGND VPWR VPWR _23582_/A sky130_fd_sc_hd__mux2_1
X_35567_ _35951_/CLK _35567_/D VGND VGND VPWR VPWR _35567_/Q sky130_fd_sc_hd__dfxtp_1
X_32779_ _36171_/CLK _32779_/D VGND VGND VPWR VPWR _32779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25320_ _25183_/X _33100_/Q _25322_/S VGND VGND VPWR VPWR _25321_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22532_ _22532_/A VGND VGND VPWR VPWR _22532_/X sky130_fd_sc_hd__buf_4
X_34518_ _34706_/CLK _34518_/D VGND VGND VPWR VPWR _34518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35498_ _35562_/CLK _35498_/D VGND VGND VPWR VPWR _35498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25251_ _25081_/X _33067_/Q _25251_/S VGND VGND VPWR VPWR _25252_/A sky130_fd_sc_hd__mux2_1
X_22463_ _22463_/A VGND VGND VPWR VPWR _22463_/X sky130_fd_sc_hd__buf_4
XFILLER_206_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34449_ _35729_/CLK _34449_/D VGND VGND VPWR VPWR _34449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24202_ _24202_/A VGND VGND VPWR VPWR _32633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21414_ _21089_/X _21412_/X _21413_/X _21094_/X VGND VGND VPWR VPWR _21414_/X sky130_fd_sc_hd__a22o_1
X_25182_ _25182_/A VGND VGND VPWR VPWR _33035_/D sky130_fd_sc_hd__clkbuf_1
X_22394_ _33791_/Q _33727_/Q _33663_/Q _33599_/Q _22149_/X _22150_/X VGND VGND VPWR
+ VPWR _22394_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36119_ _36119_/CLK _36119_/D VGND VGND VPWR VPWR _36119_/Q sky130_fd_sc_hd__dfxtp_1
X_24133_ _24133_/A VGND VGND VPWR VPWR _32600_/D sky130_fd_sc_hd__clkbuf_1
X_21345_ _33249_/Q _36129_/Q _33121_/Q _33057_/Q _21305_/X _21306_/X VGND VGND VPWR
+ VPWR _21345_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29990_ _29990_/A VGND VGND VPWR VPWR _35244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24064_ _24064_/A VGND VGND VPWR VPWR _32568_/D sky130_fd_sc_hd__clkbuf_1
X_28941_ _28941_/A VGND VGND VPWR VPWR _34778_/D sky130_fd_sc_hd__clkbuf_1
X_21276_ _32991_/Q _32927_/Q _32863_/Q _32799_/Q _21236_/X _21237_/X VGND VGND VPWR
+ VPWR _21276_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20227_ _20223_/X _20226_/X _20153_/X VGND VGND VPWR VPWR _20237_/C sky130_fd_sc_hd__o21ba_1
X_23015_ _23015_/A VGND VGND VPWR VPWR _32057_/D sky130_fd_sc_hd__clkbuf_1
X_28872_ _26959_/X _34746_/Q _28882_/S VGND VGND VPWR VPWR _28873_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27823_ _34249_/Q _24428_/X _27823_/S VGND VGND VPWR VPWR _27824_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_1199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20158_ _20158_/A VGND VGND VPWR VPWR _20158_/X sky130_fd_sc_hd__buf_4
XFILLER_172_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27754_ _34216_/Q _24326_/X _27760_/S VGND VGND VPWR VPWR _27755_/A sky130_fd_sc_hd__mux2_1
X_24966_ _24966_/A VGND VGND VPWR VPWR _32962_/D sky130_fd_sc_hd__clkbuf_1
X_20089_ _35070_/Q _35006_/Q _34942_/Q _34878_/Q _19809_/X _19810_/X VGND VGND VPWR
+ VPWR _20089_/X sky130_fd_sc_hd__mux4_1
XTAP_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26705_ _26705_/A VGND VGND VPWR VPWR _33750_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23917_ _23917_/A VGND VGND VPWR VPWR _32499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27685_ _27685_/A VGND VGND VPWR VPWR _34183_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24897_ _24987_/S VGND VGND VPWR VPWR _24916_/S sky130_fd_sc_hd__buf_4
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_501 _32009_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_512 _17938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29424_ _29424_/A VGND VGND VPWR VPWR _34976_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_523 _18004_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26636_ _25115_/X _33718_/Q _26654_/S VGND VGND VPWR VPWR _26637_/A sky130_fd_sc_hd__mux2_1
X_23848_ _23848_/A VGND VGND VPWR VPWR _32466_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_534 _20095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_545 _20134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_556 _20295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_221_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29355_ _29382_/S VGND VGND VPWR VPWR _29374_/S sky130_fd_sc_hd__buf_4
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_567 _20147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26567_ _26567_/A VGND VGND VPWR VPWR _33685_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23779_ _23779_/A VGND VGND VPWR VPWR _32434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_578 _20153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_589 _19457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16320_ _33237_/Q _36117_/Q _33109_/Q _33045_/Q _16020_/X _16021_/X VGND VGND VPWR
+ VPWR _16320_/X sky130_fd_sc_hd__mux4_1
X_28306_ _28306_/A VGND VGND VPWR VPWR _34477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25518_ _33191_/Q _24323_/X _25526_/S VGND VGND VPWR VPWR _25519_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29286_ _23139_/X _34911_/Q _29290_/S VGND VGND VPWR VPWR _29287_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26498_ _26498_/A VGND VGND VPWR VPWR _33653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28237_ _28237_/A VGND VGND VPWR VPWR _34445_/D sky130_fd_sc_hd__clkbuf_1
X_16251_ _32979_/Q _32915_/Q _32851_/Q _32787_/Q _16033_/X _16035_/X VGND VGND VPWR
+ VPWR _16251_/X sky130_fd_sc_hd__mux4_1
X_25449_ _25449_/A VGND VGND VPWR VPWR _33160_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16182_ _33233_/Q _36113_/Q _33105_/Q _33041_/Q _16020_/X _16021_/X VGND VGND VPWR
+ VPWR _16182_/X sky130_fd_sc_hd__mux4_1
X_28168_ _26915_/X _34412_/Q _28186_/S VGND VGND VPWR VPWR _28169_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27119_ _26965_/X _33916_/Q _27125_/S VGND VGND VPWR VPWR _27120_/A sky130_fd_sc_hd__mux2_1
X_28099_ _27014_/X _34380_/Q _28101_/S VGND VGND VPWR VPWR _28100_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30130_ _35311_/Q _29154_/X _30142_/S VGND VGND VPWR VPWR _30131_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19941_ _20294_/A VGND VGND VPWR VPWR _19941_/X sky130_fd_sc_hd__buf_6
XFILLER_153_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30061_ _35278_/Q _29048_/X _30079_/S VGND VGND VPWR VPWR _30062_/A sky130_fd_sc_hd__mux2_1
X_19872_ _33208_/Q _32568_/Q _35960_/Q _35896_/Q _19727_/X _19728_/X VGND VGND VPWR
+ VPWR _19872_/X sky130_fd_sc_hd__mux4_1
XFILLER_229_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18823_ _18748_/X _18821_/X _18822_/X _18753_/X VGND VGND VPWR VPWR _18823_/X sky130_fd_sc_hd__a22o_1
XTAP_6160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33820_ _35933_/CLK _33820_/D VGND VGND VPWR VPWR _33820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18754_ _18748_/X _18749_/X _18752_/X _18753_/X VGND VGND VPWR VPWR _18754_/X sky130_fd_sc_hd__a22o_1
XTAP_5470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17705_ _17860_/A VGND VGND VPWR VPWR _17705_/X sky130_fd_sc_hd__clkbuf_4
X_33751_ _35664_/CLK _33751_/D VGND VGND VPWR VPWR _33751_/Q sky130_fd_sc_hd__dfxtp_1
X_30963_ _30963_/A VGND VGND VPWR VPWR _35705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18685_ _34263_/Q _34199_/Q _34135_/Q _34071_/Q _18683_/X _18684_/X VGND VGND VPWR
+ VPWR _18685_/X sky130_fd_sc_hd__mux4_2
XFILLER_23_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32702_ _36095_/CLK _32702_/D VGND VGND VPWR VPWR _32702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17636_ _17347_/X _17634_/X _17635_/X _17350_/X VGND VGND VPWR VPWR _17636_/X sky130_fd_sc_hd__a22o_1
XFILLER_91_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33682_ _34194_/CLK _33682_/D VGND VGND VPWR VPWR _33682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30894_ _30894_/A VGND VGND VPWR VPWR _35672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35421_ _35935_/CLK _35421_/D VGND VGND VPWR VPWR _35421_/Q sky130_fd_sc_hd__dfxtp_1
X_32633_ _36090_/CLK _32633_/D VGND VGND VPWR VPWR _32633_/Q sky130_fd_sc_hd__dfxtp_1
X_17567_ _17563_/X _17566_/X _17489_/X _17490_/X VGND VGND VPWR VPWR _17584_/B sky130_fd_sc_hd__o211a_1
XFILLER_108_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19306_ _20012_/A VGND VGND VPWR VPWR _19306_/X sky130_fd_sc_hd__buf_4
X_16518_ _16443_/X _16516_/X _16517_/X _16446_/X VGND VGND VPWR VPWR _16518_/X sky130_fd_sc_hd__a22o_1
XFILLER_189_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35352_ _35481_/CLK _35352_/D VGND VGND VPWR VPWR _35352_/Q sky130_fd_sc_hd__dfxtp_1
X_32564_ _35956_/CLK _32564_/D VGND VGND VPWR VPWR _32564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17498_ _33206_/Q _32566_/Q _35958_/Q _35894_/Q _17427_/X _17428_/X VGND VGND VPWR
+ VPWR _17498_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_1038 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34303_ _34303_/CLK _34303_/D VGND VGND VPWR VPWR _34303_/Q sky130_fd_sc_hd__dfxtp_1
X_31515_ _31515_/A VGND VGND VPWR VPWR _35967_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19237_ _34790_/Q _34726_/Q _34662_/Q _34598_/Q _19235_/X _19236_/X VGND VGND VPWR
+ VPWR _19237_/X sky130_fd_sc_hd__mux4_1
X_16449_ _34520_/Q _32408_/Q _34392_/Q _34328_/Q _16166_/X _16167_/X VGND VGND VPWR
+ VPWR _16449_/X sky130_fd_sc_hd__mux4_1
X_35283_ _36211_/CLK _35283_/D VGND VGND VPWR VPWR _35283_/Q sky130_fd_sc_hd__dfxtp_1
X_32495_ _36015_/CLK _32495_/D VGND VGND VPWR VPWR _32495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34234_ _34298_/CLK _34234_/D VGND VGND VPWR VPWR _34234_/Q sky130_fd_sc_hd__dfxtp_1
X_31446_ _31446_/A VGND VGND VPWR VPWR _35934_/D sky130_fd_sc_hd__clkbuf_1
X_19168_ _19164_/X _19167_/X _19094_/X VGND VGND VPWR VPWR _19178_/C sky130_fd_sc_hd__o21ba_1
XFILLER_192_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18119_ _34568_/Q _32456_/Q _34440_/Q _34376_/Q _17931_/X _17932_/X VGND VGND VPWR
+ VPWR _18119_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34165_ _34229_/CLK _34165_/D VGND VGND VPWR VPWR _34165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31377_ _35902_/Q input43/X _31379_/S VGND VGND VPWR VPWR _31378_/A sky130_fd_sc_hd__mux2_1
X_19099_ _19452_/A VGND VGND VPWR VPWR _19099_/X sky130_fd_sc_hd__buf_4
XFILLER_173_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21130_ _33499_/Q _33435_/Q _33371_/Q _33307_/Q _21017_/X _21018_/X VGND VGND VPWR
+ VPWR _21130_/X sky130_fd_sc_hd__mux4_1
X_30328_ _30328_/A VGND VGND VPWR VPWR _35405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33116_ _36124_/CLK _33116_/D VGND VGND VPWR VPWR _33116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34096_ _34286_/CLK _34096_/D VGND VGND VPWR VPWR _34096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33047_ _36117_/CLK _33047_/D VGND VGND VPWR VPWR _33047_/Q sky130_fd_sc_hd__dfxtp_1
X_21061_ _20736_/X _21059_/X _21060_/X _20741_/X VGND VGND VPWR VPWR _21061_/X sky130_fd_sc_hd__a22o_1
X_30259_ _35372_/Q _29144_/X _30277_/S VGND VGND VPWR VPWR _30260_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20012_ _20012_/A VGND VGND VPWR VPWR _20012_/X sky130_fd_sc_hd__buf_6
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24820_ _24820_/A VGND VGND VPWR VPWR _32893_/D sky130_fd_sc_hd__clkbuf_1
X_34998_ _35257_/CLK _34998_/D VGND VGND VPWR VPWR _34998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24751_ _24751_/A VGND VGND VPWR VPWR _32860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21963_ _34546_/Q _32434_/Q _34418_/Q _34354_/Q _21825_/X _21826_/X VGND VGND VPWR
+ VPWR _21963_/X sky130_fd_sc_hd__mux4_1
X_33949_ _34205_/CLK _33949_/D VGND VGND VPWR VPWR _33949_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23702_ _23834_/S VGND VGND VPWR VPWR _23721_/S sky130_fd_sc_hd__clkbuf_8
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20914_ _22446_/A VGND VGND VPWR VPWR _20914_/X sky130_fd_sc_hd__buf_6
X_27470_ _26884_/X _34082_/Q _27488_/S VGND VGND VPWR VPWR _27471_/A sky130_fd_sc_hd__mux2_1
X_24682_ _23025_/X _32829_/Q _24686_/S VGND VGND VPWR VPWR _24683_/A sky130_fd_sc_hd__mux2_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21894_ _35056_/Q _34992_/Q _34928_/Q _34864_/Q _21756_/X _21757_/X VGND VGND VPWR
+ VPWR _21894_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26421_ _26421_/A VGND VGND VPWR VPWR _33616_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23633_ _23633_/A VGND VGND VPWR VPWR _32366_/D sky130_fd_sc_hd__clkbuf_1
X_35619_ _35811_/CLK _35619_/D VGND VGND VPWR VPWR _35619_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20845_ _20743_/X _20843_/X _20844_/X _20746_/X VGND VGND VPWR VPWR _20845_/X sky130_fd_sc_hd__a22o_1
XFILLER_154_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29140_ _29140_/A VGND VGND VPWR VPWR _34858_/D sky130_fd_sc_hd__clkbuf_1
X_26352_ _25097_/X _33584_/Q _26362_/S VGND VGND VPWR VPWR _26353_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23564_ _23696_/S VGND VGND VPWR VPWR _23583_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_39_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20776_ _20736_/X _20774_/X _20775_/X _20741_/X VGND VGND VPWR VPWR _20776_/X sky130_fd_sc_hd__a22o_1
XFILLER_195_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25303_ _25303_/A VGND VGND VPWR VPWR _33091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22515_ _33282_/Q _36162_/Q _33154_/Q _33090_/Q _22364_/X _22365_/X VGND VGND VPWR
+ VPWR _22515_/X sky130_fd_sc_hd__mux4_1
X_29071_ _34836_/Q _29070_/X _29080_/S VGND VGND VPWR VPWR _29072_/A sky130_fd_sc_hd__mux2_1
X_26283_ _24995_/X _33551_/Q _26299_/S VGND VGND VPWR VPWR _26284_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23495_ _22979_/X _32302_/Q _23509_/S VGND VGND VPWR VPWR _23496_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28022_ _26900_/X _34343_/Q _28030_/S VGND VGND VPWR VPWR _28023_/A sky130_fd_sc_hd__mux2_1
X_25234_ _25234_/A VGND VGND VPWR VPWR _33058_/D sky130_fd_sc_hd__clkbuf_1
X_22446_ _22446_/A VGND VGND VPWR VPWR _22446_/X sky130_fd_sc_hd__buf_4
XFILLER_52_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25165_ input52/X VGND VGND VPWR VPWR _25165_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_136_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22377_ _35774_/Q _35134_/Q _34494_/Q _33854_/Q _22093_/X _22094_/X VGND VGND VPWR
+ VPWR _22377_/X sky130_fd_sc_hd__mux4_1
XFILLER_198_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24116_ _24116_/A VGND VGND VPWR VPWR _32592_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21328_ _21043_/X _21326_/X _21327_/X _21046_/X VGND VGND VPWR VPWR _21328_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25096_ _25096_/A VGND VGND VPWR VPWR _33007_/D sky130_fd_sc_hd__clkbuf_1
X_29973_ _29973_/A VGND VGND VPWR VPWR _35236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28924_ _28924_/A VGND VGND VPWR VPWR _34770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21259_ _21048_/X _21257_/X _21258_/X _21053_/X VGND VGND VPWR VPWR _21259_/X sky130_fd_sc_hd__a22o_1
X_24047_ _24047_/A VGND VGND VPWR VPWR _32560_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28855_ _26934_/X _34738_/Q _28861_/S VGND VGND VPWR VPWR _28856_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_1158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27806_ _27806_/A VGND VGND VPWR VPWR _34240_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28786_ _26832_/X _34705_/Q _28798_/S VGND VGND VPWR VPWR _28787_/A sky130_fd_sc_hd__mux2_1
XTAP_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25998_ _25998_/A VGND VGND VPWR VPWR _33416_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27737_ _34208_/Q _24301_/X _27739_/S VGND VGND VPWR VPWR _27738_/A sky130_fd_sc_hd__mux2_1
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24949_ _24949_/A VGND VGND VPWR VPWR _32954_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18470_ _18387_/X _18468_/X _18469_/X _18397_/X VGND VGND VPWR VPWR _18470_/X sky130_fd_sc_hd__a22o_1
XTAP_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27668_ _27668_/A VGND VGND VPWR VPWR _34175_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_320 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_331 _32141_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_342 _36205_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17421_ _17416_/X _17418_/X _17419_/X _17420_/X VGND VGND VPWR VPWR _17421_/X sky130_fd_sc_hd__a22o_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29407_ _23117_/X _34968_/Q _29425_/S VGND VGND VPWR VPWR _29408_/A sky130_fd_sc_hd__mux2_1
X_26619_ _25091_/X _33710_/Q _26633_/S VGND VGND VPWR VPWR _26620_/A sky130_fd_sc_hd__mux2_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_353 _36206_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_364 _36207_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27599_ _27599_/A VGND VGND VPWR VPWR _34142_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_375 _36208_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_386 _36209_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_397 _36210_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17352_ _17860_/A VGND VGND VPWR VPWR _17352_/X sky130_fd_sc_hd__buf_4
XFILLER_207_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29338_ _29338_/A VGND VGND VPWR VPWR _34935_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _16074_/X _16299_/X _16302_/X _16084_/X VGND VGND VPWR VPWR _16303_/X sky130_fd_sc_hd__a22o_1
XFILLER_159_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29269_ _23114_/X _34903_/Q _29269_/S VGND VGND VPWR VPWR _29270_/A sky130_fd_sc_hd__mux2_1
X_17283_ _16994_/X _17281_/X _17282_/X _16997_/X VGND VGND VPWR VPWR _17283_/X sky130_fd_sc_hd__a22o_1
XFILLER_201_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19022_ _20232_/A VGND VGND VPWR VPWR _19022_/X sky130_fd_sc_hd__buf_4
X_31300_ _35865_/Q input3/X _31316_/S VGND VGND VPWR VPWR _31301_/A sky130_fd_sc_hd__mux2_1
X_16234_ _34514_/Q _32402_/Q _34386_/Q _34322_/Q _16166_/X _16167_/X VGND VGND VPWR
+ VPWR _16234_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32280_ _35226_/CLK _32280_/D VGND VGND VPWR VPWR _32280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31231_ _31231_/A VGND VGND VPWR VPWR _35832_/D sky130_fd_sc_hd__clkbuf_1
X_16165_ _16074_/X _16163_/X _16164_/X _16084_/X VGND VGND VPWR VPWR _16165_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_985 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31162_ _31273_/S VGND VGND VPWR VPWR _31181_/S sky130_fd_sc_hd__buf_4
X_16096_ _17773_/A VGND VGND VPWR VPWR _17159_/A sky130_fd_sc_hd__buf_12
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30113_ _35303_/Q _29129_/X _30121_/S VGND VGND VPWR VPWR _30114_/A sky130_fd_sc_hd__mux2_1
X_19924_ _19920_/X _19923_/X _19781_/X VGND VGND VPWR VPWR _19950_/A sky130_fd_sc_hd__o21ba_1
X_35970_ _35970_/CLK _35970_/D VGND VGND VPWR VPWR _35970_/Q sky130_fd_sc_hd__dfxtp_1
X_31093_ _35767_/Q _29179_/X _31109_/S VGND VGND VPWR VPWR _31094_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_1003 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30044_ _30044_/A VGND VGND VPWR VPWR _35270_/D sky130_fd_sc_hd__clkbuf_1
X_34921_ _34987_/CLK _34921_/D VGND VGND VPWR VPWR _34921_/Q sky130_fd_sc_hd__dfxtp_1
X_19855_ _20208_/A VGND VGND VPWR VPWR _19855_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_25_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18806_ _32986_/Q _32922_/Q _32858_/Q _32794_/Q _18583_/X _18584_/X VGND VGND VPWR
+ VPWR _18806_/X sky130_fd_sc_hd__mux4_1
X_34852_ _35300_/CLK _34852_/D VGND VGND VPWR VPWR _34852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19786_ _32502_/Q _32374_/Q _32054_/Q _36022_/Q _19576_/X _19717_/X VGND VGND VPWR
+ VPWR _19786_/X sky130_fd_sc_hd__mux4_1
X_16998_ _16994_/X _16995_/X _16996_/X _16997_/X VGND VGND VPWR VPWR _16998_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33803_ _35464_/CLK _33803_/D VGND VGND VPWR VPWR _33803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18737_ _18588_/X _18733_/X _18736_/X _18591_/X VGND VGND VPWR VPWR _18737_/X sky130_fd_sc_hd__a22o_1
X_34783_ _35743_/CLK _34783_/D VGND VGND VPWR VPWR _34783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31995_ _36185_/CLK _31995_/D VGND VGND VPWR VPWR _31995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33734_ _34308_/CLK _33734_/D VGND VGND VPWR VPWR _33734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18668_ _20231_/A VGND VGND VPWR VPWR _18668_/X sky130_fd_sc_hd__buf_6
X_30946_ _30946_/A VGND VGND VPWR VPWR _35697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17619_ _34298_/Q _34234_/Q _34170_/Q _34106_/Q _17442_/X _17443_/X VGND VGND VPWR
+ VPWR _17619_/X sky130_fd_sc_hd__mux4_1
X_33665_ _33729_/CLK _33665_/D VGND VGND VPWR VPWR _33665_/Q sky130_fd_sc_hd__dfxtp_1
X_30877_ _30877_/A VGND VGND VPWR VPWR _35664_/D sky130_fd_sc_hd__clkbuf_1
X_18599_ _34772_/Q _34708_/Q _34644_/Q _34580_/Q _18529_/X _18530_/X VGND VGND VPWR
+ VPWR _18599_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35404_ _35532_/CLK _35404_/D VGND VGND VPWR VPWR _35404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20630_ _22370_/A VGND VGND VPWR VPWR _22463_/A sky130_fd_sc_hd__buf_4
X_32616_ _36072_/CLK _32616_/D VGND VGND VPWR VPWR _32616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33596_ _34044_/CLK _33596_/D VGND VGND VPWR VPWR _33596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35335_ _35339_/CLK _35335_/D VGND VGND VPWR VPWR _35335_/Q sky130_fd_sc_hd__dfxtp_1
X_20561_ _18277_/X _20559_/X _20560_/X _18287_/X VGND VGND VPWR VPWR _20561_/X sky130_fd_sc_hd__a22o_1
XFILLER_221_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32547_ _35938_/CLK _32547_/D VGND VGND VPWR VPWR _32547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22300_ _22455_/A VGND VGND VPWR VPWR _22300_/X sky130_fd_sc_hd__buf_4
XFILLER_165_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35266_ _35330_/CLK _35266_/D VGND VGND VPWR VPWR _35266_/Q sky130_fd_sc_hd__dfxtp_1
X_20492_ _32779_/Q _32715_/Q _32651_/Q _36107_/Q _20278_/X _19173_/A VGND VGND VPWR
+ VPWR _20492_/X sky130_fd_sc_hd__mux4_1
X_23280_ input38/X VGND VGND VPWR VPWR _23280_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_1002 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32478_ _36065_/CLK _32478_/D VGND VGND VPWR VPWR _32478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22231_ _33018_/Q _32954_/Q _32890_/Q _32826_/Q _21942_/X _21943_/X VGND VGND VPWR
+ VPWR _22231_/X sky130_fd_sc_hd__mux4_1
X_34217_ _34279_/CLK _34217_/D VGND VGND VPWR VPWR _34217_/Q sky130_fd_sc_hd__dfxtp_1
X_31429_ _31429_/A VGND VGND VPWR VPWR _35926_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35197_ _35583_/CLK _35197_/D VGND VGND VPWR VPWR _35197_/Q sky130_fd_sc_hd__dfxtp_1
X_22162_ _33272_/Q _36152_/Q _33144_/Q _33080_/Q _22011_/X _22012_/X VGND VGND VPWR
+ VPWR _22162_/X sky130_fd_sc_hd__mux4_1
XFILLER_161_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34148_ _35992_/CLK _34148_/D VGND VGND VPWR VPWR _34148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21113_ _33178_/Q _32538_/Q _35930_/Q _35866_/Q _20968_/X _20969_/X VGND VGND VPWR
+ VPWR _21113_/X sky130_fd_sc_hd__mux4_1
XTAP_6907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26970_ _26970_/A VGND VGND VPWR VPWR _33853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22093_ _22446_/A VGND VGND VPWR VPWR _22093_/X sky130_fd_sc_hd__buf_4
XTAP_6929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34079_ _34271_/CLK _34079_/D VGND VGND VPWR VPWR _34079_/Q sky130_fd_sc_hd__dfxtp_1
X_25921_ _25921_/A VGND VGND VPWR VPWR _33379_/D sky130_fd_sc_hd__clkbuf_1
X_21044_ _34776_/Q _34712_/Q _34648_/Q _34584_/Q _20829_/X _20830_/X VGND VGND VPWR
+ VPWR _21044_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28640_ _28640_/A VGND VGND VPWR VPWR _34636_/D sky130_fd_sc_hd__clkbuf_1
X_25852_ _25156_/X _33347_/Q _25864_/S VGND VGND VPWR VPWR _25853_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24803_ _24803_/A VGND VGND VPWR VPWR _32885_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_1434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28571_ _28571_/A VGND VGND VPWR VPWR _34603_/D sky130_fd_sc_hd__clkbuf_1
X_25783_ _25053_/X _33314_/Q _25801_/S VGND VGND VPWR VPWR _25784_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22995_ _22994_/X _32051_/Q _23001_/S VGND VGND VPWR VPWR _22996_/A sky130_fd_sc_hd__mux2_1
X_27522_ _26962_/X _34107_/Q _27530_/S VGND VGND VPWR VPWR _27523_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_945 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24734_ _24734_/A VGND VGND VPWR VPWR _32852_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21946_ _21940_/X _21945_/X _21736_/X _21737_/X VGND VGND VPWR VPWR _21967_/B sky130_fd_sc_hd__o211a_1
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27453_ _26860_/X _34074_/Q _27467_/S VGND VGND VPWR VPWR _27454_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24665_ _23000_/X _32821_/Q _24665_/S VGND VGND VPWR VPWR _24666_/A sky130_fd_sc_hd__mux2_1
X_21877_ _32496_/Q _32368_/Q _32048_/Q _36016_/Q _21876_/X _21664_/X VGND VGND VPWR
+ VPWR _21877_/X sky130_fd_sc_hd__mux4_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26404_ _25174_/X _33609_/Q _26404_/S VGND VGND VPWR VPWR _26405_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23616_ _23616_/A VGND VGND VPWR VPWR _32358_/D sky130_fd_sc_hd__clkbuf_1
X_20828_ _20824_/X _20827_/X _20671_/X VGND VGND VPWR VPWR _20838_/C sky130_fd_sc_hd__o21ba_1
X_27384_ _27384_/A VGND VGND VPWR VPWR _34041_/D sky130_fd_sc_hd__clkbuf_1
X_24596_ _22898_/X _32788_/Q _24602_/S VGND VGND VPWR VPWR _24597_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29123_ input16/X VGND VGND VPWR VPWR _29123_/X sky130_fd_sc_hd__buf_2
X_26335_ _25072_/X _33576_/Q _26341_/S VGND VGND VPWR VPWR _26336_/A sky130_fd_sc_hd__mux2_1
X_23547_ _23056_/X _32327_/Q _23551_/S VGND VGND VPWR VPWR _23548_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20759_ _35536_/Q _35472_/Q _35408_/Q _35344_/Q _20658_/X _20660_/X VGND VGND VPWR
+ VPWR _20759_/X sky130_fd_sc_hd__mux4_1
XFILLER_183_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29054_ _29054_/A VGND VGND VPWR VPWR _34830_/D sky130_fd_sc_hd__clkbuf_1
X_26266_ _26266_/A VGND VGND VPWR VPWR _33543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23478_ _22954_/X _32294_/Q _23488_/S VGND VGND VPWR VPWR _23479_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28005_ _26875_/X _34335_/Q _28009_/S VGND VGND VPWR VPWR _28006_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25217_ _25217_/A VGND VGND VPWR VPWR _33050_/D sky130_fd_sc_hd__clkbuf_1
X_22429_ _22429_/A VGND VGND VPWR VPWR _22429_/X sky130_fd_sc_hd__buf_4
X_26197_ _26197_/A VGND VGND VPWR VPWR _33510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25148_ _25146_/X _33024_/Q _25175_/S VGND VGND VPWR VPWR _25149_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17970_ _17970_/A VGND VGND VPWR VPWR _32003_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_123_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29956_ _29956_/A VGND VGND VPWR VPWR _35228_/D sky130_fd_sc_hd__clkbuf_1
X_25079_ _25078_/X _33002_/Q _25082_/S VGND VGND VPWR VPWR _25080_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28907_ _27011_/X _34763_/Q _28911_/S VGND VGND VPWR VPWR _28908_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16921_ _33254_/Q _36134_/Q _33126_/Q _33062_/Q _16705_/X _16706_/X VGND VGND VPWR
+ VPWR _16921_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29887_ _35196_/Q _29194_/X _29893_/S VGND VGND VPWR VPWR _29888_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_1034 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19640_ _19355_/X _19638_/X _19639_/X _19361_/X VGND VGND VPWR VPWR _19640_/X sky130_fd_sc_hd__a22o_1
X_28838_ _26909_/X _34730_/Q _28840_/S VGND VGND VPWR VPWR _28839_/A sky130_fd_sc_hd__mux2_1
X_16852_ _17911_/A VGND VGND VPWR VPWR _16852_/X sky130_fd_sc_hd__buf_4
XFILLER_24_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19571_ _19567_/X _19570_/X _19428_/X VGND VGND VPWR VPWR _19597_/A sky130_fd_sc_hd__o21ba_1
X_16783_ _17842_/A VGND VGND VPWR VPWR _16783_/X sky130_fd_sc_hd__clkbuf_4
X_28769_ _28769_/A VGND VGND VPWR VPWR _34697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_58__f_CLK clkbuf_5_29_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_58__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_248_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18522_ _35794_/Q _32168_/Q _35666_/Q _35602_/Q _18345_/X _18346_/X VGND VGND VPWR
+ VPWR _18522_/X sky130_fd_sc_hd__mux4_1
X_30800_ _23237_/X _35628_/Q _30818_/S VGND VGND VPWR VPWR _30801_/A sky130_fd_sc_hd__mux2_1
X_31780_ _36093_/Q input42/X _31784_/S VGND VGND VPWR VPWR _31781_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30731_ _35596_/Q _29243_/X _30733_/S VGND VGND VPWR VPWR _30732_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18453_ _32976_/Q _32912_/Q _32848_/Q _32784_/Q _18333_/X _18335_/X VGND VGND VPWR
+ VPWR _18453_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_150 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_161 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_172 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _33524_/Q _33460_/Q _33396_/Q _33332_/Q _17123_/X _17124_/X VGND VGND VPWR
+ VPWR _17404_/X sky130_fd_sc_hd__mux4_1
XANTENNA_183 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18384_ _19452_/A VGND VGND VPWR VPWR _18384_/X sky130_fd_sc_hd__buf_4
X_33450_ _33512_/CLK _33450_/D VGND VGND VPWR VPWR _33450_/Q sky130_fd_sc_hd__dfxtp_1
X_30662_ _35563_/Q _29141_/X _30662_/S VGND VGND VPWR VPWR _30663_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_194 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32401_ _36204_/CLK _32401_/D VGND VGND VPWR VPWR _32401_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _34034_/Q _33970_/Q _33906_/Q _32242_/Q _17020_/X _17021_/X VGND VGND VPWR
+ VPWR _17335_/X sky130_fd_sc_hd__mux4_1
XFILLER_186_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30593_ _30593_/A VGND VGND VPWR VPWR _35530_/D sky130_fd_sc_hd__clkbuf_1
X_33381_ _33507_/CLK _33381_/D VGND VGND VPWR VPWR _33381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35120_ _35760_/CLK _35120_/D VGND VGND VPWR VPWR _35120_/Q sky130_fd_sc_hd__dfxtp_1
X_32332_ _35341_/CLK _32332_/D VGND VGND VPWR VPWR _32332_/Q sky130_fd_sc_hd__dfxtp_1
X_17266_ _34288_/Q _34224_/Q _34160_/Q _34096_/Q _17089_/X _17090_/X VGND VGND VPWR
+ VPWR _17266_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16217_ _17982_/A VGND VGND VPWR VPWR _16217_/X sky130_fd_sc_hd__buf_6
X_19005_ _20202_/A VGND VGND VPWR VPWR _19005_/X sky130_fd_sc_hd__buf_4
X_32263_ _34816_/CLK _32263_/D VGND VGND VPWR VPWR _32263_/Q sky130_fd_sc_hd__dfxtp_1
X_35051_ _35944_/CLK _35051_/D VGND VGND VPWR VPWR _35051_/Q sky130_fd_sc_hd__dfxtp_1
X_17197_ _17903_/A VGND VGND VPWR VPWR _17197_/X sky130_fd_sc_hd__clkbuf_4
X_34002_ _34197_/CLK _34002_/D VGND VGND VPWR VPWR _34002_/Q sky130_fd_sc_hd__dfxtp_1
X_31214_ _31214_/A VGND VGND VPWR VPWR _35824_/D sky130_fd_sc_hd__clkbuf_1
X_16148_ _16142_/X _16147_/X _16011_/X VGND VGND VPWR VPWR _16172_/A sky130_fd_sc_hd__o21ba_1
XFILLER_154_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32194_ _35818_/CLK _32194_/D VGND VGND VPWR VPWR _32194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31145_ _31145_/A VGND VGND VPWR VPWR _35791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16079_ _17712_/A VGND VGND VPWR VPWR _16079_/X sky130_fd_sc_hd__buf_6
XFILLER_233_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19907_ _19652_/X _19905_/X _19906_/X _19655_/X VGND VGND VPWR VPWR _19907_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35953_ _35953_/CLK _35953_/D VGND VGND VPWR VPWR _35953_/Q sky130_fd_sc_hd__dfxtp_1
X_31076_ _35759_/Q _29154_/X _31088_/S VGND VGND VPWR VPWR _31077_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30027_ _30027_/A VGND VGND VPWR VPWR _35262_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34904_ _35292_/CLK _34904_/D VGND VGND VPWR VPWR _34904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19838_ _19834_/X _19837_/X _19800_/X VGND VGND VPWR VPWR _19846_/C sky130_fd_sc_hd__o21ba_1
X_35884_ _35885_/CLK _35884_/D VGND VGND VPWR VPWR _35884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34835_ _34967_/CLK _34835_/D VGND VGND VPWR VPWR _34835_/Q sky130_fd_sc_hd__dfxtp_1
Xinput1 DW[0] VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_8
X_19769_ _19454_/X _19767_/X _19768_/X _19459_/X VGND VGND VPWR VPWR _19769_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21800_ _22506_/A VGND VGND VPWR VPWR _21800_/X sky130_fd_sc_hd__buf_2
XFILLER_83_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22780_ _35082_/Q _35018_/Q _34954_/Q _34890_/Q _20679_/X _20681_/X VGND VGND VPWR
+ VPWR _22780_/X sky130_fd_sc_hd__mux4_1
X_34766_ _35215_/CLK _34766_/D VGND VGND VPWR VPWR _34766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31978_ _35293_/CLK _31978_/D VGND VGND VPWR VPWR _31978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21731_ _33260_/Q _36140_/Q _33132_/Q _33068_/Q _21658_/X _21659_/X VGND VGND VPWR
+ VPWR _21731_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33717_ _34292_/CLK _33717_/D VGND VGND VPWR VPWR _33717_/Q sky130_fd_sc_hd__dfxtp_1
X_30929_ _30929_/A VGND VGND VPWR VPWR _35689_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34697_ _35337_/CLK _34697_/D VGND VGND VPWR VPWR _34697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24450_ _22886_/X _32720_/Q _24464_/S VGND VGND VPWR VPWR _24451_/A sky130_fd_sc_hd__mux2_1
X_33648_ _33775_/CLK _33648_/D VGND VGND VPWR VPWR _33648_/Q sky130_fd_sc_hd__dfxtp_1
X_21662_ _21655_/X _21657_/X _21660_/X _21661_/X VGND VGND VPWR VPWR _21662_/X sky130_fd_sc_hd__a22o_1
XFILLER_75_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23401_ _32259_/Q _23313_/X _23413_/S VGND VGND VPWR VPWR _23402_/A sky130_fd_sc_hd__mux2_1
X_20613_ _22361_/A VGND VGND VPWR VPWR _22501_/A sky130_fd_sc_hd__buf_12
X_24381_ _24381_/A VGND VGND VPWR VPWR _32697_/D sky130_fd_sc_hd__clkbuf_1
X_33579_ _35257_/CLK _33579_/D VGND VGND VPWR VPWR _33579_/Q sky130_fd_sc_hd__dfxtp_1
X_21593_ _21587_/X _21592_/X _21383_/X _21384_/X VGND VGND VPWR VPWR _21614_/B sky130_fd_sc_hd__o211a_1
XFILLER_162_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26120_ _25153_/X _33474_/Q _26134_/S VGND VGND VPWR VPWR _26121_/A sky130_fd_sc_hd__mux2_1
X_23332_ _23332_/A VGND VGND VPWR VPWR _32228_/D sky130_fd_sc_hd__clkbuf_1
X_35318_ _35318_/CLK _35318_/D VGND VGND VPWR VPWR _35318_/Q sky130_fd_sc_hd__dfxtp_1
X_20544_ _20544_/A VGND VGND VPWR VPWR _32140_/D sky130_fd_sc_hd__buf_4
XFILLER_137_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26051_ _26051_/A VGND VGND VPWR VPWR _33441_/D sky130_fd_sc_hd__clkbuf_1
X_35249_ _35308_/CLK _35249_/D VGND VGND VPWR VPWR _35249_/Q sky130_fd_sc_hd__dfxtp_1
X_23263_ _23263_/A VGND VGND VPWR VPWR _32205_/D sky130_fd_sc_hd__clkbuf_1
X_20475_ _20471_/X _20474_/X _20153_/A VGND VGND VPWR VPWR _20483_/C sky130_fd_sc_hd__o21ba_1
XFILLER_192_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25002_ _25001_/X _32977_/Q _25020_/S VGND VGND VPWR VPWR _25003_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22214_ _22107_/X _22212_/X _22213_/X _22112_/X VGND VGND VPWR VPWR _22214_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23194_ _23194_/A VGND VGND VPWR VPWR _32179_/D sky130_fd_sc_hd__clkbuf_1
X_29810_ _29810_/A VGND VGND VPWR VPWR _35159_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22145_ _22141_/X _22144_/X _22114_/X VGND VGND VPWR VPWR _22146_/D sky130_fd_sc_hd__o21ba_1
XFILLER_79_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29741_ _29741_/A VGND VGND VPWR VPWR _35126_/D sky130_fd_sc_hd__clkbuf_1
X_22076_ _22429_/A VGND VGND VPWR VPWR _22076_/X sky130_fd_sc_hd__buf_4
X_26953_ input37/X VGND VGND VPWR VPWR _26953_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25904_ _25904_/A VGND VGND VPWR VPWR _33371_/D sky130_fd_sc_hd__clkbuf_1
X_21027_ _32472_/Q _32344_/Q _32024_/Q _35992_/Q _20817_/X _20958_/X VGND VGND VPWR
+ VPWR _21027_/X sky130_fd_sc_hd__mux4_1
X_29672_ _35094_/Q _29076_/X _29674_/S VGND VGND VPWR VPWR _29673_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26884_ input13/X VGND VGND VPWR VPWR _26884_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_248_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28623_ _26990_/X _34628_/Q _28633_/S VGND VGND VPWR VPWR _28624_/A sky130_fd_sc_hd__mux2_1
X_25835_ _25131_/X _33339_/Q _25843_/S VGND VGND VPWR VPWR _25836_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25766_ _25029_/X _33306_/Q _25780_/S VGND VGND VPWR VPWR _25767_/A sky130_fd_sc_hd__mux2_1
X_28554_ _26888_/X _34595_/Q _28570_/S VGND VGND VPWR VPWR _28555_/A sky130_fd_sc_hd__mux2_1
X_22978_ _22978_/A VGND VGND VPWR VPWR _32045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24717_ input83/X input89/X VGND VGND VPWR VPWR _27561_/B sky130_fd_sc_hd__nand2b_4
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27505_ _26937_/X _34099_/Q _27509_/S VGND VGND VPWR VPWR _27506_/A sky130_fd_sc_hd__mux2_1
X_28485_ _28485_/A VGND VGND VPWR VPWR _34562_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21929_ _21929_/A _21929_/B _21929_/C _21929_/D VGND VGND VPWR VPWR _21930_/A sky130_fd_sc_hd__or4_1
X_25697_ _25697_/A VGND VGND VPWR VPWR _33274_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27436_ _26835_/X _34066_/Q _27446_/S VGND VGND VPWR VPWR _27437_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24648_ _24648_/A VGND VGND VPWR VPWR _32812_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27367_ _27367_/A VGND VGND VPWR VPWR _34033_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24579_ _31545_/A _26549_/C VGND VGND VPWR VPWR _27968_/A sky130_fd_sc_hd__nor2_8
XFILLER_180_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_196_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _35970_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17120_ _33772_/Q _33708_/Q _33644_/Q _33580_/Q _16843_/X _16844_/X VGND VGND VPWR
+ VPWR _17120_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29106_ _29106_/A VGND VGND VPWR VPWR _34847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26318_ _25047_/X _33568_/Q _26320_/S VGND VGND VPWR VPWR _26319_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27298_ _27298_/A VGND VGND VPWR VPWR _34000_/D sky130_fd_sc_hd__clkbuf_1
X_29037_ _29037_/A VGND VGND VPWR VPWR _34824_/D sky130_fd_sc_hd__clkbuf_1
X_17051_ _33514_/Q _33450_/Q _33386_/Q _33322_/Q _16770_/X _16771_/X VGND VGND VPWR
+ VPWR _17051_/X sky130_fd_sc_hd__mux4_1
X_26249_ _26249_/A VGND VGND VPWR VPWR _33535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16002_ _17773_/A VGND VGND VPWR VPWR _17911_/A sky130_fd_sc_hd__buf_12
XFILLER_124_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _35843_/Q _32222_/Q _35715_/Q _35651_/Q _17666_/X _17667_/X VGND VGND VPWR
+ VPWR _17953_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29939_ _29939_/A VGND VGND VPWR VPWR _35220_/D sky130_fd_sc_hd__clkbuf_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16904_ _35301_/Q _35237_/Q _35173_/Q _32293_/Q _16653_/X _16654_/X VGND VGND VPWR
+ VPWR _16904_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_120_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _36228_/CLK sky130_fd_sc_hd__clkbuf_16
X_32950_ _36086_/CLK _32950_/D VGND VGND VPWR VPWR _32950_/Q sky130_fd_sc_hd__dfxtp_1
X_17884_ _17880_/X _17883_/X _17842_/X _17843_/X VGND VGND VPWR VPWR _17899_/B sky130_fd_sc_hd__o211a_1
XFILLER_113_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19623_ _35313_/Q _35249_/Q _35185_/Q _32305_/Q _19306_/X _19307_/X VGND VGND VPWR
+ VPWR _19623_/X sky130_fd_sc_hd__mux4_1
X_31901_ _23270_/X _36150_/Q _31919_/S VGND VGND VPWR VPWR _31902_/A sky130_fd_sc_hd__mux2_1
X_16835_ _16796_/X _16833_/X _16834_/X _16799_/X VGND VGND VPWR VPWR _16835_/X sky130_fd_sc_hd__a22o_1
XFILLER_238_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32881_ _33009_/CLK _32881_/D VGND VGND VPWR VPWR _32881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34620_ _34620_/CLK _34620_/D VGND VGND VPWR VPWR _34620_/Q sky130_fd_sc_hd__dfxtp_1
X_31832_ _31832_/A VGND VGND VPWR VPWR _36117_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19554_ _19299_/X _19552_/X _19553_/X _19302_/X VGND VGND VPWR VPWR _19554_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16766_ _16766_/A VGND VGND VPWR VPWR _31969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18505_ _18505_/A VGND VGND VPWR VPWR _32081_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34551_ _35768_/CLK _34551_/D VGND VGND VPWR VPWR _34551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19485_ _19481_/X _19484_/X _19447_/X VGND VGND VPWR VPWR _19493_/C sky130_fd_sc_hd__o21ba_1
XFILLER_80_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16697_ _16489_/X _16695_/X _16696_/X _16494_/X VGND VGND VPWR VPWR _16697_/X sky130_fd_sc_hd__a22o_1
X_31763_ _36085_/Q input33/X _31763_/S VGND VGND VPWR VPWR _31764_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33502_ _34010_/CLK _33502_/D VGND VGND VPWR VPWR _33502_/Q sky130_fd_sc_hd__dfxtp_1
X_30714_ _30714_/A VGND VGND VPWR VPWR _35587_/D sky130_fd_sc_hd__clkbuf_1
X_18436_ _20155_/A VGND VGND VPWR VPWR _18436_/X sky130_fd_sc_hd__buf_4
XFILLER_146_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34482_ _35826_/CLK _34482_/D VGND VGND VPWR VPWR _34482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31694_ _36052_/Q input61/X _31700_/S VGND VGND VPWR VPWR _31695_/A sky130_fd_sc_hd__mux2_1
X_36221_ _36228_/CLK _36221_/D VGND VGND VPWR VPWR _36221_/Q sky130_fd_sc_hd__dfxtp_1
X_33433_ _34267_/CLK _33433_/D VGND VGND VPWR VPWR _33433_/Q sky130_fd_sc_hd__dfxtp_1
X_18367_ _20073_/A VGND VGND VPWR VPWR _20165_/A sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_187_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _35515_/CLK sky130_fd_sc_hd__clkbuf_16
X_30645_ _30645_/A VGND VGND VPWR VPWR _35554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36152_ _36152_/CLK _36152_/D VGND VGND VPWR VPWR _36152_/Q sky130_fd_sc_hd__dfxtp_1
X_17318_ _35569_/Q _35505_/Q _35441_/Q _35377_/Q _17250_/X _17251_/X VGND VGND VPWR
+ VPWR _17318_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33364_ _36237_/CLK _33364_/D VGND VGND VPWR VPWR _33364_/Q sky130_fd_sc_hd__dfxtp_1
X_30576_ _23310_/X _35522_/Q _30590_/S VGND VGND VPWR VPWR _30577_/A sky130_fd_sc_hd__mux2_1
X_18298_ _20095_/A VGND VGND VPWR VPWR _18298_/X sky130_fd_sc_hd__buf_4
XFILLER_200_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35103_ _35296_/CLK _35103_/D VGND VGND VPWR VPWR _35103_/Q sky130_fd_sc_hd__dfxtp_1
X_32315_ _35580_/CLK _32315_/D VGND VGND VPWR VPWR _32315_/Q sky130_fd_sc_hd__dfxtp_1
X_17249_ _16994_/X _17247_/X _17248_/X _16997_/X VGND VGND VPWR VPWR _17249_/X sky130_fd_sc_hd__a22o_1
X_36083_ _36141_/CLK _36083_/D VGND VGND VPWR VPWR _36083_/Q sky130_fd_sc_hd__dfxtp_1
X_33295_ _33490_/CLK _33295_/D VGND VGND VPWR VPWR _33295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20260_ _20005_/X _20258_/X _20259_/X _20008_/X VGND VGND VPWR VPWR _20260_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35034_ _35034_/CLK _35034_/D VGND VGND VPWR VPWR _35034_/Q sky130_fd_sc_hd__dfxtp_1
X_32246_ _36150_/CLK _32246_/D VGND VGND VPWR VPWR _32246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20191_ _20187_/X _20190_/X _20153_/X VGND VGND VPWR VPWR _20199_/C sky130_fd_sc_hd__o21ba_1
XFILLER_66_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32177_ _36063_/CLK _32177_/D VGND VGND VPWR VPWR _32177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31128_ _35784_/Q _29231_/X _31130_/S VGND VGND VPWR VPWR _31129_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_111_CLK clkbuf_6_20__f_CLK/X VGND VGND VPWR VPWR _34638_/CLK sky130_fd_sc_hd__clkbuf_16
X_23950_ _23044_/X _32515_/Q _23962_/S VGND VGND VPWR VPWR _23951_/A sky130_fd_sc_hd__mux2_1
XTAP_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35936_ _35937_/CLK _35936_/D VGND VGND VPWR VPWR _35936_/Q sky130_fd_sc_hd__dfxtp_1
X_31059_ _35751_/Q _29129_/X _31067_/S VGND VGND VPWR VPWR _31060_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22901_ input62/X VGND VGND VPWR VPWR _22901_/X sky130_fd_sc_hd__buf_4
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35867_ _35931_/CLK _35867_/D VGND VGND VPWR VPWR _35867_/Q sky130_fd_sc_hd__dfxtp_1
X_23881_ _22941_/X _32482_/Q _23899_/S VGND VGND VPWR VPWR _23882_/A sky130_fd_sc_hd__mux2_1
X_25620_ _33238_/Q _24270_/X _25622_/S VGND VGND VPWR VPWR _25621_/A sky130_fd_sc_hd__mux2_1
X_34818_ _34819_/CLK _34818_/D VGND VGND VPWR VPWR _34818_/Q sky130_fd_sc_hd__dfxtp_1
X_22832_ _35596_/Q _35532_/Q _35468_/Q _35404_/Q _22556_/X _22557_/X VGND VGND VPWR
+ VPWR _22832_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35798_ _35799_/CLK _35798_/D VGND VGND VPWR VPWR _35798_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_908 _27018_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_919 _26996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_41__f_CLK clkbuf_5_20_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_41__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_225_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25551_ _25551_/A VGND VGND VPWR VPWR _33206_/D sky130_fd_sc_hd__clkbuf_1
X_22763_ _33290_/Q _36170_/Q _33162_/Q _33098_/Q _20628_/X _21757_/A VGND VGND VPWR
+ VPWR _22763_/X sky130_fd_sc_hd__mux4_1
X_34749_ _36029_/CLK _34749_/D VGND VGND VPWR VPWR _34749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24502_ _22963_/X _32745_/Q _24506_/S VGND VGND VPWR VPWR _24503_/A sky130_fd_sc_hd__mux2_1
X_21714_ _34539_/Q _32427_/Q _34411_/Q _34347_/Q _21472_/X _21473_/X VGND VGND VPWR
+ VPWR _21714_/X sky130_fd_sc_hd__mux4_1
X_28270_ _28270_/A VGND VGND VPWR VPWR _34460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25482_ _33174_/Q _24270_/X _25484_/S VGND VGND VPWR VPWR _25483_/A sky130_fd_sc_hd__mux2_1
X_22694_ _22694_/A VGND VGND VPWR VPWR _36231_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27221_ _26915_/X _33964_/Q _27239_/S VGND VGND VPWR VPWR _27222_/A sky130_fd_sc_hd__mux2_1
X_24433_ _24433_/A VGND VGND VPWR VPWR _32714_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_178_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _36107_/CLK sky130_fd_sc_hd__clkbuf_16
X_21645_ _21641_/X _21644_/X _21408_/X VGND VGND VPWR VPWR _21646_/D sky130_fd_sc_hd__o21ba_1
XFILLER_244_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27152_ _27014_/X _33932_/Q _27154_/S VGND VGND VPWR VPWR _27153_/A sky130_fd_sc_hd__mux2_1
X_24364_ _32692_/Q _24363_/X _24367_/S VGND VGND VPWR VPWR _24365_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_50 _32119_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21576_ _21576_/A _21576_/B _21576_/C _21576_/D VGND VGND VPWR VPWR _21577_/A sky130_fd_sc_hd__or4_4
XANTENNA_61 _32126_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_72 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26103_ _25128_/X _33466_/Q _26113_/S VGND VGND VPWR VPWR _26104_/A sky130_fd_sc_hd__mux2_1
X_23315_ _23315_/A VGND VGND VPWR VPWR _32222_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20527_ _19454_/A _20525_/X _20526_/X _19459_/A VGND VGND VPWR VPWR _20527_/X sky130_fd_sc_hd__a22o_1
XANTENNA_83 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27083_ _26912_/X _33899_/Q _27083_/S VGND VGND VPWR VPWR _27084_/A sky130_fd_sc_hd__mux2_1
XANTENNA_94 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24295_ input8/X VGND VGND VPWR VPWR _24295_/X sky130_fd_sc_hd__buf_4
XFILLER_21_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26034_ _25026_/X _33433_/Q _26050_/S VGND VGND VPWR VPWR _26035_/A sky130_fd_sc_hd__mux2_1
X_23246_ _23246_/A VGND VGND VPWR VPWR _32199_/D sky130_fd_sc_hd__clkbuf_1
X_20458_ _33546_/Q _33482_/Q _33418_/Q _33354_/Q _18333_/X _18335_/X VGND VGND VPWR
+ VPWR _20458_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_350_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _34291_/CLK sky130_fd_sc_hd__clkbuf_16
X_23177_ _23177_/A VGND VGND VPWR VPWR _32171_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20389_ _34567_/Q _32455_/Q _34439_/Q _34375_/Q _20231_/X _20232_/X VGND VGND VPWR
+ VPWR _20389_/X sky130_fd_sc_hd__mux4_1
XFILLER_234_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1307 _16990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1318 input45/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22128_ _32503_/Q _32375_/Q _32055_/Q _36023_/Q _21876_/X _22017_/X VGND VGND VPWR
+ VPWR _22128_/X sky130_fd_sc_hd__mux4_1
XTAP_6534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput190 _36216_/Q VGND VGND VPWR VPWR D2[42] sky130_fd_sc_hd__buf_2
XTAP_5800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27985_ _27985_/A VGND VGND VPWR VPWR _34325_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_1329 _20158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29724_ _29724_/A VGND VGND VPWR VPWR _35118_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_102_CLK clkbuf_leaf_99_CLK/A VGND VGND VPWR VPWR _35028_/CLK sky130_fd_sc_hd__clkbuf_16
X_26936_ _26936_/A VGND VGND VPWR VPWR _33842_/D sky130_fd_sc_hd__clkbuf_1
X_22059_ _21947_/X _22057_/X _22058_/X _21950_/X VGND VGND VPWR VPWR _22059_/X sky130_fd_sc_hd__a22o_1
XFILLER_82_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29655_ _29787_/S VGND VGND VPWR VPWR _29674_/S sky130_fd_sc_hd__buf_4
XFILLER_248_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26867_ _26866_/X _33820_/Q _26882_/S VGND VGND VPWR VPWR _26868_/A sky130_fd_sc_hd__mux2_1
XTAP_5899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28606_ _26965_/X _34620_/Q _28612_/S VGND VGND VPWR VPWR _28607_/A sky130_fd_sc_hd__mux2_1
X_16620_ _35037_/Q _34973_/Q _34909_/Q _34845_/Q _16450_/X _16451_/X VGND VGND VPWR
+ VPWR _16620_/X sky130_fd_sc_hd__mux4_1
X_25818_ _25106_/X _33331_/Q _25822_/S VGND VGND VPWR VPWR _25819_/A sky130_fd_sc_hd__mux2_1
X_26798_ _26798_/A VGND VGND VPWR VPWR _33794_/D sky130_fd_sc_hd__clkbuf_1
X_29586_ _35053_/Q _29148_/X _29602_/S VGND VGND VPWR VPWR _29587_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16551_ _35291_/Q _35227_/Q _35163_/Q _32283_/Q _16300_/X _16301_/X VGND VGND VPWR
+ VPWR _16551_/X sky130_fd_sc_hd__mux4_1
X_25749_ _25004_/X _33298_/Q _25759_/S VGND VGND VPWR VPWR _25750_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28537_ _26863_/X _34587_/Q _28549_/S VGND VGND VPWR VPWR _28538_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19270_ _35303_/Q _35239_/Q _35175_/Q _32295_/Q _18953_/X _18954_/X VGND VGND VPWR
+ VPWR _19270_/X sky130_fd_sc_hd__mux4_1
X_16482_ _16443_/X _16480_/X _16481_/X _16446_/X VGND VGND VPWR VPWR _16482_/X sky130_fd_sc_hd__a22o_1
X_28468_ _28468_/A VGND VGND VPWR VPWR _34554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18221_ _18217_/X _18220_/X _17834_/A VGND VGND VPWR VPWR _18243_/A sky130_fd_sc_hd__o21ba_1
X_27419_ _27419_/A VGND VGND VPWR VPWR _34058_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_169_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _36045_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28399_ _28399_/A VGND VGND VPWR VPWR _34521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30430_ _23294_/X _35453_/Q _30434_/S VGND VGND VPWR VPWR _30431_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18152_ _18148_/X _18151_/X _17867_/X VGND VGND VPWR VPWR _18153_/D sky130_fd_sc_hd__o21ba_1
XFILLER_178_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17103_ _17099_/X _17102_/X _16783_/X _16784_/X VGND VGND VPWR VPWR _17118_/B sky130_fd_sc_hd__o211a_1
X_18083_ _33223_/Q _32583_/Q _35975_/Q _35911_/Q _17780_/X _17781_/X VGND VGND VPWR
+ VPWR _18083_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30361_ _23130_/X _35420_/Q _30371_/S VGND VGND VPWR VPWR _30362_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17034_ _16994_/X _17032_/X _17033_/X _16997_/X VGND VGND VPWR VPWR _17034_/X sky130_fd_sc_hd__a22o_1
X_32100_ _35552_/CLK _32100_/D VGND VGND VPWR VPWR _32100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33080_ _36088_/CLK _33080_/D VGND VGND VPWR VPWR _33080_/Q sky130_fd_sc_hd__dfxtp_1
X_30292_ _35388_/Q _29194_/X _30298_/S VGND VGND VPWR VPWR _30293_/A sky130_fd_sc_hd__mux2_1
X_32031_ _36129_/CLK _32031_/D VGND VGND VPWR VPWR _32031_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_341_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _34039_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ _18981_/X _18984_/X _18741_/X VGND VGND VPWR VPWR _18993_/C sky130_fd_sc_hd__o21ba_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17936_ _17930_/X _17935_/X _17867_/X VGND VGND VPWR VPWR _17937_/D sky130_fd_sc_hd__o21ba_1
XFILLER_152_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33982_ _34046_/CLK _33982_/D VGND VGND VPWR VPWR _33982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35721_ _35848_/CLK _35721_/D VGND VGND VPWR VPWR _35721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32933_ _36069_/CLK _32933_/D VGND VGND VPWR VPWR _32933_/Q sky130_fd_sc_hd__dfxtp_1
X_17867_ _17867_/A VGND VGND VPWR VPWR _17867_/X sky130_fd_sc_hd__clkbuf_4
X_19606_ _32753_/Q _32689_/Q _32625_/Q _36081_/Q _19572_/X _19356_/X VGND VGND VPWR
+ VPWR _19606_/X sky130_fd_sc_hd__mux4_1
X_35652_ _35845_/CLK _35652_/D VGND VGND VPWR VPWR _35652_/Q sky130_fd_sc_hd__dfxtp_1
X_16818_ _16814_/X _16817_/X _16775_/X VGND VGND VPWR VPWR _16840_/A sky130_fd_sc_hd__o21ba_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32864_ _36001_/CLK _32864_/D VGND VGND VPWR VPWR _32864_/Q sky130_fd_sc_hd__dfxtp_1
X_17798_ _17548_/X _17794_/X _17797_/X _17553_/X VGND VGND VPWR VPWR _17798_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34603_ _34986_/CLK _34603_/D VGND VGND VPWR VPWR _34603_/Q sky130_fd_sc_hd__dfxtp_1
X_31815_ _31815_/A _31815_/B VGND VGND VPWR VPWR _31948_/S sky130_fd_sc_hd__nand2_8
X_19537_ _34031_/Q _33967_/Q _33903_/Q _32239_/Q _19320_/X _19321_/X VGND VGND VPWR
+ VPWR _19537_/X sky130_fd_sc_hd__mux4_1
X_35583_ _35583_/CLK _35583_/D VGND VGND VPWR VPWR _35583_/Q sky130_fd_sc_hd__dfxtp_1
X_16749_ _16710_/X _16747_/X _16748_/X _16714_/X VGND VGND VPWR VPWR _16749_/X sky130_fd_sc_hd__a22o_1
X_32795_ _36118_/CLK _32795_/D VGND VGND VPWR VPWR _32795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34534_ _35942_/CLK _34534_/D VGND VGND VPWR VPWR _34534_/Q sky130_fd_sc_hd__dfxtp_1
X_31746_ _31746_/A VGND VGND VPWR VPWR _36076_/D sky130_fd_sc_hd__clkbuf_1
X_19468_ _33517_/Q _33453_/Q _33389_/Q _33325_/Q _19423_/X _19424_/X VGND VGND VPWR
+ VPWR _19468_/X sky130_fd_sc_hd__mux4_2
XFILLER_59_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18419_ _18415_/X _18418_/X _18340_/X _18342_/X VGND VGND VPWR VPWR _18434_/B sky130_fd_sc_hd__o211a_1
XFILLER_222_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34465_ _35743_/CLK _34465_/D VGND VGND VPWR VPWR _34465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31677_ _31677_/A VGND VGND VPWR VPWR _36044_/D sky130_fd_sc_hd__clkbuf_1
X_19399_ _19355_/X _19397_/X _19398_/X _19361_/X VGND VGND VPWR VPWR _19399_/X sky130_fd_sc_hd__a22o_1
XFILLER_37_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36204_ _36204_/CLK _36204_/D VGND VGND VPWR VPWR _36204_/Q sky130_fd_sc_hd__dfxtp_1
X_33416_ _34306_/CLK _33416_/D VGND VGND VPWR VPWR _33416_/Q sky130_fd_sc_hd__dfxtp_1
X_21430_ _33187_/Q _32547_/Q _35939_/Q _35875_/Q _21321_/X _21322_/X VGND VGND VPWR
+ VPWR _21430_/X sky130_fd_sc_hd__mux4_1
X_30628_ _30628_/A VGND VGND VPWR VPWR _35546_/D sky130_fd_sc_hd__clkbuf_1
X_34396_ _35166_/CLK _34396_/D VGND VGND VPWR VPWR _34396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36135_ _36135_/CLK _36135_/D VGND VGND VPWR VPWR _36135_/Q sky130_fd_sc_hd__dfxtp_1
X_33347_ _34050_/CLK _33347_/D VGND VGND VPWR VPWR _33347_/Q sky130_fd_sc_hd__dfxtp_1
X_21361_ _34529_/Q _32417_/Q _34401_/Q _34337_/Q _21119_/X _21120_/X VGND VGND VPWR
+ VPWR _21361_/X sky130_fd_sc_hd__mux4_1
X_30559_ _23283_/X _35514_/Q _30569_/S VGND VGND VPWR VPWR _30560_/A sky130_fd_sc_hd__mux2_1
X_23100_ _32146_/Q _23099_/X _23115_/S VGND VGND VPWR VPWR _23101_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20312_ _32773_/Q _32709_/Q _32645_/Q _36101_/Q _20278_/X _20062_/X VGND VGND VPWR
+ VPWR _20312_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput70 R1[5] VGND VGND VPWR VPWR input70/X sky130_fd_sc_hd__buf_2
X_24080_ _23034_/X _32576_/Q _24098_/S VGND VGND VPWR VPWR _24081_/A sky130_fd_sc_hd__mux2_1
X_36066_ _36067_/CLK _36066_/D VGND VGND VPWR VPWR _36066_/Q sky130_fd_sc_hd__dfxtp_1
Xinput81 R3[4] VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__buf_2
X_33278_ _34046_/CLK _33278_/D VGND VGND VPWR VPWR _33278_/Q sky130_fd_sc_hd__dfxtp_1
X_21292_ _21288_/X _21291_/X _21055_/X VGND VGND VPWR VPWR _21293_/D sky130_fd_sc_hd__o21ba_1
X_35017_ _35781_/CLK _35017_/D VGND VGND VPWR VPWR _35017_/Q sky130_fd_sc_hd__dfxtp_1
X_23031_ input44/X VGND VGND VPWR VPWR _23031_/X sky130_fd_sc_hd__clkbuf_4
X_32229_ _35464_/CLK _32229_/D VGND VGND VPWR VPWR _32229_/Q sky130_fd_sc_hd__dfxtp_1
X_20243_ _34051_/Q _33987_/Q _33923_/Q _32259_/Q _20026_/X _20027_/X VGND VGND VPWR
+ VPWR _20243_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_332_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _36024_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20174_ _33537_/Q _33473_/Q _33409_/Q _33345_/Q _20129_/X _20130_/X VGND VGND VPWR
+ VPWR _20174_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1097 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24982_ _24982_/A VGND VGND VPWR VPWR _32970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27770_ _27770_/A VGND VGND VPWR VPWR _34223_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23933_ _23019_/X _32507_/Q _23941_/S VGND VGND VPWR VPWR _23934_/A sky130_fd_sc_hd__mux2_1
X_26721_ _33758_/Q _24295_/X _26727_/S VGND VGND VPWR VPWR _26722_/A sky130_fd_sc_hd__mux2_1
X_35919_ _35919_/CLK _35919_/D VGND VGND VPWR VPWR _35919_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26652_ _25140_/X _33726_/Q _26654_/S VGND VGND VPWR VPWR _26653_/A sky130_fd_sc_hd__mux2_1
XTAP_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29440_ _23223_/X _34984_/Q _29446_/S VGND VGND VPWR VPWR _29441_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23864_ _22917_/X _32474_/Q _23878_/S VGND VGND VPWR VPWR _23865_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_705 _22532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_716 _22453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25603_ _25735_/S VGND VGND VPWR VPWR _25622_/S sky130_fd_sc_hd__buf_4
XFILLER_84_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22815_ _33804_/Q _33740_/Q _33676_/Q _33612_/Q _20620_/X _20621_/X VGND VGND VPWR
+ VPWR _22815_/X sky130_fd_sc_hd__mux4_1
X_29371_ _29371_/A VGND VGND VPWR VPWR _34951_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_727 _20838_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_399_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _35500_/CLK sky130_fd_sc_hd__clkbuf_16
X_26583_ _25038_/X _33693_/Q _26591_/S VGND VGND VPWR VPWR _26584_/A sky130_fd_sc_hd__mux2_1
X_23795_ _23016_/X _32442_/Q _23805_/S VGND VGND VPWR VPWR _23796_/A sky130_fd_sc_hd__mux2_1
XANTENNA_738 _21545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_749 _22393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25534_ _25534_/A VGND VGND VPWR VPWR _33198_/D sky130_fd_sc_hd__clkbuf_1
X_28322_ _28322_/A VGND VGND VPWR VPWR _34485_/D sky130_fd_sc_hd__clkbuf_1
X_22746_ _34825_/Q _34761_/Q _34697_/Q _34633_/Q _22594_/X _22595_/X VGND VGND VPWR
+ VPWR _22746_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28253_ _28253_/A VGND VGND VPWR VPWR _34452_/D sky130_fd_sc_hd__clkbuf_1
X_25465_ _25597_/S VGND VGND VPWR VPWR _25484_/S sky130_fd_sc_hd__buf_4
X_22677_ _22369_/X _22675_/X _22676_/X _22373_/X VGND VGND VPWR VPWR _22677_/X sky130_fd_sc_hd__a22o_1
XFILLER_201_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27204_ _26891_/X _33956_/Q _27218_/S VGND VGND VPWR VPWR _27205_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24416_ input51/X VGND VGND VPWR VPWR _24416_/X sky130_fd_sc_hd__buf_4
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21628_ _32489_/Q _32361_/Q _32041_/Q _36009_/Q _21523_/X _21311_/X VGND VGND VPWR
+ VPWR _21628_/X sky130_fd_sc_hd__mux4_1
X_28184_ _26940_/X _34420_/Q _28186_/S VGND VGND VPWR VPWR _28185_/A sky130_fd_sc_hd__mux2_1
X_25396_ _25094_/X _33135_/Q _25408_/S VGND VGND VPWR VPWR _25397_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27135_ _27135_/A VGND VGND VPWR VPWR _33923_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24347_ _24347_/A VGND VGND VPWR VPWR _32686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21559_ _21555_/X _21558_/X _21383_/X _21384_/X VGND VGND VPWR VPWR _21576_/B sky130_fd_sc_hd__o211a_1
XFILLER_126_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27066_ _27066_/A VGND VGND VPWR VPWR _33890_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24278_ _32664_/Q _24276_/X _24305_/S VGND VGND VPWR VPWR _24279_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26017_ _25001_/X _33425_/Q _26029_/S VGND VGND VPWR VPWR _26018_/A sky130_fd_sc_hd__mux2_1
XTAP_7010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23229_ _32194_/Q _23228_/X _23235_/S VGND VGND VPWR VPWR _23230_/A sky130_fd_sc_hd__mux2_1
XTAP_7021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_323_CLK clkbuf_6_38__f_CLK/X VGND VGND VPWR VPWR _35956_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_7032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1104 _17400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1115 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1126 input63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1137 _18283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18770_ _32985_/Q _32921_/Q _32857_/Q _32793_/Q _18583_/X _18584_/X VGND VGND VPWR
+ VPWR _18770_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1148 _18789_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15982_ _16059_/A VGND VGND VPWR VPWR _17903_/A sky130_fd_sc_hd__buf_12
X_27968_ _27968_/A _28778_/B VGND VGND VPWR VPWR _28101_/S sky130_fd_sc_hd__nand2_8
XTAP_5630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1159 _22395_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29707_ _29707_/A VGND VGND VPWR VPWR _35110_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17721_ _17721_/A VGND VGND VPWR VPWR _31996_/D sky130_fd_sc_hd__clkbuf_4
X_26919_ input25/X VGND VGND VPWR VPWR _26919_/X sky130_fd_sc_hd__buf_4
XTAP_5674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27899_ _27899_/A VGND VGND VPWR VPWR _34284_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29638_ _35078_/Q _29225_/X _29644_/S VGND VGND VPWR VPWR _29639_/A sky130_fd_sc_hd__mux2_1
XTAP_4973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ _33787_/Q _33723_/Q _33659_/Q _33595_/Q _17549_/X _17550_/X VGND VGND VPWR
+ VPWR _17652_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16603_ _32477_/Q _32349_/Q _32029_/Q _35997_/Q _16570_/X _16358_/X VGND VGND VPWR
+ VPWR _16603_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17583_ _17577_/X _17582_/X _17514_/X VGND VGND VPWR VPWR _17584_/D sky130_fd_sc_hd__o21ba_1
X_29569_ _35045_/Q _29123_/X _29581_/S VGND VGND VPWR VPWR _29570_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31600_ _31600_/A VGND VGND VPWR VPWR _36007_/D sky130_fd_sc_hd__clkbuf_1
X_19322_ _34025_/Q _33961_/Q _33897_/Q _32226_/Q _19320_/X _19321_/X VGND VGND VPWR
+ VPWR _19322_/X sky130_fd_sc_hd__mux4_1
X_16534_ _32731_/Q _32667_/Q _32603_/Q _36059_/Q _16213_/X _16350_/X VGND VGND VPWR
+ VPWR _16534_/X sky130_fd_sc_hd__mux4_1
X_32580_ _35971_/CLK _32580_/D VGND VGND VPWR VPWR _32580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31531_ _23327_/X _35975_/Q _31535_/S VGND VGND VPWR VPWR _31532_/A sky130_fd_sc_hd__mux2_1
X_19253_ _32743_/Q _32679_/Q _32615_/Q _36071_/Q _19219_/X _19003_/X VGND VGND VPWR
+ VPWR _19253_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16465_ _16461_/X _16464_/X _16422_/X VGND VGND VPWR VPWR _16487_/A sky130_fd_sc_hd__o21ba_1
XFILLER_223_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18204_ _15997_/X _18202_/X _18203_/X _16003_/X VGND VGND VPWR VPWR _18204_/X sky130_fd_sc_hd__a22o_1
XPHY_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34250_ _35851_/CLK _34250_/D VGND VGND VPWR VPWR _34250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16396_ _16357_/X _16394_/X _16395_/X _16361_/X VGND VGND VPWR VPWR _16396_/X sky130_fd_sc_hd__a22o_1
X_31462_ _23217_/X _35942_/Q _31472_/S VGND VGND VPWR VPWR _31463_/A sky130_fd_sc_hd__mux2_1
X_19184_ _34021_/Q _33957_/Q _33893_/Q _32182_/Q _18967_/X _18968_/X VGND VGND VPWR
+ VPWR _19184_/X sky130_fd_sc_hd__mux4_1
XPHY_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33201_ _35889_/CLK _33201_/D VGND VGND VPWR VPWR _33201_/Q sky130_fd_sc_hd__dfxtp_1
X_18135_ _32521_/Q _32393_/Q _32073_/Q _36041_/Q _17982_/X _17007_/A VGND VGND VPWR
+ VPWR _18135_/X sky130_fd_sc_hd__mux4_1
X_30413_ _23267_/X _35445_/Q _30413_/S VGND VGND VPWR VPWR _30414_/A sky130_fd_sc_hd__mux2_1
X_34181_ _34308_/CLK _34181_/D VGND VGND VPWR VPWR _34181_/Q sky130_fd_sc_hd__dfxtp_1
X_31393_ _31393_/A VGND VGND VPWR VPWR _35909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33132_ _36141_/CLK _33132_/D VGND VGND VPWR VPWR _33132_/Q sky130_fd_sc_hd__dfxtp_1
X_18066_ _34311_/Q _34247_/Q _34183_/Q _34119_/Q _17795_/X _17796_/X VGND VGND VPWR
+ VPWR _18066_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30344_ _23105_/X _35412_/Q _30350_/S VGND VGND VPWR VPWR _30345_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_5__f_CLK clkbuf_5_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_5__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_17017_ _34281_/Q _34217_/Q _34153_/Q _34089_/Q _16736_/X _16737_/X VGND VGND VPWR
+ VPWR _17017_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_314_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _34809_/CLK sky130_fd_sc_hd__clkbuf_16
X_30275_ _35380_/Q _29169_/X _30277_/S VGND VGND VPWR VPWR _30276_/A sky130_fd_sc_hd__mux2_1
X_33063_ _36135_/CLK _33063_/D VGND VGND VPWR VPWR _33063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32014_ _35982_/CLK _32014_/D VGND VGND VPWR VPWR _32014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18968_ _20147_/A VGND VGND VPWR VPWR _18968_/X sky130_fd_sc_hd__buf_4
XFILLER_101_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17919_ _17769_/X _17917_/X _17918_/X _17773_/X VGND VGND VPWR VPWR _17919_/X sky130_fd_sc_hd__a22o_1
XFILLER_152_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33965_ _35958_/CLK _33965_/D VGND VGND VPWR VPWR _33965_/Q sky130_fd_sc_hd__dfxtp_1
X_18899_ _18895_/X _18898_/X _18722_/X VGND VGND VPWR VPWR _18923_/A sky130_fd_sc_hd__o21ba_1
XFILLER_227_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35704_ _35766_/CLK _35704_/D VGND VGND VPWR VPWR _35704_/Q sky130_fd_sc_hd__dfxtp_1
X_20930_ _33173_/Q _32533_/Q _35925_/Q _35861_/Q _20663_/X _20665_/X VGND VGND VPWR
+ VPWR _20930_/X sky130_fd_sc_hd__mux4_1
X_32916_ _35002_/CLK _32916_/D VGND VGND VPWR VPWR _32916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33896_ _34153_/CLK _33896_/D VGND VGND VPWR VPWR _33896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35635_ _35827_/CLK _35635_/D VGND VGND VPWR VPWR _35635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20861_ _20656_/X _20859_/X _20860_/X _20668_/X VGND VGND VPWR VPWR _20861_/X sky130_fd_sc_hd__a22o_1
X_32847_ _35985_/CLK _32847_/D VGND VGND VPWR VPWR _32847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22600_ _35076_/Q _35012_/Q _34948_/Q _34884_/Q _22462_/X _22463_/X VGND VGND VPWR
+ VPWR _22600_/X sky130_fd_sc_hd__mux4_1
XFILLER_207_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23580_ _23580_/A VGND VGND VPWR VPWR _32341_/D sky130_fd_sc_hd__clkbuf_1
X_35566_ _35949_/CLK _35566_/D VGND VGND VPWR VPWR _35566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32778_ _36172_/CLK _32778_/D VGND VGND VPWR VPWR _32778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20792_ _22447_/A VGND VGND VPWR VPWR _20792_/X sky130_fd_sc_hd__buf_4
XFILLER_81_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22531_ _22531_/A VGND VGND VPWR VPWR _22531_/X sky130_fd_sc_hd__buf_6
X_34517_ _36196_/CLK _34517_/D VGND VGND VPWR VPWR _34517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_928 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31729_ _31729_/A VGND VGND VPWR VPWR _36068_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35497_ _35819_/CLK _35497_/D VGND VGND VPWR VPWR _35497_/Q sky130_fd_sc_hd__dfxtp_1
X_25250_ _25250_/A VGND VGND VPWR VPWR _33066_/D sky130_fd_sc_hd__clkbuf_1
X_22462_ _22462_/A VGND VGND VPWR VPWR _22462_/X sky130_fd_sc_hd__buf_4
XFILLER_206_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34448_ _35279_/CLK _34448_/D VGND VGND VPWR VPWR _34448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24201_ _23013_/X _32633_/Q _24213_/S VGND VGND VPWR VPWR _24202_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21413_ _34275_/Q _34211_/Q _34147_/Q _34083_/Q _21336_/X _21337_/X VGND VGND VPWR
+ VPWR _21413_/X sky130_fd_sc_hd__mux4_1
X_25181_ _25180_/X _33035_/Q _25187_/S VGND VGND VPWR VPWR _25182_/A sky130_fd_sc_hd__mux2_1
X_34379_ _35147_/CLK _34379_/D VGND VGND VPWR VPWR _34379_/Q sky130_fd_sc_hd__dfxtp_1
X_22393_ _22393_/A VGND VGND VPWR VPWR _36222_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36118_ _36118_/CLK _36118_/D VGND VGND VPWR VPWR _36118_/Q sky130_fd_sc_hd__dfxtp_1
X_24132_ _22910_/X _32600_/Q _24150_/S VGND VGND VPWR VPWR _24133_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21344_ _32737_/Q _32673_/Q _32609_/Q _36065_/Q _21166_/X _21303_/X VGND VGND VPWR
+ VPWR _21344_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36049_ _36049_/CLK _36049_/D VGND VGND VPWR VPWR _36049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24063_ _23010_/X _32568_/Q _24077_/S VGND VGND VPWR VPWR _24064_/A sky130_fd_sc_hd__mux2_1
X_28940_ _34778_/Q _24283_/X _28954_/S VGND VGND VPWR VPWR _28941_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_305_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _34620_/CLK sky130_fd_sc_hd__clkbuf_16
X_21275_ _32479_/Q _32351_/Q _32031_/Q _35999_/Q _21170_/X _20958_/X VGND VGND VPWR
+ VPWR _21275_/X sky130_fd_sc_hd__mux4_1
X_23014_ _23013_/X _32057_/Q _23032_/S VGND VGND VPWR VPWR _23015_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20226_ _20005_/X _20224_/X _20225_/X _20008_/X VGND VGND VPWR VPWR _20226_/X sky130_fd_sc_hd__a22o_1
XFILLER_172_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28871_ _28871_/A VGND VGND VPWR VPWR _34745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27822_ _27822_/A VGND VGND VPWR VPWR _34248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20157_ _35328_/Q _35264_/Q _35200_/Q _32320_/Q _20012_/X _20013_/X VGND VGND VPWR
+ VPWR _20157_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24965_ _23041_/X _32962_/Q _24979_/S VGND VGND VPWR VPWR _24966_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27753_ _27753_/A VGND VGND VPWR VPWR _34215_/D sky130_fd_sc_hd__clkbuf_1
X_20088_ _34558_/Q _32446_/Q _34430_/Q _34366_/Q _19878_/X _19879_/X VGND VGND VPWR
+ VPWR _20088_/X sky130_fd_sc_hd__mux4_1
XTAP_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26704_ _33750_/Q _24270_/X _26706_/S VGND VGND VPWR VPWR _26705_/A sky130_fd_sc_hd__mux2_1
XTAP_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23916_ _22994_/X _32499_/Q _23920_/S VGND VGND VPWR VPWR _23917_/A sky130_fd_sc_hd__mux2_1
X_27684_ _34183_/Q _24422_/X _27688_/S VGND VGND VPWR VPWR _27685_/A sky130_fd_sc_hd__mux2_1
XTAP_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24896_ _24896_/A VGND VGND VPWR VPWR _32929_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_502 _17792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29423_ _23142_/X _34976_/Q _29425_/S VGND VGND VPWR VPWR _29424_/A sky130_fd_sc_hd__mux2_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_513 _17938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26635_ _26683_/S VGND VGND VPWR VPWR _26654_/S sky130_fd_sc_hd__buf_4
X_23847_ _22892_/X _32466_/Q _23857_/S VGND VGND VPWR VPWR _23848_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_524 _18004_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_535 _20095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_546 _20162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29354_ _29354_/A VGND VGND VPWR VPWR _34943_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_557 _20295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26566_ _25013_/X _33685_/Q _26570_/S VGND VGND VPWR VPWR _26567_/A sky130_fd_sc_hd__mux2_1
XANTENNA_568 _20147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23778_ _22991_/X _32434_/Q _23784_/S VGND VGND VPWR VPWR _23779_/A sky130_fd_sc_hd__mux2_1
XANTENNA_579 _20153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28305_ _34477_/Q _24342_/X _28321_/S VGND VGND VPWR VPWR _28306_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22729_ _34057_/Q _33993_/Q _33929_/Q _32265_/Q _20658_/X _20660_/X VGND VGND VPWR
+ VPWR _22729_/X sky130_fd_sc_hd__mux4_1
XFILLER_214_895 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25517_ _25517_/A VGND VGND VPWR VPWR _33190_/D sky130_fd_sc_hd__clkbuf_1
X_29285_ _29285_/A VGND VGND VPWR VPWR _34910_/D sky130_fd_sc_hd__clkbuf_1
X_26497_ _25112_/X _33653_/Q _26497_/S VGND VGND VPWR VPWR _26498_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16250_ _32467_/Q _32339_/Q _32019_/Q _35987_/Q _16217_/X _17863_/A VGND VGND VPWR
+ VPWR _16250_/X sky130_fd_sc_hd__mux4_1
X_28236_ _27017_/X _34445_/Q _28236_/S VGND VGND VPWR VPWR _28237_/A sky130_fd_sc_hd__mux2_1
X_25448_ _25171_/X _33160_/Q _25450_/S VGND VGND VPWR VPWR _25449_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16181_ _32721_/Q _32657_/Q _32593_/Q _36049_/Q _17862_/A _17713_/A VGND VGND VPWR
+ VPWR _16181_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28167_ _28236_/S VGND VGND VPWR VPWR _28186_/S sky130_fd_sc_hd__buf_4
X_25379_ _25069_/X _33127_/Q _25387_/S VGND VGND VPWR VPWR _25380_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27118_ _27118_/A VGND VGND VPWR VPWR _33915_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28098_ _28098_/A VGND VGND VPWR VPWR _34379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19940_ _19936_/X _19939_/X _19800_/X VGND VGND VPWR VPWR _19950_/C sky130_fd_sc_hd__o21ba_1
XFILLER_114_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27049_ _27049_/A VGND VGND VPWR VPWR _33882_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30060_ _30192_/S VGND VGND VPWR VPWR _30079_/S sky130_fd_sc_hd__buf_6
XFILLER_141_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19871_ _35576_/Q _35512_/Q _35448_/Q _35384_/Q _19550_/X _19551_/X VGND VGND VPWR
+ VPWR _19871_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18822_ _35034_/Q _34970_/Q _34906_/Q _34842_/Q _18750_/X _18751_/X VGND VGND VPWR
+ VPWR _18822_/X sky130_fd_sc_hd__mux4_1
XTAP_6150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18753_ _19459_/A VGND VGND VPWR VPWR _18753_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_95_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17704_ _17700_/X _17701_/X _17702_/X _17703_/X VGND VGND VPWR VPWR _17704_/X sky130_fd_sc_hd__a22o_1
X_33750_ _34259_/CLK _33750_/D VGND VGND VPWR VPWR _33750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18684_ _20257_/A VGND VGND VPWR VPWR _18684_/X sky130_fd_sc_hd__buf_4
X_30962_ _35705_/Q _29185_/X _30974_/S VGND VGND VPWR VPWR _30963_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32701_ _36095_/CLK _32701_/D VGND VGND VPWR VPWR _32701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17635_ _35770_/Q _35130_/Q _34490_/Q _33850_/Q _17493_/X _17494_/X VGND VGND VPWR
+ VPWR _17635_/X sky130_fd_sc_hd__mux4_1
X_33681_ _34194_/CLK _33681_/D VGND VGND VPWR VPWR _33681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30893_ _35672_/Q _29082_/X _30911_/S VGND VGND VPWR VPWR _30894_/A sky130_fd_sc_hd__mux2_1
X_35420_ _35869_/CLK _35420_/D VGND VGND VPWR VPWR _35420_/Q sky130_fd_sc_hd__dfxtp_1
X_32632_ _36089_/CLK _32632_/D VGND VGND VPWR VPWR _32632_/Q sky130_fd_sc_hd__dfxtp_1
X_17566_ _17416_/X _17564_/X _17565_/X _17420_/X VGND VGND VPWR VPWR _17566_/X sky130_fd_sc_hd__a22o_1
XFILLER_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19305_ _34792_/Q _34728_/Q _34664_/Q _34600_/Q _19235_/X _19236_/X VGND VGND VPWR
+ VPWR _19305_/X sky130_fd_sc_hd__mux4_1
XFILLER_205_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35351_ _35863_/CLK _35351_/D VGND VGND VPWR VPWR _35351_/Q sky130_fd_sc_hd__dfxtp_1
X_16517_ _35290_/Q _35226_/Q _35162_/Q _32282_/Q _16300_/X _16301_/X VGND VGND VPWR
+ VPWR _16517_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32563_ _35955_/CLK _32563_/D VGND VGND VPWR VPWR _32563_/Q sky130_fd_sc_hd__dfxtp_1
X_17497_ _35574_/Q _35510_/Q _35446_/Q _35382_/Q _17250_/X _17251_/X VGND VGND VPWR
+ VPWR _17497_/X sky130_fd_sc_hd__mux4_1
XFILLER_231_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34302_ _34302_/CLK _34302_/D VGND VGND VPWR VPWR _34302_/Q sky130_fd_sc_hd__dfxtp_1
X_31514_ _23300_/X _35967_/Q _31514_/S VGND VGND VPWR VPWR _31515_/A sky130_fd_sc_hd__mux2_1
X_19236_ _20295_/A VGND VGND VPWR VPWR _19236_/X sky130_fd_sc_hd__clkbuf_4
X_35282_ _35282_/CLK _35282_/D VGND VGND VPWR VPWR _35282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16448_ _17154_/A VGND VGND VPWR VPWR _16448_/X sky130_fd_sc_hd__buf_4
XFILLER_158_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1069 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32494_ _36015_/CLK _32494_/D VGND VGND VPWR VPWR _32494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34233_ _34296_/CLK _34233_/D VGND VGND VPWR VPWR _34233_/Q sky130_fd_sc_hd__dfxtp_1
X_31445_ _23136_/X _35934_/Q _31451_/S VGND VGND VPWR VPWR _31446_/A sky130_fd_sc_hd__mux2_1
X_19167_ _18946_/X _19165_/X _19166_/X _18949_/X VGND VGND VPWR VPWR _19167_/X sky130_fd_sc_hd__a22o_1
X_16379_ _16375_/X _16378_/X _16100_/X VGND VGND VPWR VPWR _16380_/D sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_91_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _36191_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18118_ _17855_/X _18116_/X _18117_/X _17858_/X VGND VGND VPWR VPWR _18118_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34164_ _34228_/CLK _34164_/D VGND VGND VPWR VPWR _34164_/Q sky130_fd_sc_hd__dfxtp_1
X_31376_ _31376_/A VGND VGND VPWR VPWR _35901_/D sky130_fd_sc_hd__clkbuf_1
X_19098_ _35298_/Q _35234_/Q _35170_/Q _32290_/Q _18953_/X _18954_/X VGND VGND VPWR
+ VPWR _19098_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33115_ _34265_/CLK _33115_/D VGND VGND VPWR VPWR _33115_/Q sky130_fd_sc_hd__dfxtp_1
X_30327_ _35405_/Q _29246_/X _30327_/S VGND VGND VPWR VPWR _30328_/A sky130_fd_sc_hd__mux2_1
X_18049_ _35846_/Q _32225_/Q _35718_/Q _35654_/Q _15989_/X _15991_/X VGND VGND VPWR
+ VPWR _18049_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34095_ _34286_/CLK _34095_/D VGND VGND VPWR VPWR _34095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33046_ _36117_/CLK _33046_/D VGND VGND VPWR VPWR _33046_/Q sky130_fd_sc_hd__dfxtp_1
X_21060_ _34265_/Q _34201_/Q _34137_/Q _34073_/Q _20983_/X _20984_/X VGND VGND VPWR
+ VPWR _21060_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_1162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30258_ _30327_/S VGND VGND VPWR VPWR _30277_/S sky130_fd_sc_hd__buf_6
XFILLER_63_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20011_ _34812_/Q _34748_/Q _34684_/Q _34620_/Q _19941_/X _19942_/X VGND VGND VPWR
+ VPWR _20011_/X sky130_fd_sc_hd__mux4_1
X_30189_ _30189_/A VGND VGND VPWR VPWR _35339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34997_ _34997_/CLK _34997_/D VGND VGND VPWR VPWR _34997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24750_ _22923_/X _32860_/Q _24760_/S VGND VGND VPWR VPWR _24751_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21962_ _21749_/X _21958_/X _21961_/X _21752_/X VGND VGND VPWR VPWR _21962_/X sky130_fd_sc_hd__a22o_1
X_33948_ _34205_/CLK _33948_/D VGND VGND VPWR VPWR _33948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23701_ _28778_/B _30465_/B VGND VGND VPWR VPWR _23834_/S sky130_fd_sc_hd__nand2_8
XFILLER_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20913_ _33493_/Q _33429_/Q _33365_/Q _33301_/Q _20598_/X _20599_/X VGND VGND VPWR
+ VPWR _20913_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24681_ _24681_/A VGND VGND VPWR VPWR _32828_/D sky130_fd_sc_hd__clkbuf_1
X_33879_ _36220_/CLK _33879_/D VGND VGND VPWR VPWR _33879_/Q sky130_fd_sc_hd__dfxtp_1
X_21893_ _34544_/Q _32432_/Q _34416_/Q _34352_/Q _21825_/X _21826_/X VGND VGND VPWR
+ VPWR _21893_/X sky130_fd_sc_hd__mux4_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26420_ _24998_/X _33616_/Q _26434_/S VGND VGND VPWR VPWR _26421_/A sky130_fd_sc_hd__mux2_1
X_35618_ _35811_/CLK _35618_/D VGND VGND VPWR VPWR _35618_/Q sky130_fd_sc_hd__dfxtp_1
X_23632_ _32366_/Q _23244_/X _23646_/S VGND VGND VPWR VPWR _23633_/A sky130_fd_sc_hd__mux2_1
X_20844_ _34003_/Q _33939_/Q _33875_/Q _32147_/Q _20708_/X _20709_/X VGND VGND VPWR
+ VPWR _20844_/X sky130_fd_sc_hd__mux4_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_20_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_20_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_214_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26351_ _26351_/A VGND VGND VPWR VPWR _33583_/D sky130_fd_sc_hd__clkbuf_1
X_23563_ _31680_/B _25462_/A VGND VGND VPWR VPWR _23696_/S sky130_fd_sc_hd__nor2_8
X_35549_ _35935_/CLK _35549_/D VGND VGND VPWR VPWR _35549_/Q sky130_fd_sc_hd__dfxtp_1
X_20775_ _34257_/Q _34193_/Q _34129_/Q _34065_/Q _20605_/X _20607_/X VGND VGND VPWR
+ VPWR _20775_/X sky130_fd_sc_hd__mux4_1
XFILLER_243_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25302_ _25156_/X _33091_/Q _25314_/S VGND VGND VPWR VPWR _25303_/A sky130_fd_sc_hd__mux2_1
X_22514_ _32770_/Q _32706_/Q _32642_/Q _36098_/Q _22225_/X _22362_/X VGND VGND VPWR
+ VPWR _22514_/X sky130_fd_sc_hd__mux4_1
X_26282_ _26282_/A VGND VGND VPWR VPWR _33550_/D sky130_fd_sc_hd__clkbuf_1
X_29070_ input61/X VGND VGND VPWR VPWR _29070_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23494_ _23494_/A VGND VGND VPWR VPWR _32301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28021_ _28021_/A VGND VGND VPWR VPWR _34342_/D sky130_fd_sc_hd__clkbuf_1
X_25233_ _25053_/X _33058_/Q _25251_/S VGND VGND VPWR VPWR _25234_/A sky130_fd_sc_hd__mux2_1
X_22445_ _35840_/Q _32219_/Q _35712_/Q _35648_/Q _22266_/X _22267_/X VGND VGND VPWR
+ VPWR _22445_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_82_CLK clkbuf_leaf_87_CLK/A VGND VGND VPWR VPWR _35797_/CLK sky130_fd_sc_hd__clkbuf_16
X_25164_ _25164_/A VGND VGND VPWR VPWR _33029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22376_ _35838_/Q _32217_/Q _35710_/Q _35646_/Q _22266_/X _22267_/X VGND VGND VPWR
+ VPWR _22376_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24115_ _22886_/X _32592_/Q _24129_/S VGND VGND VPWR VPWR _24116_/A sky130_fd_sc_hd__mux2_1
X_21327_ _35296_/Q _35232_/Q _35168_/Q _32288_/Q _21253_/X _21254_/X VGND VGND VPWR
+ VPWR _21327_/X sky130_fd_sc_hd__mux4_1
X_25095_ _25094_/X _33007_/Q _25113_/S VGND VGND VPWR VPWR _25096_/A sky130_fd_sc_hd__mux2_1
X_29972_ _35236_/Q _29120_/X _29986_/S VGND VGND VPWR VPWR _29973_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28923_ _34770_/Q _24258_/X _28933_/S VGND VGND VPWR VPWR _28924_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24046_ _22985_/X _32560_/Q _24056_/S VGND VGND VPWR VPWR _24047_/A sky130_fd_sc_hd__mux2_1
X_21258_ _35038_/Q _34974_/Q _34910_/Q _34846_/Q _21050_/X _21051_/X VGND VGND VPWR
+ VPWR _21258_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20209_ _33538_/Q _33474_/Q _33410_/Q _33346_/Q _20129_/X _20130_/X VGND VGND VPWR
+ VPWR _20209_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28854_ _28854_/A VGND VGND VPWR VPWR _34737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21189_ _21048_/X _21187_/X _21188_/X _21053_/X VGND VGND VPWR VPWR _21189_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_948 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27805_ _34240_/Q _24400_/X _27823_/S VGND VGND VPWR VPWR _27806_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28785_ _28785_/A VGND VGND VPWR VPWR _34704_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25997_ _25171_/X _33416_/Q _25999_/S VGND VGND VPWR VPWR _25998_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_1262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27736_ _27736_/A VGND VGND VPWR VPWR _34207_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24948_ _23016_/X _32954_/Q _24958_/S VGND VGND VPWR VPWR _24949_/A sky130_fd_sc_hd__mux2_1
XTAP_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_310 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27667_ _34175_/Q _24397_/X _27667_/S VGND VGND VPWR VPWR _27668_/A sky130_fd_sc_hd__mux2_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24879_ _22914_/X _32921_/Q _24895_/S VGND VGND VPWR VPWR _24880_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_321 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_332 _32141_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29406_ _29517_/S VGND VGND VPWR VPWR _29425_/S sky130_fd_sc_hd__buf_4
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _17911_/A VGND VGND VPWR VPWR _17420_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_343 _36205_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26618_ _26618_/A VGND VGND VPWR VPWR _33709_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_354 _36206_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_365 _36207_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27598_ _34142_/Q _24295_/X _27604_/S VGND VGND VPWR VPWR _27599_/A sky130_fd_sc_hd__mux2_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_376 _36208_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29337_ _23274_/X _34935_/Q _29353_/S VGND VGND VPWR VPWR _29338_/A sky130_fd_sc_hd__mux2_1
XANTENNA_387 _36209_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _17347_/X _17348_/X _17349_/X _17350_/X VGND VGND VPWR VPWR _17351_/X sky130_fd_sc_hd__a22o_1
X_26549_ input85/X input84/X _26549_/C VGND VGND VPWR VPWR _31815_/A sky130_fd_sc_hd__nor3_4
XANTENNA_398 _36210_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _35284_/Q _35220_/Q _35156_/Q _32276_/Q _16300_/X _16301_/X VGND VGND VPWR
+ VPWR _16302_/X sky130_fd_sc_hd__mux4_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29268_ _29268_/A VGND VGND VPWR VPWR _34902_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17282_ _35760_/Q _35120_/Q _34480_/Q _33840_/Q _17140_/X _17141_/X VGND VGND VPWR
+ VPWR _17282_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19021_ _20231_/A VGND VGND VPWR VPWR _19021_/X sky130_fd_sc_hd__buf_6
X_28219_ _28219_/A VGND VGND VPWR VPWR _34436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16233_ _16074_/X _16231_/X _16232_/X _16084_/X VGND VGND VPWR VPWR _16233_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29199_ _29199_/A VGND VGND VPWR VPWR _34877_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_73_CLK clkbuf_leaf_73_CLK/A VGND VGND VPWR VPWR _36050_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_103_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31230_ _35832_/Q input37/X _31244_/S VGND VGND VPWR VPWR _31231_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16164_ _35280_/Q _35216_/Q _35152_/Q _32272_/Q _16079_/X _16081_/X VGND VGND VPWR
+ VPWR _16164_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_18__f_CLK clkbuf_5_9_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_87_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_86_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1075 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16095_ _35022_/Q _34958_/Q _34894_/Q _34830_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _16095_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31161_ _31161_/A VGND VGND VPWR VPWR _35799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19923_ _19855_/X _19921_/X _19922_/X _19858_/X VGND VGND VPWR VPWR _19923_/X sky130_fd_sc_hd__a22o_1
X_30112_ _30112_/A VGND VGND VPWR VPWR _35302_/D sky130_fd_sc_hd__clkbuf_1
X_31092_ _31092_/A VGND VGND VPWR VPWR _35766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30043_ _35270_/Q _29225_/X _30049_/S VGND VGND VPWR VPWR _30044_/A sky130_fd_sc_hd__mux2_1
X_34920_ _35302_/CLK _34920_/D VGND VGND VPWR VPWR _34920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19854_ _19848_/X _19851_/X _19852_/X _19853_/X VGND VGND VPWR VPWR _19854_/X sky130_fd_sc_hd__a22o_1
XFILLER_218_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18805_ _32474_/Q _32346_/Q _32026_/Q _35994_/Q _18517_/X _18658_/X VGND VGND VPWR
+ VPWR _18805_/X sky130_fd_sc_hd__mux4_1
XFILLER_205_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34851_ _35299_/CLK _34851_/D VGND VGND VPWR VPWR _34851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19785_ _19708_/X _19783_/X _19784_/X _19714_/X VGND VGND VPWR VPWR _19785_/X sky130_fd_sc_hd__a22o_1
X_16997_ _17858_/A VGND VGND VPWR VPWR _16997_/X sky130_fd_sc_hd__buf_4
XFILLER_37_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33802_ _34251_/CLK _33802_/D VGND VGND VPWR VPWR _33802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18736_ _35736_/Q _35096_/Q _34456_/Q _33816_/Q _18734_/X _18735_/X VGND VGND VPWR
+ VPWR _18736_/X sky130_fd_sc_hd__mux4_1
XTAP_5290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34782_ _34782_/CLK _34782_/D VGND VGND VPWR VPWR _34782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31994_ _34205_/CLK _31994_/D VGND VGND VPWR VPWR _31994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33733_ _34308_/CLK _33733_/D VGND VGND VPWR VPWR _33733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18667_ _35542_/Q _35478_/Q _35414_/Q _35350_/Q _18491_/X _18492_/X VGND VGND VPWR
+ VPWR _18667_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30945_ _35697_/Q _29160_/X _30953_/S VGND VGND VPWR VPWR _30946_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17618_ _33786_/Q _33722_/Q _33658_/Q _33594_/Q _17549_/X _17550_/X VGND VGND VPWR
+ VPWR _17618_/X sky130_fd_sc_hd__mux4_1
X_33664_ _33729_/CLK _33664_/D VGND VGND VPWR VPWR _33664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30876_ _35664_/Q _29058_/X _30890_/S VGND VGND VPWR VPWR _30877_/A sky130_fd_sc_hd__mux2_1
X_18598_ _18592_/X _18597_/X _18371_/X VGND VGND VPWR VPWR _18608_/C sky130_fd_sc_hd__o21ba_1
XFILLER_225_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35403_ _35851_/CLK _35403_/D VGND VGND VPWR VPWR _35403_/Q sky130_fd_sc_hd__dfxtp_1
X_32615_ _33255_/CLK _32615_/D VGND VGND VPWR VPWR _32615_/Q sky130_fd_sc_hd__dfxtp_1
X_17549_ _17902_/A VGND VGND VPWR VPWR _17549_/X sky130_fd_sc_hd__buf_4
X_33595_ _33723_/CLK _33595_/D VGND VGND VPWR VPWR _33595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35334_ _35334_/CLK _35334_/D VGND VGND VPWR VPWR _35334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20560_ _35789_/Q _35149_/Q _34509_/Q _33869_/Q _18408_/X _18409_/X VGND VGND VPWR
+ VPWR _20560_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32546_ _35298_/CLK _32546_/D VGND VGND VPWR VPWR _32546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19219_ _20278_/A VGND VGND VPWR VPWR _19219_/X sky130_fd_sc_hd__buf_8
X_35265_ _35328_/CLK _35265_/D VGND VGND VPWR VPWR _35265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20491_ _20487_/X _20490_/X _20134_/A VGND VGND VPWR VPWR _20513_/A sky130_fd_sc_hd__o21ba_1
XFILLER_203_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32477_ _34146_/CLK _32477_/D VGND VGND VPWR VPWR _32477_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_64_CLK clkbuf_leaf_66_CLK/A VGND VGND VPWR VPWR _33507_/CLK sky130_fd_sc_hd__clkbuf_16
X_22230_ _32506_/Q _32378_/Q _32058_/Q _36026_/Q _22229_/X _22017_/X VGND VGND VPWR
+ VPWR _22230_/X sky130_fd_sc_hd__mux4_1
X_34216_ _34279_/CLK _34216_/D VGND VGND VPWR VPWR _34216_/Q sky130_fd_sc_hd__dfxtp_1
X_31428_ _23111_/X _35926_/Q _31430_/S VGND VGND VPWR VPWR _31429_/A sky130_fd_sc_hd__mux2_1
X_35196_ _35583_/CLK _35196_/D VGND VGND VPWR VPWR _35196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22161_ _32760_/Q _32696_/Q _32632_/Q _36088_/Q _21872_/X _22009_/X VGND VGND VPWR
+ VPWR _22161_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34147_ _35992_/CLK _34147_/D VGND VGND VPWR VPWR _34147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31359_ _31359_/A VGND VGND VPWR VPWR _35893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21112_ _35546_/Q _35482_/Q _35418_/Q _35354_/Q _20791_/X _20792_/X VGND VGND VPWR
+ VPWR _21112_/X sky130_fd_sc_hd__mux4_1
XFILLER_246_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34078_ _36200_/CLK _34078_/D VGND VGND VPWR VPWR _34078_/Q sky130_fd_sc_hd__dfxtp_1
X_22092_ _35830_/Q _32208_/Q _35702_/Q _35638_/Q _21913_/X _21914_/X VGND VGND VPWR
+ VPWR _22092_/X sky130_fd_sc_hd__mux4_1
XTAP_6919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33029_ _36100_/CLK _33029_/D VGND VGND VPWR VPWR _33029_/Q sky130_fd_sc_hd__dfxtp_1
X_25920_ _25057_/X _33379_/Q _25936_/S VGND VGND VPWR VPWR _25921_/A sky130_fd_sc_hd__mux2_1
X_21043_ _21749_/A VGND VGND VPWR VPWR _21043_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25851_ _25851_/A VGND VGND VPWR VPWR _33346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24802_ _23000_/X _32885_/Q _24802_/S VGND VGND VPWR VPWR _24803_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28570_ _26912_/X _34603_/Q _28570_/S VGND VGND VPWR VPWR _28571_/A sky130_fd_sc_hd__mux2_1
X_25782_ _25872_/S VGND VGND VPWR VPWR _25801_/S sky130_fd_sc_hd__buf_4
X_22994_ input31/X VGND VGND VPWR VPWR _22994_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_210_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27521_ _27521_/A VGND VGND VPWR VPWR _34106_/D sky130_fd_sc_hd__clkbuf_1
X_24733_ _22898_/X _32852_/Q _24739_/S VGND VGND VPWR VPWR _24734_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21945_ _21663_/X _21941_/X _21944_/X _21667_/X VGND VGND VPWR VPWR _21945_/X sky130_fd_sc_hd__a22o_1
XFILLER_216_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27452_ _27452_/A VGND VGND VPWR VPWR _34073_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24664_ _24664_/A VGND VGND VPWR VPWR _32820_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21876_ _22582_/A VGND VGND VPWR VPWR _21876_/X sky130_fd_sc_hd__buf_6
XFILLER_242_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26403_ _26403_/A VGND VGND VPWR VPWR _33608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23615_ _32358_/Q _23217_/X _23625_/S VGND VGND VPWR VPWR _23616_/A sky130_fd_sc_hd__mux2_1
X_20827_ _20656_/X _20825_/X _20826_/X _20668_/X VGND VGND VPWR VPWR _20827_/X sky130_fd_sc_hd__a22o_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24595_ _24595_/A VGND VGND VPWR VPWR _32787_/D sky130_fd_sc_hd__clkbuf_1
X_27383_ _34041_/Q _24379_/X _27395_/S VGND VGND VPWR VPWR _27384_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29122_ _29122_/A VGND VGND VPWR VPWR _34852_/D sky130_fd_sc_hd__clkbuf_1
X_23546_ _23546_/A VGND VGND VPWR VPWR _32326_/D sky130_fd_sc_hd__clkbuf_1
X_26334_ _26334_/A VGND VGND VPWR VPWR _33575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20758_ _20644_/X _20756_/X _20757_/X _20654_/X VGND VGND VPWR VPWR _20758_/X sky130_fd_sc_hd__a22o_1
XFILLER_211_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26265_ _25168_/X _33543_/Q _26269_/S VGND VGND VPWR VPWR _26266_/A sky130_fd_sc_hd__mux2_1
X_29053_ _34830_/Q _29048_/X _29080_/S VGND VGND VPWR VPWR _29054_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23477_ _23477_/A VGND VGND VPWR VPWR _32293_/D sky130_fd_sc_hd__clkbuf_1
X_20689_ _22362_/A VGND VGND VPWR VPWR _21473_/A sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_55_CLK clkbuf_leaf_57_CLK/A VGND VGND VPWR VPWR _33635_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28004_ _28004_/A VGND VGND VPWR VPWR _34334_/D sky130_fd_sc_hd__clkbuf_1
X_25216_ _25029_/X _33050_/Q _25230_/S VGND VGND VPWR VPWR _25217_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22428_ _22148_/X _22426_/X _22427_/X _22153_/X VGND VGND VPWR VPWR _22428_/X sky130_fd_sc_hd__a22o_1
XFILLER_137_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26196_ _25066_/X _33510_/Q _26206_/S VGND VGND VPWR VPWR _26197_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25147_ _25187_/S VGND VGND VPWR VPWR _25175_/S sky130_fd_sc_hd__buf_6
XFILLER_13_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22359_ _22155_/X _22357_/X _22358_/X _22158_/X VGND VGND VPWR VPWR _22359_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1048 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29955_ _35228_/Q _29095_/X _29965_/S VGND VGND VPWR VPWR _29956_/A sky130_fd_sc_hd__mux2_1
X_25078_ input21/X VGND VGND VPWR VPWR _25078_/X sky130_fd_sc_hd__buf_2
XFILLER_3_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28906_ _28906_/A VGND VGND VPWR VPWR _34762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24029_ _22960_/X _32552_/Q _24035_/S VGND VGND VPWR VPWR _24030_/A sky130_fd_sc_hd__mux2_1
X_16920_ _32742_/Q _32678_/Q _32614_/Q _36070_/Q _16919_/X _16703_/X VGND VGND VPWR
+ VPWR _16920_/X sky130_fd_sc_hd__mux4_1
X_29886_ _29886_/A VGND VGND VPWR VPWR _35195_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28837_ _28837_/A VGND VGND VPWR VPWR _34729_/D sky130_fd_sc_hd__clkbuf_1
X_16851_ _34020_/Q _33956_/Q _33892_/Q _32171_/Q _16667_/X _16668_/X VGND VGND VPWR
+ VPWR _16851_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_1046 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19570_ _19502_/X _19568_/X _19569_/X _19505_/X VGND VGND VPWR VPWR _19570_/X sky130_fd_sc_hd__a22o_1
X_28768_ _27005_/X _34697_/Q _28768_/S VGND VGND VPWR VPWR _28769_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16782_ _16710_/X _16780_/X _16781_/X _16714_/X VGND VGND VPWR VPWR _16782_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18521_ _18516_/X _18520_/X _18340_/X _18342_/X VGND VGND VPWR VPWR _18538_/B sky130_fd_sc_hd__o211a_1
XFILLER_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27719_ _27719_/A VGND VGND VPWR VPWR _34199_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28699_ _26903_/X _34664_/Q _28705_/S VGND VGND VPWR VPWR _28700_/A sky130_fd_sc_hd__mux2_1
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30730_ _30730_/A VGND VGND VPWR VPWR _35595_/D sky130_fd_sc_hd__clkbuf_1
X_18452_ _32464_/Q _32336_/Q _32016_/Q _35984_/Q _18328_/X _20163_/A VGND VGND VPWR
+ VPWR _18452_/X sky130_fd_sc_hd__mux4_1
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_151 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_162 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17403_ _17195_/X _17401_/X _17402_/X _17200_/X VGND VGND VPWR VPWR _17403_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_173 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18383_ _20067_/A VGND VGND VPWR VPWR _19452_/A sky130_fd_sc_hd__buf_12
XFILLER_18_1112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30661_ _30661_/A VGND VGND VPWR VPWR _35562_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_195 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32400_ _35281_/CLK _32400_/D VGND VGND VPWR VPWR _32400_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _33522_/Q _33458_/Q _33394_/Q _33330_/Q _17123_/X _17124_/X VGND VGND VPWR
+ VPWR _17334_/X sky130_fd_sc_hd__mux4_1
X_33380_ _33702_/CLK _33380_/D VGND VGND VPWR VPWR _33380_/Q sky130_fd_sc_hd__dfxtp_1
X_30592_ _23336_/X _35530_/Q _30598_/S VGND VGND VPWR VPWR _30593_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32331_ _35147_/CLK _32331_/D VGND VGND VPWR VPWR _32331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17265_ _33776_/Q _33712_/Q _33648_/Q _33584_/Q _17196_/X _17197_/X VGND VGND VPWR
+ VPWR _17265_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_CLK clkbuf_6_6__f_CLK/X VGND VGND VPWR VPWR _35481_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19004_ _32736_/Q _32672_/Q _32608_/Q _36064_/Q _18866_/X _19003_/X VGND VGND VPWR
+ VPWR _19004_/X sky130_fd_sc_hd__mux4_1
X_16216_ _16014_/X _16214_/X _16215_/X _16023_/X VGND VGND VPWR VPWR _16216_/X sky130_fd_sc_hd__a22o_1
X_35050_ _35050_/CLK _35050_/D VGND VGND VPWR VPWR _35050_/Q sky130_fd_sc_hd__dfxtp_1
X_32262_ _34306_/CLK _32262_/D VGND VGND VPWR VPWR _32262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17196_ _17902_/A VGND VGND VPWR VPWR _17196_/X sky130_fd_sc_hd__buf_4
X_34001_ _34001_/CLK _34001_/D VGND VGND VPWR VPWR _34001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31213_ _35824_/Q input28/X _31223_/S VGND VGND VPWR VPWR _31214_/A sky130_fd_sc_hd__mux2_1
X_16147_ _16143_/X _16144_/X _16145_/X _16146_/X VGND VGND VPWR VPWR _16147_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32193_ _34087_/CLK _32193_/D VGND VGND VPWR VPWR _32193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31144_ _35791_/Q input12/X _31160_/S VGND VGND VPWR VPWR _31145_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16078_ _17978_/A VGND VGND VPWR VPWR _17712_/A sky130_fd_sc_hd__buf_12
XFILLER_64_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19906_ _33209_/Q _32569_/Q _35961_/Q _35897_/Q _19727_/X _19728_/X VGND VGND VPWR
+ VPWR _19906_/X sky130_fd_sc_hd__mux4_1
X_31075_ _31075_/A VGND VGND VPWR VPWR _35758_/D sky130_fd_sc_hd__clkbuf_1
X_35952_ _35952_/CLK _35952_/D VGND VGND VPWR VPWR _35952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34903_ _34967_/CLK _34903_/D VGND VGND VPWR VPWR _34903_/Q sky130_fd_sc_hd__dfxtp_1
X_30026_ _35262_/Q _29200_/X _30028_/S VGND VGND VPWR VPWR _30027_/A sky130_fd_sc_hd__mux2_1
X_19837_ _19652_/X _19835_/X _19836_/X _19655_/X VGND VGND VPWR VPWR _19837_/X sky130_fd_sc_hd__a22o_1
X_35883_ _35947_/CLK _35883_/D VGND VGND VPWR VPWR _35883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34834_ _35026_/CLK _34834_/D VGND VGND VPWR VPWR _34834_/Q sky130_fd_sc_hd__dfxtp_1
Xinput2 DW[10] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__buf_6
X_19768_ _35061_/Q _34997_/Q _34933_/Q _34869_/Q _19456_/X _19457_/X VGND VGND VPWR
+ VPWR _19768_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18719_ _33496_/Q _33432_/Q _33368_/Q _33304_/Q _18717_/X _18718_/X VGND VGND VPWR
+ VPWR _18719_/X sky130_fd_sc_hd__mux4_1
X_34765_ _35341_/CLK _34765_/D VGND VGND VPWR VPWR _34765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31977_ _35293_/CLK _31977_/D VGND VGND VPWR VPWR _31977_/Q sky130_fd_sc_hd__dfxtp_1
X_19699_ _19699_/A _19699_/B _19699_/C _19699_/D VGND VGND VPWR VPWR _19700_/A sky130_fd_sc_hd__or4_2
XFILLER_232_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21730_ _32748_/Q _32684_/Q _32620_/Q _36076_/Q _21519_/X _21656_/X VGND VGND VPWR
+ VPWR _21730_/X sky130_fd_sc_hd__mux4_1
X_33716_ _33780_/CLK _33716_/D VGND VGND VPWR VPWR _33716_/Q sky130_fd_sc_hd__dfxtp_1
X_30928_ _35689_/Q _29135_/X _30932_/S VGND VGND VPWR VPWR _30929_/A sky130_fd_sc_hd__mux2_1
X_34696_ _35334_/CLK _34696_/D VGND VGND VPWR VPWR _34696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33647_ _33775_/CLK _33647_/D VGND VGND VPWR VPWR _33647_/Q sky130_fd_sc_hd__dfxtp_1
X_21661_ _22506_/A VGND VGND VPWR VPWR _21661_/X sky130_fd_sc_hd__buf_6
XFILLER_240_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30859_ _30859_/A VGND VGND VPWR VPWR _35656_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23400_ _23400_/A VGND VGND VPWR VPWR _32258_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20612_ _20593_/X _20609_/X _20611_/X VGND VGND VPWR VPWR _20702_/A sky130_fd_sc_hd__o21ba_1
XFILLER_51_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24380_ _32697_/Q _24379_/X _24398_/S VGND VGND VPWR VPWR _24381_/A sky130_fd_sc_hd__mux2_1
X_33578_ _34281_/CLK _33578_/D VGND VGND VPWR VPWR _33578_/Q sky130_fd_sc_hd__dfxtp_1
X_21592_ _21310_/X _21588_/X _21591_/X _21314_/X VGND VGND VPWR VPWR _21592_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23331_ _32228_/Q _23330_/X _23334_/S VGND VGND VPWR VPWR _23332_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35317_ _35574_/CLK _35317_/D VGND VGND VPWR VPWR _35317_/Q sky130_fd_sc_hd__dfxtp_1
X_20543_ _20543_/A _20543_/B _20543_/C _20543_/D VGND VGND VPWR VPWR _20544_/A sky130_fd_sc_hd__or4_1
X_32529_ _34317_/CLK _32529_/D VGND VGND VPWR VPWR _32529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_37_CLK clkbuf_6_7__f_CLK/X VGND VGND VPWR VPWR _36123_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_192_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26050_ _25050_/X _33441_/Q _26050_/S VGND VGND VPWR VPWR _26051_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35248_ _35757_/CLK _35248_/D VGND VGND VPWR VPWR _35248_/Q sky130_fd_sc_hd__dfxtp_1
X_23262_ _32205_/Q _23261_/X _23268_/S VGND VGND VPWR VPWR _23263_/A sky130_fd_sc_hd__mux2_1
X_20474_ _18297_/X _20472_/X _20473_/X _18303_/X VGND VGND VPWR VPWR _20474_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25001_ input34/X VGND VGND VPWR VPWR _25001_/X sky130_fd_sc_hd__buf_4
XFILLER_69_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22213_ _35065_/Q _35001_/Q _34937_/Q _34873_/Q _22109_/X _22110_/X VGND VGND VPWR
+ VPWR _22213_/X sky130_fd_sc_hd__mux4_1
XFILLER_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35179_ _35179_/CLK _35179_/D VGND VGND VPWR VPWR _35179_/Q sky130_fd_sc_hd__dfxtp_1
X_23193_ _32179_/Q _23130_/X _23206_/S VGND VGND VPWR VPWR _23194_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22144_ _22107_/X _22142_/X _22143_/X _22112_/X VGND VGND VPWR VPWR _22144_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29740_ _35126_/Q _29175_/X _29758_/S VGND VGND VPWR VPWR _29741_/A sky130_fd_sc_hd__mux2_1
XTAP_6738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26952_ _26952_/A VGND VGND VPWR VPWR _33847_/D sky130_fd_sc_hd__clkbuf_1
X_22075_ _21795_/X _22073_/X _22074_/X _21800_/X VGND VGND VPWR VPWR _22075_/X sky130_fd_sc_hd__a22o_1
XFILLER_248_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25903_ _25032_/X _33371_/Q _25915_/S VGND VGND VPWR VPWR _25904_/A sky130_fd_sc_hd__mux2_1
X_21026_ _20949_/X _21024_/X _21025_/X _20955_/X VGND VGND VPWR VPWR _21026_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29671_ _29671_/A VGND VGND VPWR VPWR _35093_/D sky130_fd_sc_hd__clkbuf_1
X_26883_ _26883_/A VGND VGND VPWR VPWR _33825_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28622_ _28622_/A VGND VGND VPWR VPWR _34627_/D sky130_fd_sc_hd__clkbuf_1
X_25834_ _25834_/A VGND VGND VPWR VPWR _33338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28553_ _28553_/A VGND VGND VPWR VPWR _34594_/D sky130_fd_sc_hd__clkbuf_1
X_25765_ _25765_/A VGND VGND VPWR VPWR _33305_/D sky130_fd_sc_hd__clkbuf_1
X_22977_ _22976_/X _32045_/Q _23001_/S VGND VGND VPWR VPWR _22978_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27504_ _27504_/A VGND VGND VPWR VPWR _34098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1014 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24716_ _24716_/A VGND VGND VPWR VPWR _32845_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28484_ _26984_/X _34562_/Q _28498_/S VGND VGND VPWR VPWR _28485_/A sky130_fd_sc_hd__mux2_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21928_ _21924_/X _21927_/X _21761_/X VGND VGND VPWR VPWR _21929_/D sky130_fd_sc_hd__o21ba_1
X_25696_ _33274_/Q _24382_/X _25706_/S VGND VGND VPWR VPWR _25697_/A sky130_fd_sc_hd__mux2_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27435_ _27435_/A VGND VGND VPWR VPWR _34065_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24647_ _22972_/X _32812_/Q _24665_/S VGND VGND VPWR VPWR _24648_/A sky130_fd_sc_hd__mux2_1
X_21859_ _34543_/Q _32431_/Q _34415_/Q _34351_/Q _21825_/X _21826_/X VGND VGND VPWR
+ VPWR _21859_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27366_ _34033_/Q _24354_/X _27374_/S VGND VGND VPWR VPWR _27367_/A sky130_fd_sc_hd__mux2_1
X_24578_ _24578_/A VGND VGND VPWR VPWR _32781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29105_ _34847_/Q _29104_/X _29111_/S VGND VGND VPWR VPWR _29106_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26317_ _26317_/A VGND VGND VPWR VPWR _33567_/D sky130_fd_sc_hd__clkbuf_1
X_23529_ _23529_/A VGND VGND VPWR VPWR _32318_/D sky130_fd_sc_hd__clkbuf_1
X_27297_ _34000_/Q _24252_/X _27311_/S VGND VGND VPWR VPWR _27298_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_28_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _33946_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29036_ _34824_/Q _24425_/X _29038_/S VGND VGND VPWR VPWR _29037_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17050_ _16842_/X _17048_/X _17049_/X _16847_/X VGND VGND VPWR VPWR _17050_/X sky130_fd_sc_hd__a22o_1
X_26248_ _25143_/X _33535_/Q _26248_/S VGND VGND VPWR VPWR _26249_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16001_ input68/X input67/X VGND VGND VPWR VPWR _17773_/A sky130_fd_sc_hd__nor2b_4
XFILLER_87_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1023 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26179_ _25041_/X _33502_/Q _26185_/S VGND VGND VPWR VPWR _26180_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17952_ _17948_/X _17951_/X _17842_/X _17843_/X VGND VGND VPWR VPWR _17969_/B sky130_fd_sc_hd__o211a_1
XFILLER_151_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29938_ _35220_/Q _29070_/X _29944_/S VGND VGND VPWR VPWR _29939_/A sky130_fd_sc_hd__mux2_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16903_ _34789_/Q _34725_/Q _34661_/Q _34597_/Q _16582_/X _16583_/X VGND VGND VPWR
+ VPWR _16903_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17883_ _17769_/X _17881_/X _17882_/X _17773_/X VGND VGND VPWR VPWR _17883_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_918 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29869_ _29869_/A VGND VGND VPWR VPWR _35187_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31900_ _31948_/S VGND VGND VPWR VPWR _31919_/S sky130_fd_sc_hd__buf_4
X_19622_ _34801_/Q _34737_/Q _34673_/Q _34609_/Q _19588_/X _19589_/X VGND VGND VPWR
+ VPWR _19622_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16834_ _35299_/Q _35235_/Q _35171_/Q _32291_/Q _16653_/X _16654_/X VGND VGND VPWR
+ VPWR _16834_/X sky130_fd_sc_hd__mux4_1
X_32880_ _33009_/CLK _32880_/D VGND VGND VPWR VPWR _32880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31831_ _23108_/X _36117_/Q _31835_/S VGND VGND VPWR VPWR _31832_/A sky130_fd_sc_hd__mux2_1
X_19553_ _33199_/Q _32559_/Q _35951_/Q _35887_/Q _19374_/X _19375_/X VGND VGND VPWR
+ VPWR _19553_/X sky130_fd_sc_hd__mux4_1
XFILLER_24_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16765_ _16765_/A _16765_/B _16765_/C _16765_/D VGND VGND VPWR VPWR _16766_/A sky130_fd_sc_hd__or4_1
XFILLER_98_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18504_ _18504_/A _18504_/B _18504_/C _18504_/D VGND VGND VPWR VPWR _18505_/A sky130_fd_sc_hd__or4_4
X_34550_ _35768_/CLK _34550_/D VGND VGND VPWR VPWR _34550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19484_ _19299_/X _19482_/X _19483_/X _19302_/X VGND VGND VPWR VPWR _19484_/X sky130_fd_sc_hd__a22o_1
X_31762_ _31762_/A VGND VGND VPWR VPWR _36084_/D sky130_fd_sc_hd__clkbuf_1
X_16696_ _34272_/Q _34208_/Q _34144_/Q _34080_/Q _16383_/X _16384_/X VGND VGND VPWR
+ VPWR _16696_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33501_ _34202_/CLK _33501_/D VGND VGND VPWR VPWR _33501_/Q sky130_fd_sc_hd__dfxtp_1
X_30713_ _35587_/Q _29216_/X _30725_/S VGND VGND VPWR VPWR _30714_/A sky130_fd_sc_hd__mux2_1
X_18435_ _18435_/A VGND VGND VPWR VPWR _32079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34481_ _35760_/CLK _34481_/D VGND VGND VPWR VPWR _34481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31693_ _31693_/A VGND VGND VPWR VPWR _36051_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36220_ _36220_/CLK _36220_/D VGND VGND VPWR VPWR _36220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33432_ _34267_/CLK _33432_/D VGND VGND VPWR VPWR _33432_/Q sky130_fd_sc_hd__dfxtp_1
X_18366_ _33166_/Q _32526_/Q _35918_/Q _35854_/Q _18363_/X _18365_/X VGND VGND VPWR
+ VPWR _18366_/X sky130_fd_sc_hd__mux4_1
X_30644_ _35554_/Q _29113_/X _30662_/S VGND VGND VPWR VPWR _30645_/A sky130_fd_sc_hd__mux2_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36151_ _36152_/CLK _36151_/D VGND VGND VPWR VPWR _36151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17317_ _16994_/X _17315_/X _17316_/X _16997_/X VGND VGND VPWR VPWR _17317_/X sky130_fd_sc_hd__a22o_1
X_33363_ _36232_/CLK _33363_/D VGND VGND VPWR VPWR _33363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18297_ _20160_/A VGND VGND VPWR VPWR _18297_/X sky130_fd_sc_hd__buf_4
XFILLER_187_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30575_ _30575_/A VGND VGND VPWR VPWR _35521_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_19_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _34777_/CLK sky130_fd_sc_hd__clkbuf_16
X_35102_ _35743_/CLK _35102_/D VGND VGND VPWR VPWR _35102_/Q sky130_fd_sc_hd__dfxtp_1
X_32314_ _35577_/CLK _32314_/D VGND VGND VPWR VPWR _32314_/Q sky130_fd_sc_hd__dfxtp_1
X_17248_ _35759_/Q _35119_/Q _34479_/Q _33839_/Q _17140_/X _17141_/X VGND VGND VPWR
+ VPWR _17248_/X sky130_fd_sc_hd__mux4_1
X_36082_ _36141_/CLK _36082_/D VGND VGND VPWR VPWR _36082_/Q sky130_fd_sc_hd__dfxtp_1
X_33294_ _33490_/CLK _33294_/D VGND VGND VPWR VPWR _33294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35033_ _35034_/CLK _35033_/D VGND VGND VPWR VPWR _35033_/Q sky130_fd_sc_hd__dfxtp_1
X_32245_ _36149_/CLK _32245_/D VGND VGND VPWR VPWR _32245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17179_ _35821_/Q _32198_/Q _35693_/Q _35629_/Q _16960_/X _16961_/X VGND VGND VPWR
+ VPWR _17179_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20190_ _20005_/X _20188_/X _20189_/X _20008_/X VGND VGND VPWR VPWR _20190_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32176_ _36063_/CLK _32176_/D VGND VGND VPWR VPWR _32176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31127_ _31127_/A VGND VGND VPWR VPWR _35783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35935_ _35935_/CLK _35935_/D VGND VGND VPWR VPWR _35935_/Q sky130_fd_sc_hd__dfxtp_1
X_31058_ _31058_/A VGND VGND VPWR VPWR _35750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22900_ _22900_/A VGND VGND VPWR VPWR _32020_/D sky130_fd_sc_hd__clkbuf_1
X_30009_ _30057_/S VGND VGND VPWR VPWR _30028_/S sky130_fd_sc_hd__buf_4
XFILLER_29_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23880_ _23970_/S VGND VGND VPWR VPWR _23899_/S sky130_fd_sc_hd__buf_4
XTAP_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35866_ _35931_/CLK _35866_/D VGND VGND VPWR VPWR _35866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22831_ _20577_/X _22829_/X _22830_/X _20587_/X VGND VGND VPWR VPWR _22831_/X sky130_fd_sc_hd__a22o_1
X_34817_ _34817_/CLK _34817_/D VGND VGND VPWR VPWR _34817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35797_ _35797_/CLK _35797_/D VGND VGND VPWR VPWR _35797_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_909 _27018_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22762_ _32778_/Q _32714_/Q _32650_/Q _36106_/Q _22578_/X _21473_/A VGND VGND VPWR
+ VPWR _22762_/X sky130_fd_sc_hd__mux4_1
XFILLER_112_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25550_ _33206_/Q _24369_/X _25568_/S VGND VGND VPWR VPWR _25551_/A sky130_fd_sc_hd__mux2_1
X_34748_ _35707_/CLK _34748_/D VGND VGND VPWR VPWR _34748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21713_ _21396_/X _21711_/X _21712_/X _21399_/X VGND VGND VPWR VPWR _21713_/X sky130_fd_sc_hd__a22o_1
X_24501_ _24501_/A VGND VGND VPWR VPWR _32744_/D sky130_fd_sc_hd__clkbuf_1
X_25481_ _25481_/A VGND VGND VPWR VPWR _33173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22693_ _22693_/A _22693_/B _22693_/C _22693_/D VGND VGND VPWR VPWR _22694_/A sky130_fd_sc_hd__or4_4
XFILLER_227_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34679_ _34745_/CLK _34679_/D VGND VGND VPWR VPWR _34679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27220_ _27289_/S VGND VGND VPWR VPWR _27239_/S sky130_fd_sc_hd__buf_4
XFILLER_244_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24432_ _32714_/Q _24431_/X _24441_/S VGND VGND VPWR VPWR _24433_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21644_ _21401_/X _21642_/X _21643_/X _21406_/X VGND VGND VPWR VPWR _21644_/X sky130_fd_sc_hd__a22o_1
XFILLER_36_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27151_ _27151_/A VGND VGND VPWR VPWR _33931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24363_ input32/X VGND VGND VPWR VPWR _24363_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_40 _32118_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21575_ _21571_/X _21574_/X _21408_/X VGND VGND VPWR VPWR _21576_/D sky130_fd_sc_hd__o21ba_1
XFILLER_240_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_51 _32119_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23314_ _32222_/Q _23313_/X _23334_/S VGND VGND VPWR VPWR _23315_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26102_ _26102_/A VGND VGND VPWR VPWR _33465_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_62 _32126_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20526_ _33036_/Q _32972_/Q _32908_/Q _32844_/Q _18280_/X _18283_/X VGND VGND VPWR
+ VPWR _20526_/X sky130_fd_sc_hd__mux4_1
XANTENNA_73 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27082_ _27082_/A VGND VGND VPWR VPWR _33898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_84 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24294_ _24294_/A VGND VGND VPWR VPWR _32669_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_95 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26033_ _26033_/A VGND VGND VPWR VPWR _33432_/D sky130_fd_sc_hd__clkbuf_1
X_23245_ _32199_/Q _23244_/X _23268_/S VGND VGND VPWR VPWR _23246_/A sky130_fd_sc_hd__mux2_1
X_20457_ _20201_/X _20455_/X _20456_/X _20206_/X VGND VGND VPWR VPWR _20457_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23176_ _32171_/Q _23175_/X _23350_/S VGND VGND VPWR VPWR _23177_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20388_ _20155_/X _20386_/X _20387_/X _20158_/X VGND VGND VPWR VPWR _20388_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22127_ _22008_/X _22125_/X _22126_/X _22014_/X VGND VGND VPWR VPWR _22127_/X sky130_fd_sc_hd__a22o_1
XTAP_6524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1308 _17055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1319 input52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27984_ _26844_/X _34325_/Q _27988_/S VGND VGND VPWR VPWR _27985_/A sky130_fd_sc_hd__mux2_1
XTAP_6546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput180 _36207_/Q VGND VGND VPWR VPWR D2[33] sky130_fd_sc_hd__buf_2
Xoutput191 _36217_/Q VGND VGND VPWR VPWR D2[43] sky130_fd_sc_hd__buf_2
XTAP_5812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29723_ _35118_/Q _29151_/X _29737_/S VGND VGND VPWR VPWR _29724_/A sky130_fd_sc_hd__mux2_1
XTAP_6568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26935_ _26934_/X _33842_/Q _26944_/S VGND VGND VPWR VPWR _26936_/A sky130_fd_sc_hd__mux2_1
X_22058_ _35765_/Q _35125_/Q _34485_/Q _33845_/Q _21740_/X _21741_/X VGND VGND VPWR
+ VPWR _22058_/X sky130_fd_sc_hd__mux4_1
XTAP_6579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21009_ _35031_/Q _34967_/Q _34903_/Q _34839_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _21009_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29654_ _29924_/A _31275_/B VGND VGND VPWR VPWR _29787_/S sky130_fd_sc_hd__nor2_8
XTAP_5867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26866_ input6/X VGND VGND VPWR VPWR _26866_/X sky130_fd_sc_hd__buf_4
XTAP_5889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28605_ _28605_/A VGND VGND VPWR VPWR _34619_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25817_ _25817_/A VGND VGND VPWR VPWR _33330_/D sky130_fd_sc_hd__clkbuf_1
X_29585_ _29585_/A VGND VGND VPWR VPWR _35052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26797_ _33794_/Q _24407_/X _26811_/S VGND VGND VPWR VPWR _26798_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28536_ _28536_/A VGND VGND VPWR VPWR _34586_/D sky130_fd_sc_hd__clkbuf_1
X_16550_ _34779_/Q _34715_/Q _34651_/Q _34587_/Q _16229_/X _16230_/X VGND VGND VPWR
+ VPWR _16550_/X sky130_fd_sc_hd__mux4_1
X_25748_ _25748_/A VGND VGND VPWR VPWR _33297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28467_ _26959_/X _34554_/Q _28477_/S VGND VGND VPWR VPWR _28468_/A sky130_fd_sc_hd__mux2_1
X_16481_ _35289_/Q _35225_/Q _35161_/Q _32281_/Q _16300_/X _16301_/X VGND VGND VPWR
+ VPWR _16481_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25679_ _33266_/Q _24357_/X _25685_/S VGND VGND VPWR VPWR _25680_/A sky130_fd_sc_hd__mux2_1
X_18220_ _16026_/X _18218_/X _18219_/X _16037_/X VGND VGND VPWR VPWR _18220_/X sky130_fd_sc_hd__a22o_1
X_27418_ _34058_/Q _24431_/X _27424_/S VGND VGND VPWR VPWR _27419_/A sky130_fd_sc_hd__mux2_1
X_28398_ _26857_/X _34521_/Q _28414_/S VGND VGND VPWR VPWR _28399_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18151_ _17860_/X _18149_/X _18150_/X _17865_/X VGND VGND VPWR VPWR _18151_/X sky130_fd_sc_hd__a22o_1
XFILLER_141_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27349_ _34025_/Q _24329_/X _27353_/S VGND VGND VPWR VPWR _27350_/A sky130_fd_sc_hd__mux2_1
X_17102_ _17063_/X _17100_/X _17101_/X _17067_/X VGND VGND VPWR VPWR _17102_/X sky130_fd_sc_hd__a22o_1
XFILLER_129_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18082_ _35591_/Q _35527_/Q _35463_/Q _35399_/Q _17956_/X _17957_/X VGND VGND VPWR
+ VPWR _18082_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30360_ _30360_/A VGND VGND VPWR VPWR _35419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29019_ _29046_/S VGND VGND VPWR VPWR _29038_/S sky130_fd_sc_hd__buf_4
X_17033_ _35753_/Q _35113_/Q _34473_/Q _33833_/Q _16787_/X _16788_/X VGND VGND VPWR
+ VPWR _17033_/X sky130_fd_sc_hd__mux4_1
X_30291_ _30291_/A VGND VGND VPWR VPWR _35387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32030_ _36065_/CLK _32030_/D VGND VGND VPWR VPWR _32030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ _18946_/X _18982_/X _18983_/X _18949_/X VGND VGND VPWR VPWR _18984_/X sky130_fd_sc_hd__a22o_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ _17860_/X _17933_/X _17934_/X _17865_/X VGND VGND VPWR VPWR _17935_/X sky130_fd_sc_hd__a22o_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33981_ _34046_/CLK _33981_/D VGND VGND VPWR VPWR _33981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35720_ _35848_/CLK _35720_/D VGND VGND VPWR VPWR _35720_/Q sky130_fd_sc_hd__dfxtp_1
X_32932_ _36067_/CLK _32932_/D VGND VGND VPWR VPWR _32932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17866_ _17860_/X _17861_/X _17864_/X _17865_/X VGND VGND VPWR VPWR _17866_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _35164_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1040 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19605_ _19601_/X _19604_/X _19428_/X VGND VGND VPWR VPWR _19629_/A sky130_fd_sc_hd__o21ba_1
X_16817_ _16496_/X _16815_/X _16816_/X _16499_/X VGND VGND VPWR VPWR _16817_/X sky130_fd_sc_hd__a22o_1
X_35651_ _35845_/CLK _35651_/D VGND VGND VPWR VPWR _35651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32863_ _36062_/CLK _32863_/D VGND VGND VPWR VPWR _32863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17797_ _34303_/Q _34239_/Q _34175_/Q _34111_/Q _17795_/X _17796_/X VGND VGND VPWR
+ VPWR _17797_/X sky130_fd_sc_hd__mux4_1
X_31814_ _31814_/A VGND VGND VPWR VPWR _36109_/D sky130_fd_sc_hd__clkbuf_1
X_19536_ _33519_/Q _33455_/Q _33391_/Q _33327_/Q _19423_/X _19424_/X VGND VGND VPWR
+ VPWR _19536_/X sky130_fd_sc_hd__mux4_1
X_34602_ _34794_/CLK _34602_/D VGND VGND VPWR VPWR _34602_/Q sky130_fd_sc_hd__dfxtp_1
X_35582_ _35710_/CLK _35582_/D VGND VGND VPWR VPWR _35582_/Q sky130_fd_sc_hd__dfxtp_1
X_16748_ _32993_/Q _32929_/Q _32865_/Q _32801_/Q _16636_/X _16637_/X VGND VGND VPWR
+ VPWR _16748_/X sky130_fd_sc_hd__mux4_1
X_32794_ _33244_/CLK _32794_/D VGND VGND VPWR VPWR _32794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34533_ _35942_/CLK _34533_/D VGND VGND VPWR VPWR _34533_/Q sky130_fd_sc_hd__dfxtp_1
X_31745_ _36076_/Q input24/X _31763_/S VGND VGND VPWR VPWR _31746_/A sky130_fd_sc_hd__mux2_1
X_19467_ _19142_/X _19465_/X _19466_/X _19147_/X VGND VGND VPWR VPWR _19467_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16679_ _35807_/Q _32183_/Q _35679_/Q _35615_/Q _16607_/X _16608_/X VGND VGND VPWR
+ VPWR _16679_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18418_ _18326_/X _18416_/X _18417_/X _18337_/X VGND VGND VPWR VPWR _18418_/X sky130_fd_sc_hd__a22o_1
X_34464_ _35743_/CLK _34464_/D VGND VGND VPWR VPWR _34464_/Q sky130_fd_sc_hd__dfxtp_1
X_31676_ _36044_/Q input59/X _31678_/S VGND VGND VPWR VPWR _31677_/A sky130_fd_sc_hd__mux2_1
X_19398_ _33259_/Q _36139_/Q _33131_/Q _33067_/Q _19358_/X _19359_/X VGND VGND VPWR
+ VPWR _19398_/X sky130_fd_sc_hd__mux4_1
XFILLER_146_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33415_ _33544_/CLK _33415_/D VGND VGND VPWR VPWR _33415_/Q sky130_fd_sc_hd__dfxtp_1
X_36203_ _36204_/CLK _36203_/D VGND VGND VPWR VPWR _36203_/Q sky130_fd_sc_hd__dfxtp_1
X_18349_ _20294_/A VGND VGND VPWR VPWR _18349_/X sky130_fd_sc_hd__buf_6
X_30627_ _35546_/Q _29089_/X _30641_/S VGND VGND VPWR VPWR _30628_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34395_ _34970_/CLK _34395_/D VGND VGND VPWR VPWR _34395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36134_ _36134_/CLK _36134_/D VGND VGND VPWR VPWR _36134_/Q sky130_fd_sc_hd__dfxtp_1
X_33346_ _34050_/CLK _33346_/D VGND VGND VPWR VPWR _33346_/Q sky130_fd_sc_hd__dfxtp_1
X_21360_ _21043_/X _21358_/X _21359_/X _21046_/X VGND VGND VPWR VPWR _21360_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30558_ _30558_/A VGND VGND VPWR VPWR _35513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20311_ _20307_/X _20310_/X _20134_/X VGND VGND VPWR VPWR _20333_/A sky130_fd_sc_hd__o21ba_2
X_36065_ _36065_/CLK _36065_/D VGND VGND VPWR VPWR _36065_/Q sky130_fd_sc_hd__dfxtp_1
X_33277_ _36157_/CLK _33277_/D VGND VGND VPWR VPWR _33277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21291_ _21048_/X _21289_/X _21290_/X _21053_/X VGND VGND VPWR VPWR _21291_/X sky130_fd_sc_hd__a22o_1
Xinput60 DW[63] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__buf_12
Xinput71 R2[0] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30489_ _30489_/A VGND VGND VPWR VPWR _35480_/D sky130_fd_sc_hd__clkbuf_1
Xinput82 R3[5] VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__buf_2
X_35016_ _35079_/CLK _35016_/D VGND VGND VPWR VPWR _35016_/Q sky130_fd_sc_hd__dfxtp_1
X_23030_ _23030_/A VGND VGND VPWR VPWR _32062_/D sky130_fd_sc_hd__clkbuf_1
X_32228_ _35848_/CLK _32228_/D VGND VGND VPWR VPWR _32228_/Q sky130_fd_sc_hd__dfxtp_1
X_20242_ _33539_/Q _33475_/Q _33411_/Q _33347_/Q _20129_/X _20130_/X VGND VGND VPWR
+ VPWR _20242_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20173_ _19848_/X _20171_/X _20172_/X _19853_/X VGND VGND VPWR VPWR _20173_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32159_ _34016_/CLK _32159_/D VGND VGND VPWR VPWR _32159_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24981_ _23065_/X _32970_/Q _24987_/S VGND VGND VPWR VPWR _24982_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26720_ _26720_/A VGND VGND VPWR VPWR _33757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35918_ _35919_/CLK _35918_/D VGND VGND VPWR VPWR _35918_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23932_ _23932_/A VGND VGND VPWR VPWR _32506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26651_ _26651_/A VGND VGND VPWR VPWR _33725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35849_ _35849_/CLK _35849_/D VGND VGND VPWR VPWR _35849_/Q sky130_fd_sc_hd__dfxtp_1
X_23863_ _23863_/A VGND VGND VPWR VPWR _32473_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25602_ _25602_/A _31140_/B VGND VGND VPWR VPWR _25735_/S sky130_fd_sc_hd__nor2_8
XANTENNA_706 _22532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29370_ _23327_/X _34951_/Q _29374_/S VGND VGND VPWR VPWR _29371_/A sky130_fd_sc_hd__mux2_1
X_22814_ _22814_/A VGND VGND VPWR VPWR _36235_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_717 _22453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_728 _20870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26582_ _26582_/A VGND VGND VPWR VPWR _33692_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23794_ _23794_/A VGND VGND VPWR VPWR _32441_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_739 _21577_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28321_ _34485_/Q _24366_/X _28321_/S VGND VGND VPWR VPWR _28322_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25533_ _33198_/Q _24345_/X _25547_/S VGND VGND VPWR VPWR _25534_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22745_ _22741_/X _22744_/X _22453_/X VGND VGND VPWR VPWR _22753_/C sky130_fd_sc_hd__o21ba_1
XFILLER_129_1254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28252_ _34452_/Q _24264_/X _28258_/S VGND VGND VPWR VPWR _28253_/A sky130_fd_sc_hd__mux2_1
X_22676_ _33031_/Q _32967_/Q _32903_/Q _32839_/Q _20580_/X _20583_/X VGND VGND VPWR
+ VPWR _22676_/X sky130_fd_sc_hd__mux4_1
X_25464_ _31275_/B _30600_/B VGND VGND VPWR VPWR _25597_/S sky130_fd_sc_hd__nor2_8
XFILLER_129_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27203_ _27203_/A VGND VGND VPWR VPWR _33955_/D sky130_fd_sc_hd__clkbuf_1
X_24415_ _24415_/A VGND VGND VPWR VPWR _32708_/D sky130_fd_sc_hd__clkbuf_1
X_21627_ _21302_/X _21625_/X _21626_/X _21308_/X VGND VGND VPWR VPWR _21627_/X sky130_fd_sc_hd__a22o_1
X_28183_ _28183_/A VGND VGND VPWR VPWR _34419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25395_ _25395_/A VGND VGND VPWR VPWR _33134_/D sky130_fd_sc_hd__clkbuf_1
X_27134_ _26987_/X _33923_/Q _27146_/S VGND VGND VPWR VPWR _27135_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24346_ _32686_/Q _24345_/X _24367_/S VGND VGND VPWR VPWR _24347_/A sky130_fd_sc_hd__mux2_1
X_21558_ _21310_/X _21556_/X _21557_/X _21314_/X VGND VGND VPWR VPWR _21558_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20509_ _34571_/Q _32459_/Q _34443_/Q _34379_/Q _20231_/X _20232_/X VGND VGND VPWR
+ VPWR _20509_/X sky130_fd_sc_hd__mux4_1
X_24277_ _24441_/S VGND VGND VPWR VPWR _24305_/S sky130_fd_sc_hd__buf_6
X_27065_ _26884_/X _33890_/Q _27083_/S VGND VGND VPWR VPWR _27066_/A sky130_fd_sc_hd__mux2_1
X_21489_ _21302_/X _21487_/X _21488_/X _21308_/X VGND VGND VPWR VPWR _21489_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26016_ _26016_/A VGND VGND VPWR VPWR _33424_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23228_ input20/X VGND VGND VPWR VPWR _23228_/X sky130_fd_sc_hd__buf_4
XFILLER_84_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23159_ _31140_/A _29924_/A VGND VGND VPWR VPWR _23346_/S sky130_fd_sc_hd__nor2_8
XTAP_7055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1105 _17400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1116 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1127 input8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1138 _20206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15981_ input66/X VGND VGND VPWR VPWR _16059_/A sky130_fd_sc_hd__buf_8
XTAP_6365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27967_ _27967_/A VGND VGND VPWR VPWR _34317_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_1149 _19428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_212_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17720_ _17720_/A _17720_/B _17720_/C _17720_/D VGND VGND VPWR VPWR _17721_/A sky130_fd_sc_hd__or4_2
X_29706_ _35110_/Q _29126_/X _29716_/S VGND VGND VPWR VPWR _29707_/A sky130_fd_sc_hd__mux2_1
XTAP_6398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26918_ _26918_/A VGND VGND VPWR VPWR _33836_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27898_ _34284_/Q _24338_/X _27916_/S VGND VGND VPWR VPWR _27899_/A sky130_fd_sc_hd__mux2_1
XTAP_4941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29637_ _29637_/A VGND VGND VPWR VPWR _35077_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ _17651_/A VGND VGND VPWR VPWR _31994_/D sky130_fd_sc_hd__clkbuf_4
XTAP_4963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26849_ _26849_/A VGND VGND VPWR VPWR _33814_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16602_ _16349_/X _16600_/X _16601_/X _16355_/X VGND VGND VPWR VPWR _16602_/X sky130_fd_sc_hd__a22o_1
X_17582_ _17507_/X _17580_/X _17581_/X _17512_/X VGND VGND VPWR VPWR _17582_/X sky130_fd_sc_hd__a22o_1
X_29568_ _29568_/A VGND VGND VPWR VPWR _35044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19321_ _20147_/A VGND VGND VPWR VPWR _19321_/X sky130_fd_sc_hd__buf_6
X_28519_ _28519_/A VGND VGND VPWR VPWR _34578_/D sky130_fd_sc_hd__clkbuf_1
X_16533_ _16529_/X _16532_/X _16422_/X VGND VGND VPWR VPWR _16557_/A sky130_fd_sc_hd__o21ba_1
XFILLER_232_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29499_ _23316_/X _35012_/Q _29509_/S VGND VGND VPWR VPWR _29500_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31530_ _31530_/A VGND VGND VPWR VPWR _35974_/D sky130_fd_sc_hd__clkbuf_1
X_19252_ _19248_/X _19251_/X _19075_/X VGND VGND VPWR VPWR _19276_/A sky130_fd_sc_hd__o21ba_1
X_16464_ _16143_/X _16462_/X _16463_/X _16146_/X VGND VGND VPWR VPWR _16464_/X sky130_fd_sc_hd__a22o_1
XFILLER_92_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18203_ _33227_/Q _32587_/Q _35979_/Q _35915_/Q _16075_/X _16076_/X VGND VGND VPWR
+ VPWR _18203_/X sky130_fd_sc_hd__mux4_1
XPHY_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19183_ _33509_/Q _33445_/Q _33381_/Q _33317_/Q _19070_/X _19071_/X VGND VGND VPWR
+ VPWR _19183_/X sky130_fd_sc_hd__mux4_1
X_31461_ _31461_/A VGND VGND VPWR VPWR _35941_/D sky130_fd_sc_hd__clkbuf_1
XPHY_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16395_ _32983_/Q _32919_/Q _32855_/Q _32791_/Q _16283_/X _16284_/X VGND VGND VPWR
+ VPWR _16395_/X sky130_fd_sc_hd__mux4_1
XPHY_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33200_ _36013_/CLK _33200_/D VGND VGND VPWR VPWR _33200_/Q sky130_fd_sc_hd__dfxtp_1
X_18134_ _17149_/A _18132_/X _18133_/X _17152_/A VGND VGND VPWR VPWR _18134_/X sky130_fd_sc_hd__a22o_1
X_30412_ _30412_/A VGND VGND VPWR VPWR _35444_/D sky130_fd_sc_hd__clkbuf_1
X_34180_ _34310_/CLK _34180_/D VGND VGND VPWR VPWR _34180_/Q sky130_fd_sc_hd__dfxtp_1
X_31392_ _35909_/Q input51/X _31400_/S VGND VGND VPWR VPWR _31393_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33131_ _36139_/CLK _33131_/D VGND VGND VPWR VPWR _33131_/Q sky130_fd_sc_hd__dfxtp_1
X_18065_ _33799_/Q _33735_/Q _33671_/Q _33607_/Q _17902_/X _17903_/X VGND VGND VPWR
+ VPWR _18065_/X sky130_fd_sc_hd__mux4_1
X_30343_ _30343_/A VGND VGND VPWR VPWR _35411_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17016_ _33769_/Q _33705_/Q _33641_/Q _33577_/Q _16843_/X _16844_/X VGND VGND VPWR
+ VPWR _17016_/X sky130_fd_sc_hd__mux4_1
X_33062_ _36135_/CLK _33062_/D VGND VGND VPWR VPWR _33062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30274_ _30274_/A VGND VGND VPWR VPWR _35379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32013_ _36185_/CLK _32013_/D VGND VGND VPWR VPWR _32013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18967_ _20146_/A VGND VGND VPWR VPWR _18967_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_224_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17918_ _33026_/Q _32962_/Q _32898_/Q _32834_/Q _17695_/X _17696_/X VGND VGND VPWR
+ VPWR _17918_/X sky130_fd_sc_hd__mux4_1
XFILLER_230_1246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33964_ _35574_/CLK _33964_/D VGND VGND VPWR VPWR _33964_/Q sky130_fd_sc_hd__dfxtp_1
X_18898_ _18796_/X _18896_/X _18897_/X _18799_/X VGND VGND VPWR VPWR _18898_/X sky130_fd_sc_hd__a22o_1
XFILLER_152_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35703_ _35831_/CLK _35703_/D VGND VGND VPWR VPWR _35703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17849_ _17700_/X _17845_/X _17848_/X _17703_/X VGND VGND VPWR VPWR _17849_/X sky130_fd_sc_hd__a22o_1
X_32915_ _35986_/CLK _32915_/D VGND VGND VPWR VPWR _32915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33895_ _34087_/CLK _33895_/D VGND VGND VPWR VPWR _33895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20860_ _33171_/Q _32531_/Q _35923_/Q _35859_/Q _20663_/X _20665_/X VGND VGND VPWR
+ VPWR _20860_/X sky130_fd_sc_hd__mux4_1
X_32846_ _35982_/CLK _32846_/D VGND VGND VPWR VPWR _32846_/Q sky130_fd_sc_hd__dfxtp_1
X_35634_ _35826_/CLK _35634_/D VGND VGND VPWR VPWR _35634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19519_ _33198_/Q _32558_/Q _35950_/Q _35886_/Q _19374_/X _19375_/X VGND VGND VPWR
+ VPWR _19519_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32777_ _36105_/CLK _32777_/D VGND VGND VPWR VPWR _32777_/Q sky130_fd_sc_hd__dfxtp_1
X_20791_ _22446_/A VGND VGND VPWR VPWR _20791_/X sky130_fd_sc_hd__buf_6
X_35565_ _35949_/CLK _35565_/D VGND VGND VPWR VPWR _35565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_250_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _34053_/CLK sky130_fd_sc_hd__clkbuf_16
X_22530_ _22455_/X _22528_/X _22529_/X _22458_/X VGND VGND VPWR VPWR _22530_/X sky130_fd_sc_hd__a22o_1
X_34516_ _34706_/CLK _34516_/D VGND VGND VPWR VPWR _34516_/Q sky130_fd_sc_hd__dfxtp_1
X_31728_ _36068_/Q input15/X _31742_/S VGND VGND VPWR VPWR _31729_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35496_ _35819_/CLK _35496_/D VGND VGND VPWR VPWR _35496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22461_ _34560_/Q _32448_/Q _34432_/Q _34368_/Q _22178_/X _22179_/X VGND VGND VPWR
+ VPWR _22461_/X sky130_fd_sc_hd__mux4_1
XFILLER_206_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34447_ _35279_/CLK _34447_/D VGND VGND VPWR VPWR _34447_/Q sky130_fd_sc_hd__dfxtp_1
X_31659_ _31659_/A VGND VGND VPWR VPWR _36035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24200_ _24200_/A VGND VGND VPWR VPWR _32632_/D sky130_fd_sc_hd__clkbuf_1
X_21412_ _33763_/Q _33699_/Q _33635_/Q _33571_/Q _21090_/X _21091_/X VGND VGND VPWR
+ VPWR _21412_/X sky130_fd_sc_hd__mux4_1
X_25180_ input58/X VGND VGND VPWR VPWR _25180_/X sky130_fd_sc_hd__buf_2
X_34378_ _35339_/CLK _34378_/D VGND VGND VPWR VPWR _34378_/Q sky130_fd_sc_hd__dfxtp_1
X_22392_ _22392_/A _22392_/B _22392_/C _22392_/D VGND VGND VPWR VPWR _22393_/A sky130_fd_sc_hd__or4_4
XFILLER_120_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24131_ _24242_/S VGND VGND VPWR VPWR _24150_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_11_1310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36117_ _36117_/CLK _36117_/D VGND VGND VPWR VPWR _36117_/Q sky130_fd_sc_hd__dfxtp_1
X_33329_ _34033_/CLK _33329_/D VGND VGND VPWR VPWR _33329_/Q sky130_fd_sc_hd__dfxtp_1
X_21343_ _21339_/X _21342_/X _21022_/X VGND VGND VPWR VPWR _21365_/A sky130_fd_sc_hd__o21ba_1
XFILLER_175_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24062_ _24062_/A VGND VGND VPWR VPWR _32567_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36048_ _36048_/CLK _36048_/D VGND VGND VPWR VPWR _36048_/Q sky130_fd_sc_hd__dfxtp_1
X_21274_ _20949_/X _21272_/X _21273_/X _20955_/X VGND VGND VPWR VPWR _21274_/X sky130_fd_sc_hd__a22o_1
XFILLER_239_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23013_ input38/X VGND VGND VPWR VPWR _23013_/X sky130_fd_sc_hd__clkbuf_4
X_20225_ _33218_/Q _32578_/Q _35970_/Q _35906_/Q _20080_/X _20081_/X VGND VGND VPWR
+ VPWR _20225_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28870_ _26956_/X _34745_/Q _28882_/S VGND VGND VPWR VPWR _28871_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27821_ _34248_/Q _24425_/X _27823_/S VGND VGND VPWR VPWR _27822_/A sky130_fd_sc_hd__mux2_1
X_20156_ _34816_/Q _34752_/Q _34688_/Q _34624_/Q _19941_/X _19942_/X VGND VGND VPWR
+ VPWR _20156_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27752_ _34215_/Q _24323_/X _27760_/S VGND VGND VPWR VPWR _27753_/A sky130_fd_sc_hd__mux2_1
X_24964_ _24964_/A VGND VGND VPWR VPWR _32961_/D sky130_fd_sc_hd__clkbuf_1
X_20087_ _19802_/X _20085_/X _20086_/X _19805_/X VGND VGND VPWR VPWR _20087_/X sky130_fd_sc_hd__a22o_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26703_ _26703_/A VGND VGND VPWR VPWR _33749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23915_ _23915_/A VGND VGND VPWR VPWR _32498_/D sky130_fd_sc_hd__clkbuf_1
X_27683_ _27683_/A VGND VGND VPWR VPWR _34182_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24895_ _22938_/X _32929_/Q _24895_/S VGND VGND VPWR VPWR _24896_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29422_ _29422_/A VGND VGND VPWR VPWR _34975_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26634_ _26634_/A VGND VGND VPWR VPWR _33717_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_503 _17793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_514 _17938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23846_ _23846_/A VGND VGND VPWR VPWR _32465_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_525 _18004_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_536 _20096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29353_ _23300_/X _34943_/Q _29353_/S VGND VGND VPWR VPWR _29354_/A sky130_fd_sc_hd__mux2_1
XANTENNA_547 _20162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26565_ _26565_/A VGND VGND VPWR VPWR _33684_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_558 _20295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20989_ _20743_/X _20987_/X _20988_/X _20746_/X VGND VGND VPWR VPWR _20989_/X sky130_fd_sc_hd__a22o_1
XFILLER_129_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23777_ _23777_/A VGND VGND VPWR VPWR _32433_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_569 _20147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_241_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _34817_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28304_ _28304_/A VGND VGND VPWR VPWR _34476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_918 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25516_ _33190_/Q _24320_/X _25526_/S VGND VGND VPWR VPWR _25517_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22728_ _33545_/Q _33481_/Q _33417_/Q _33353_/Q _22429_/X _22430_/X VGND VGND VPWR
+ VPWR _22728_/X sky130_fd_sc_hd__mux4_1
X_29284_ _23136_/X _34910_/Q _29290_/S VGND VGND VPWR VPWR _29285_/A sky130_fd_sc_hd__mux2_1
X_26496_ _26496_/A VGND VGND VPWR VPWR _33652_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28235_ _28235_/A VGND VGND VPWR VPWR _34444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25447_ _25447_/A VGND VGND VPWR VPWR _33159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22659_ _34566_/Q _32454_/Q _34438_/Q _34374_/Q _22531_/X _22532_/X VGND VGND VPWR
+ VPWR _22659_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16180_ _16176_/X _16179_/X _16011_/X VGND VGND VPWR VPWR _16204_/A sky130_fd_sc_hd__o21ba_1
XFILLER_173_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28166_ _28166_/A VGND VGND VPWR VPWR _34411_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25378_ _25378_/A VGND VGND VPWR VPWR _33126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27117_ _26962_/X _33915_/Q _27125_/S VGND VGND VPWR VPWR _27118_/A sky130_fd_sc_hd__mux2_1
X_24329_ input20/X VGND VGND VPWR VPWR _24329_/X sky130_fd_sc_hd__buf_4
X_28097_ _27011_/X _34379_/Q _28101_/S VGND VGND VPWR VPWR _28098_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27048_ _26860_/X _33882_/Q _27062_/S VGND VGND VPWR VPWR _27049_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19870_ _19647_/X _19868_/X _19869_/X _19650_/X VGND VGND VPWR VPWR _19870_/X sky130_fd_sc_hd__a22o_1
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18821_ _34522_/Q _32410_/Q _34394_/Q _34330_/Q _18819_/X _18820_/X VGND VGND VPWR
+ VPWR _18821_/X sky130_fd_sc_hd__mux4_1
XTAP_6140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28999_ _34806_/Q _24369_/X _29017_/S VGND VGND VPWR VPWR _29000_/A sky130_fd_sc_hd__mux2_1
XTAP_6162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18752_ _35032_/Q _34968_/Q _34904_/Q _34840_/Q _18750_/X _18751_/X VGND VGND VPWR
+ VPWR _18752_/X sky130_fd_sc_hd__mux4_1
XTAP_5450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17703_ _17858_/A VGND VGND VPWR VPWR _17703_/X sky130_fd_sc_hd__buf_4
XFILLER_248_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18683_ _20256_/A VGND VGND VPWR VPWR _18683_/X sky130_fd_sc_hd__buf_6
X_30961_ _30961_/A VGND VGND VPWR VPWR _35704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32700_ _36156_/CLK _32700_/D VGND VGND VPWR VPWR _32700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_480_CLK clkbuf_6_3__f_CLK/X VGND VGND VPWR VPWR _35864_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17634_ _35834_/Q _32212_/Q _35706_/Q _35642_/Q _17313_/X _17314_/X VGND VGND VPWR
+ VPWR _17634_/X sky130_fd_sc_hd__mux4_1
X_33680_ _34194_/CLK _33680_/D VGND VGND VPWR VPWR _33680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30892_ _31003_/S VGND VGND VPWR VPWR _30911_/S sky130_fd_sc_hd__buf_4
XFILLER_63_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32631_ _36087_/CLK _32631_/D VGND VGND VPWR VPWR _32631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17565_ _33016_/Q _32952_/Q _32888_/Q _32824_/Q _17342_/X _17343_/X VGND VGND VPWR
+ VPWR _17565_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_232_CLK clkbuf_6_60__f_CLK/X VGND VGND VPWR VPWR _36103_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_205_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19304_ _19298_/X _19303_/X _19094_/X VGND VGND VPWR VPWR _19314_/C sky130_fd_sc_hd__o21ba_1
XFILLER_72_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35350_ _35927_/CLK _35350_/D VGND VGND VPWR VPWR _35350_/Q sky130_fd_sc_hd__dfxtp_1
X_16516_ _34778_/Q _34714_/Q _34650_/Q _34586_/Q _16229_/X _16230_/X VGND VGND VPWR
+ VPWR _16516_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32562_ _36141_/CLK _32562_/D VGND VGND VPWR VPWR _32562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17496_ _17347_/X _17492_/X _17495_/X _17350_/X VGND VGND VPWR VPWR _17496_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31513_ _31513_/A VGND VGND VPWR VPWR _35966_/D sky130_fd_sc_hd__clkbuf_1
X_34301_ _36157_/CLK _34301_/D VGND VGND VPWR VPWR _34301_/Q sky130_fd_sc_hd__dfxtp_1
X_19235_ _20294_/A VGND VGND VPWR VPWR _19235_/X sky130_fd_sc_hd__buf_6
X_35281_ _35281_/CLK _35281_/D VGND VGND VPWR VPWR _35281_/Q sky130_fd_sc_hd__dfxtp_1
X_16447_ _16443_/X _16444_/X _16445_/X _16446_/X VGND VGND VPWR VPWR _16447_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32493_ _36013_/CLK _32493_/D VGND VGND VPWR VPWR _32493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34232_ _34296_/CLK _34232_/D VGND VGND VPWR VPWR _34232_/Q sky130_fd_sc_hd__dfxtp_1
X_19166_ _33188_/Q _32548_/Q _35940_/Q _35876_/Q _19021_/X _19022_/X VGND VGND VPWR
+ VPWR _19166_/X sky130_fd_sc_hd__mux4_1
X_31444_ _31444_/A VGND VGND VPWR VPWR _35933_/D sky130_fd_sc_hd__clkbuf_1
X_16378_ _16087_/X _16376_/X _16377_/X _16097_/X VGND VGND VPWR VPWR _16378_/X sky130_fd_sc_hd__a22o_1
XFILLER_223_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18117_ _35336_/Q _35272_/Q _35208_/Q _32328_/Q _16088_/X _16090_/X VGND VGND VPWR
+ VPWR _18117_/X sky130_fd_sc_hd__mux4_1
X_34163_ _34291_/CLK _34163_/D VGND VGND VPWR VPWR _34163_/Q sky130_fd_sc_hd__dfxtp_1
X_31375_ _35901_/Q input42/X _31379_/S VGND VGND VPWR VPWR _31376_/A sky130_fd_sc_hd__mux2_1
X_19097_ _34786_/Q _34722_/Q _34658_/Q _34594_/Q _18882_/X _18883_/X VGND VGND VPWR
+ VPWR _19097_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33114_ _36124_/CLK _33114_/D VGND VGND VPWR VPWR _33114_/Q sky130_fd_sc_hd__dfxtp_1
X_30326_ _30326_/A VGND VGND VPWR VPWR _35404_/D sky130_fd_sc_hd__clkbuf_1
X_18048_ _18044_/X _18047_/X _17842_/X _17843_/X VGND VGND VPWR VPWR _18063_/B sky130_fd_sc_hd__o211a_1
XFILLER_133_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34094_ _34222_/CLK _34094_/D VGND VGND VPWR VPWR _34094_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_299_CLK clkbuf_6_50__f_CLK/X VGND VGND VPWR VPWR _35965_/CLK sky130_fd_sc_hd__clkbuf_16
X_33045_ _36117_/CLK _33045_/D VGND VGND VPWR VPWR _33045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30257_ _30257_/A VGND VGND VPWR VPWR _35371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20010_ _20004_/X _20009_/X _19800_/X VGND VGND VPWR VPWR _20020_/C sky130_fd_sc_hd__o21ba_1
XFILLER_113_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30188_ _35339_/Q _29240_/X _30192_/S VGND VGND VPWR VPWR _30189_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19999_ _19993_/X _19998_/X _19789_/X _19790_/X VGND VGND VPWR VPWR _20020_/B sky130_fd_sc_hd__o211a_1
XFILLER_87_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34996_ _35061_/CLK _34996_/D VGND VGND VPWR VPWR _34996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33947_ _36194_/CLK _33947_/D VGND VGND VPWR VPWR _33947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21961_ _35314_/Q _35250_/Q _35186_/Q _32306_/Q _21959_/X _21960_/X VGND VGND VPWR
+ VPWR _21961_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_999 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23700_ _26549_/C _25462_/A VGND VGND VPWR VPWR _30465_/B sky130_fd_sc_hd__nor2_8
Xclkbuf_leaf_471_CLK clkbuf_6_8__f_CLK/X VGND VGND VPWR VPWR _35555_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20912_ _20736_/X _20910_/X _20911_/X _20741_/X VGND VGND VPWR VPWR _20912_/X sky130_fd_sc_hd__a22o_1
X_24680_ _23022_/X _32828_/Q _24686_/S VGND VGND VPWR VPWR _24681_/A sky130_fd_sc_hd__mux2_1
X_21892_ _21749_/X _21890_/X _21891_/X _21752_/X VGND VGND VPWR VPWR _21892_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33878_ _34006_/CLK _33878_/D VGND VGND VPWR VPWR _33878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ _33491_/Q _33427_/Q _33363_/Q _33299_/Q _20598_/X _20599_/X VGND VGND VPWR
+ VPWR _20843_/X sky130_fd_sc_hd__mux4_1
X_23631_ _23631_/A VGND VGND VPWR VPWR _32365_/D sky130_fd_sc_hd__clkbuf_1
X_35617_ _35807_/CLK _35617_/D VGND VGND VPWR VPWR _35617_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32829_ _32959_/CLK _32829_/D VGND VGND VPWR VPWR _32829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_223_CLK clkbuf_6_55__f_CLK/X VGND VGND VPWR VPWR _35075_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26350_ _25094_/X _33583_/Q _26362_/S VGND VGND VPWR VPWR _26351_/A sky130_fd_sc_hd__mux2_1
X_20774_ _33745_/Q _33681_/Q _33617_/Q _33553_/Q _20737_/X _20738_/X VGND VGND VPWR
+ VPWR _20774_/X sky130_fd_sc_hd__mux4_1
X_23562_ input84/X input85/X VGND VGND VPWR VPWR _25462_/A sky130_fd_sc_hd__nand2b_4
X_35548_ _35933_/CLK _35548_/D VGND VGND VPWR VPWR _35548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25301_ _25301_/A VGND VGND VPWR VPWR _33090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22513_ _22507_/X _22512_/X _22434_/X VGND VGND VPWR VPWR _22537_/A sky130_fd_sc_hd__o21ba_1
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26281_ _24989_/X _33550_/Q _26299_/S VGND VGND VPWR VPWR _26282_/A sky130_fd_sc_hd__mux2_1
X_23493_ _22976_/X _32301_/Q _23509_/S VGND VGND VPWR VPWR _23494_/A sky130_fd_sc_hd__mux2_1
X_35479_ _35863_/CLK _35479_/D VGND VGND VPWR VPWR _35479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28020_ _26897_/X _34342_/Q _28030_/S VGND VGND VPWR VPWR _28021_/A sky130_fd_sc_hd__mux2_1
X_22444_ _22438_/X _22441_/X _22442_/X _22443_/X VGND VGND VPWR VPWR _22469_/B sky130_fd_sc_hd__o211a_1
X_25232_ _25322_/S VGND VGND VPWR VPWR _25251_/S sky130_fd_sc_hd__buf_4
XFILLER_183_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25163_ _25162_/X _33029_/Q _25175_/S VGND VGND VPWR VPWR _25164_/A sky130_fd_sc_hd__mux2_1
X_22375_ _22368_/X _22374_/X _22089_/X _22090_/X VGND VGND VPWR VPWR _22392_/B sky130_fd_sc_hd__o211a_1
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1022 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24114_ _24114_/A VGND VGND VPWR VPWR _32591_/D sky130_fd_sc_hd__clkbuf_1
X_21326_ _34784_/Q _34720_/Q _34656_/Q _34592_/Q _21182_/X _21183_/X VGND VGND VPWR
+ VPWR _21326_/X sky130_fd_sc_hd__mux4_1
X_25094_ input27/X VGND VGND VPWR VPWR _25094_/X sky130_fd_sc_hd__buf_2
X_29971_ _29971_/A VGND VGND VPWR VPWR _35235_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28922_ _28922_/A VGND VGND VPWR VPWR _34769_/D sky130_fd_sc_hd__clkbuf_1
X_21257_ _34526_/Q _32414_/Q _34398_/Q _34334_/Q _21119_/X _21120_/X VGND VGND VPWR
+ VPWR _21257_/X sky130_fd_sc_hd__mux4_1
X_24045_ _24045_/A VGND VGND VPWR VPWR _32559_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20208_ _20208_/A VGND VGND VPWR VPWR _20208_/X sky130_fd_sc_hd__clkbuf_8
X_28853_ _26931_/X _34737_/Q _28861_/S VGND VGND VPWR VPWR _28854_/A sky130_fd_sc_hd__mux2_1
X_21188_ _35036_/Q _34972_/Q _34908_/Q _34844_/Q _21050_/X _21051_/X VGND VGND VPWR
+ VPWR _21188_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27804_ _27831_/S VGND VGND VPWR VPWR _27823_/S sky130_fd_sc_hd__clkbuf_8
X_20139_ _32512_/Q _32384_/Q _32064_/Q _36032_/Q _19929_/X _20070_/X VGND VGND VPWR
+ VPWR _20139_/X sky130_fd_sc_hd__mux4_1
X_28784_ _26829_/X _34704_/Q _28798_/S VGND VGND VPWR VPWR _28785_/A sky130_fd_sc_hd__mux2_1
XTAP_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25996_ _25996_/A VGND VGND VPWR VPWR _33415_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27735_ _34207_/Q _24298_/X _27739_/S VGND VGND VPWR VPWR _27736_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24947_ _24947_/A VGND VGND VPWR VPWR _32953_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_462_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _34859_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27666_ _27666_/A VGND VGND VPWR VPWR _34174_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1004 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24878_ _24878_/A VGND VGND VPWR VPWR _32920_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_300 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_311 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29405_ _29405_/A VGND VGND VPWR VPWR _34967_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_322 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_333 _32141_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26617_ _25088_/X _33709_/Q _26633_/S VGND VGND VPWR VPWR _26618_/A sky130_fd_sc_hd__mux2_1
XTAP_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23829_ _23829_/A VGND VGND VPWR VPWR _32458_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_344 _36205_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27597_ _27597_/A VGND VGND VPWR VPWR _34141_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_355 _36206_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_214_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _35078_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_366 _36207_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_377 _36208_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29336_ _29336_/A VGND VGND VPWR VPWR _34934_/D sky130_fd_sc_hd__clkbuf_1
X_17350_ _17858_/A VGND VGND VPWR VPWR _17350_/X sky130_fd_sc_hd__buf_4
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_388 _36209_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26548_ _26548_/A VGND VGND VPWR VPWR _33677_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_399 _36210_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16301_ _17007_/A VGND VGND VPWR VPWR _16301_/X sky130_fd_sc_hd__buf_4
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29267_ _23111_/X _34902_/Q _29269_/S VGND VGND VPWR VPWR _29268_/A sky130_fd_sc_hd__mux2_1
X_17281_ _35824_/Q _32201_/Q _35696_/Q _35632_/Q _16960_/X _16961_/X VGND VGND VPWR
+ VPWR _17281_/X sky130_fd_sc_hd__mux4_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26479_ _25084_/X _33644_/Q _26497_/S VGND VGND VPWR VPWR _26480_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19020_ _35552_/Q _35488_/Q _35424_/Q _35360_/Q _18844_/X _18845_/X VGND VGND VPWR
+ VPWR _19020_/X sky130_fd_sc_hd__mux4_1
X_28218_ _26990_/X _34436_/Q _28228_/S VGND VGND VPWR VPWR _28219_/A sky130_fd_sc_hd__mux2_1
X_16232_ _35282_/Q _35218_/Q _35154_/Q _32274_/Q _16079_/X _16081_/X VGND VGND VPWR
+ VPWR _16232_/X sky130_fd_sc_hd__mux4_1
XFILLER_146_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29198_ _34877_/Q _29197_/X _29204_/S VGND VGND VPWR VPWR _29199_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16163_ _34768_/Q _34704_/Q _34640_/Q _34576_/Q _16075_/X _16076_/X VGND VGND VPWR
+ VPWR _16163_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28149_ _26888_/X _34403_/Q _28165_/S VGND VGND VPWR VPWR _28150_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31160_ _35799_/Q input64/X _31160_/S VGND VGND VPWR VPWR _31161_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16094_ _17157_/A VGND VGND VPWR VPWR _16094_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_181_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30111_ _35302_/Q _29126_/X _30121_/S VGND VGND VPWR VPWR _30112_/A sky130_fd_sc_hd__mux2_1
X_19922_ _34042_/Q _33978_/Q _33914_/Q _32250_/Q _19673_/X _19674_/X VGND VGND VPWR
+ VPWR _19922_/X sky130_fd_sc_hd__mux4_1
XFILLER_170_968 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31091_ _35766_/Q _29175_/X _31109_/S VGND VGND VPWR VPWR _31092_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30042_ _30042_/A VGND VGND VPWR VPWR _35269_/D sky130_fd_sc_hd__clkbuf_1
X_19853_ _20206_/A VGND VGND VPWR VPWR _19853_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18804_ _18649_/X _18802_/X _18803_/X _18655_/X VGND VGND VPWR VPWR _18804_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34850_ _35299_/CLK _34850_/D VGND VGND VPWR VPWR _34850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16996_ _35752_/Q _35112_/Q _34472_/Q _33832_/Q _16787_/X _16788_/X VGND VGND VPWR
+ VPWR _16996_/X sky130_fd_sc_hd__mux4_1
X_19784_ _33270_/Q _36150_/Q _33142_/Q _33078_/Q _19711_/X _19712_/X VGND VGND VPWR
+ VPWR _19784_/X sky130_fd_sc_hd__mux4_1
XFILLER_205_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33801_ _34817_/CLK _33801_/D VGND VGND VPWR VPWR _33801_/Q sky130_fd_sc_hd__dfxtp_1
X_18735_ _20295_/A VGND VGND VPWR VPWR _18735_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34781_ _34781_/CLK _34781_/D VGND VGND VPWR VPWR _34781_/Q sky130_fd_sc_hd__dfxtp_1
X_31993_ _36200_/CLK _31993_/D VGND VGND VPWR VPWR _31993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_453_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _35239_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33732_ _33795_/CLK _33732_/D VGND VGND VPWR VPWR _33732_/Q sky130_fd_sc_hd__dfxtp_1
X_18666_ _18588_/X _18664_/X _18665_/X _18591_/X VGND VGND VPWR VPWR _18666_/X sky130_fd_sc_hd__a22o_1
X_30944_ _30944_/A VGND VGND VPWR VPWR _35696_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17617_ _17617_/A VGND VGND VPWR VPWR _31993_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_224_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30875_ _30875_/A VGND VGND VPWR VPWR _35663_/D sky130_fd_sc_hd__clkbuf_1
X_33663_ _33793_/CLK _33663_/D VGND VGND VPWR VPWR _33663_/Q sky130_fd_sc_hd__dfxtp_1
X_18597_ _18593_/X _18594_/X _18595_/X _18596_/X VGND VGND VPWR VPWR _18597_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_205_CLK clkbuf_6_52__f_CLK/X VGND VGND VPWR VPWR _35909_/CLK sky130_fd_sc_hd__clkbuf_16
X_35402_ _35852_/CLK _35402_/D VGND VGND VPWR VPWR _35402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17548_ _17901_/A VGND VGND VPWR VPWR _17548_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_162_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32614_ _36070_/CLK _32614_/D VGND VGND VPWR VPWR _32614_/Q sky130_fd_sc_hd__dfxtp_1
X_33594_ _33787_/CLK _33594_/D VGND VGND VPWR VPWR _33594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35333_ _35333_/CLK _35333_/D VGND VGND VPWR VPWR _35333_/Q sky130_fd_sc_hd__dfxtp_1
X_32545_ _35938_/CLK _32545_/D VGND VGND VPWR VPWR _32545_/Q sky130_fd_sc_hd__dfxtp_1
X_17479_ _34038_/Q _33974_/Q _33910_/Q _32246_/Q _17373_/X _17374_/X VGND VGND VPWR
+ VPWR _17479_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19218_ _19214_/X _19217_/X _19075_/X VGND VGND VPWR VPWR _19244_/A sky130_fd_sc_hd__o21ba_1
X_35264_ _35328_/CLK _35264_/D VGND VGND VPWR VPWR _35264_/Q sky130_fd_sc_hd__dfxtp_1
X_20490_ _20208_/X _20488_/X _20489_/X _20211_/X VGND VGND VPWR VPWR _20490_/X sky130_fd_sc_hd__a22o_1
XFILLER_165_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32476_ _32860_/CLK _32476_/D VGND VGND VPWR VPWR _32476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31427_ _31427_/A VGND VGND VPWR VPWR _35925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_943 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34215_ _34279_/CLK _34215_/D VGND VGND VPWR VPWR _34215_/Q sky130_fd_sc_hd__dfxtp_1
X_19149_ _20208_/A VGND VGND VPWR VPWR _19149_/X sky130_fd_sc_hd__clkbuf_4
X_35195_ _35580_/CLK _35195_/D VGND VGND VPWR VPWR _35195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22160_ _22154_/X _22159_/X _22081_/X VGND VGND VPWR VPWR _22184_/A sky130_fd_sc_hd__o21ba_1
X_34146_ _34146_/CLK _34146_/D VGND VGND VPWR VPWR _34146_/Q sky130_fd_sc_hd__dfxtp_1
X_31358_ _35893_/Q input33/X _31358_/S VGND VGND VPWR VPWR _31359_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21111_ _20888_/X _21109_/X _21110_/X _20891_/X VGND VGND VPWR VPWR _21111_/X sky130_fd_sc_hd__a22o_1
X_30309_ _35396_/Q _29219_/X _30319_/S VGND VGND VPWR VPWR _30310_/A sky130_fd_sc_hd__mux2_1
X_22091_ _22085_/X _22088_/X _22089_/X _22090_/X VGND VGND VPWR VPWR _22116_/B sky130_fd_sc_hd__o211a_1
X_34077_ _36200_/CLK _34077_/D VGND VGND VPWR VPWR _34077_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31289_ _35860_/Q input61/X _31295_/S VGND VGND VPWR VPWR _31290_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33028_ _36039_/CLK _33028_/D VGND VGND VPWR VPWR _33028_/Q sky130_fd_sc_hd__dfxtp_1
X_21042_ _21037_/X _21040_/X _21041_/X VGND VGND VPWR VPWR _21057_/C sky130_fd_sc_hd__o21ba_1
XFILLER_141_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25850_ _25153_/X _33346_/Q _25864_/S VGND VGND VPWR VPWR _25851_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24801_ _24801_/A VGND VGND VPWR VPWR _32884_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25781_ _25781_/A VGND VGND VPWR VPWR _33313_/D sky130_fd_sc_hd__clkbuf_1
X_34979_ _35299_/CLK _34979_/D VGND VGND VPWR VPWR _34979_/Q sky130_fd_sc_hd__dfxtp_1
X_22993_ _22993_/A VGND VGND VPWR VPWR _32050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27520_ _26959_/X _34106_/Q _27530_/S VGND VGND VPWR VPWR _27521_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_444_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _36070_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_215_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24732_ _24732_/A VGND VGND VPWR VPWR _32851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21944_ _33010_/Q _32946_/Q _32882_/Q _32818_/Q _21942_/X _21943_/X VGND VGND VPWR
+ VPWR _21944_/X sky130_fd_sc_hd__mux4_1
XFILLER_227_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27451_ _26857_/X _34073_/Q _27467_/S VGND VGND VPWR VPWR _27452_/A sky130_fd_sc_hd__mux2_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24663_ _22997_/X _32820_/Q _24665_/S VGND VGND VPWR VPWR _24664_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_6_24__f_CLK clkbuf_5_12_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_73_CLK/A sky130_fd_sc_hd__clkbuf_16
X_21875_ _21655_/X _21873_/X _21874_/X _21661_/X VGND VGND VPWR VPWR _21875_/X sky130_fd_sc_hd__a22o_1
XFILLER_208_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26402_ _25171_/X _33608_/Q _26404_/S VGND VGND VPWR VPWR _26403_/A sky130_fd_sc_hd__mux2_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23614_ _23614_/A VGND VGND VPWR VPWR _32357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20826_ _33170_/Q _32530_/Q _35922_/Q _35858_/Q _20663_/X _20665_/X VGND VGND VPWR
+ VPWR _20826_/X sky130_fd_sc_hd__mux4_1
X_27382_ _27382_/A VGND VGND VPWR VPWR _34040_/D sky130_fd_sc_hd__clkbuf_1
X_24594_ _22895_/X _32787_/Q _24602_/S VGND VGND VPWR VPWR _24595_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29121_ _34852_/Q _29120_/X _29142_/S VGND VGND VPWR VPWR _29122_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26333_ _25069_/X _33575_/Q _26341_/S VGND VGND VPWR VPWR _26334_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23545_ _23053_/X _32326_/Q _23551_/S VGND VGND VPWR VPWR _23546_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20757_ _35728_/Q _35088_/Q _34448_/Q _33808_/Q _20649_/X _20651_/X VGND VGND VPWR
+ VPWR _20757_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29052_ _29247_/S VGND VGND VPWR VPWR _29080_/S sky130_fd_sc_hd__buf_4
XFILLER_52_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26264_ _26264_/A VGND VGND VPWR VPWR _33542_/D sky130_fd_sc_hd__clkbuf_1
X_20688_ _22312_/A VGND VGND VPWR VPWR _20688_/X sky130_fd_sc_hd__buf_6
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23476_ _22951_/X _32293_/Q _23488_/S VGND VGND VPWR VPWR _23477_/A sky130_fd_sc_hd__mux2_1
X_28003_ _26872_/X _34334_/Q _28009_/S VGND VGND VPWR VPWR _28004_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25215_ _25215_/A VGND VGND VPWR VPWR _33049_/D sky130_fd_sc_hd__clkbuf_1
X_22427_ _34304_/Q _34240_/Q _34176_/Q _34112_/Q _22395_/X _22396_/X VGND VGND VPWR
+ VPWR _22427_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26195_ _26195_/A VGND VGND VPWR VPWR _33509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25146_ input46/X VGND VGND VPWR VPWR _25146_/X sky130_fd_sc_hd__buf_2
X_22358_ _34046_/Q _33982_/Q _33918_/Q _32254_/Q _22326_/X _22327_/X VGND VGND VPWR
+ VPWR _22358_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21309_ _21302_/X _21304_/X _21307_/X _21308_/X VGND VGND VPWR VPWR _21309_/X sky130_fd_sc_hd__a22o_1
X_22289_ _22155_/X _22287_/X _22288_/X _22158_/X VGND VGND VPWR VPWR _22289_/X sky130_fd_sc_hd__a22o_1
XFILLER_3_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29954_ _29954_/A VGND VGND VPWR VPWR _35227_/D sky130_fd_sc_hd__clkbuf_1
X_25077_ _25077_/A VGND VGND VPWR VPWR _33001_/D sky130_fd_sc_hd__clkbuf_1
X_28905_ _27008_/X _34762_/Q _28911_/S VGND VGND VPWR VPWR _28906_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24028_ _24028_/A VGND VGND VPWR VPWR _32551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29885_ _35195_/Q _29191_/X _29893_/S VGND VGND VPWR VPWR _29886_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16850_ _33508_/Q _33444_/Q _33380_/Q _33316_/Q _16770_/X _16771_/X VGND VGND VPWR
+ VPWR _16850_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28836_ _26906_/X _34729_/Q _28840_/S VGND VGND VPWR VPWR _28837_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28767_ _28767_/A VGND VGND VPWR VPWR _34696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16781_ _32994_/Q _32930_/Q _32866_/Q _32802_/Q _16636_/X _16637_/X VGND VGND VPWR
+ VPWR _16781_/X sky130_fd_sc_hd__mux4_1
X_25979_ _25979_/A VGND VGND VPWR VPWR _33407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18520_ _18326_/X _18518_/X _18519_/X _18337_/X VGND VGND VPWR VPWR _18520_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_435_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _34279_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_219_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27718_ _34199_/Q _24273_/X _27718_/S VGND VGND VPWR VPWR _27719_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28698_ _28698_/A VGND VGND VPWR VPWR _34663_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_963 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18451_ _18314_/X _18449_/X _18450_/X _18323_/X VGND VGND VPWR VPWR _18451_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27649_ _34166_/Q _24369_/X _27667_/S VGND VGND VPWR VPWR _27650_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_130 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_152 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _34292_/Q _34228_/Q _34164_/Q _34100_/Q _17089_/X _17090_/X VGND VGND VPWR
+ VPWR _17402_/X sky130_fd_sc_hd__mux4_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _35278_/Q _35214_/Q _35150_/Q _32270_/Q _18379_/X _18381_/X VGND VGND VPWR
+ VPWR _18382_/X sky130_fd_sc_hd__mux4_1
XANTENNA_163 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30660_ _35562_/Q _29138_/X _30662_/S VGND VGND VPWR VPWR _30661_/A sky130_fd_sc_hd__mux2_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_185 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_196 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29319_ _29319_/A VGND VGND VPWR VPWR _34926_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _17195_/X _17331_/X _17332_/X _17200_/X VGND VGND VPWR VPWR _17333_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30591_ _30591_/A VGND VGND VPWR VPWR _35529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32330_ _35147_/CLK _32330_/D VGND VGND VPWR VPWR _32330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17264_ _17264_/A VGND VGND VPWR VPWR _31983_/D sky130_fd_sc_hd__clkbuf_1
X_19003_ _20062_/A VGND VGND VPWR VPWR _19003_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_179_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16215_ _33234_/Q _36114_/Q _33106_/Q _33042_/Q _16020_/X _16021_/X VGND VGND VPWR
+ VPWR _16215_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32261_ _34057_/CLK _32261_/D VGND VGND VPWR VPWR _32261_/Q sky130_fd_sc_hd__dfxtp_1
X_17195_ _17901_/A VGND VGND VPWR VPWR _17195_/X sky130_fd_sc_hd__buf_2
X_34000_ _34004_/CLK _34000_/D VGND VGND VPWR VPWR _34000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31212_ _31212_/A VGND VGND VPWR VPWR _35823_/D sky130_fd_sc_hd__clkbuf_1
X_16146_ _17865_/A VGND VGND VPWR VPWR _16146_/X sky130_fd_sc_hd__buf_4
XFILLER_143_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32192_ _35818_/CLK _32192_/D VGND VGND VPWR VPWR _32192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31143_ _31143_/A VGND VGND VPWR VPWR _35790_/D sky130_fd_sc_hd__clkbuf_1
X_16077_ _34766_/Q _34702_/Q _34638_/Q _34574_/Q _16075_/X _16076_/X VGND VGND VPWR
+ VPWR _16077_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19905_ _35577_/Q _35513_/Q _35449_/Q _35385_/Q _19903_/X _19904_/X VGND VGND VPWR
+ VPWR _19905_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31074_ _35758_/Q _29151_/X _31088_/S VGND VGND VPWR VPWR _31075_/A sky130_fd_sc_hd__mux2_1
X_35951_ _35951_/CLK _35951_/D VGND VGND VPWR VPWR _35951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34902_ _35028_/CLK _34902_/D VGND VGND VPWR VPWR _34902_/Q sky130_fd_sc_hd__dfxtp_1
X_30025_ _30025_/A VGND VGND VPWR VPWR _35261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19836_ _33207_/Q _32567_/Q _35959_/Q _35895_/Q _19727_/X _19728_/X VGND VGND VPWR
+ VPWR _19836_/X sky130_fd_sc_hd__mux4_1
X_35882_ _35946_/CLK _35882_/D VGND VGND VPWR VPWR _35882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34833_ _36211_/CLK _34833_/D VGND VGND VPWR VPWR _34833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19767_ _34549_/Q _32437_/Q _34421_/Q _34357_/Q _19525_/X _19526_/X VGND VGND VPWR
+ VPWR _19767_/X sky130_fd_sc_hd__mux4_1
Xinput3 DW[11] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__buf_8
X_16979_ _34280_/Q _34216_/Q _34152_/Q _34088_/Q _16736_/X _16737_/X VGND VGND VPWR
+ VPWR _16979_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_426_CLK clkbuf_6_36__f_CLK/X VGND VGND VPWR VPWR _36009_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18718_ _20096_/A VGND VGND VPWR VPWR _18718_/X sky130_fd_sc_hd__buf_4
XFILLER_37_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34764_ _35340_/CLK _34764_/D VGND VGND VPWR VPWR _34764_/Q sky130_fd_sc_hd__dfxtp_1
X_31976_ _35034_/CLK _31976_/D VGND VGND VPWR VPWR _31976_/Q sky130_fd_sc_hd__dfxtp_1
X_19698_ _19694_/X _19697_/X _19461_/X VGND VGND VPWR VPWR _19699_/D sky130_fd_sc_hd__o21ba_1
XFILLER_225_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33715_ _33779_/CLK _33715_/D VGND VGND VPWR VPWR _33715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18649_ _20201_/A VGND VGND VPWR VPWR _18649_/X sky130_fd_sc_hd__clkbuf_4
X_30927_ _30927_/A VGND VGND VPWR VPWR _35688_/D sky130_fd_sc_hd__clkbuf_1
X_34695_ _34822_/CLK _34695_/D VGND VGND VPWR VPWR _34695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30858_ _23330_/X _35656_/Q _30860_/S VGND VGND VPWR VPWR _30859_/A sky130_fd_sc_hd__mux2_1
X_33646_ _34288_/CLK _33646_/D VGND VGND VPWR VPWR _33646_/Q sky130_fd_sc_hd__dfxtp_1
X_21660_ _33258_/Q _36138_/Q _33130_/Q _33066_/Q _21658_/X _21659_/X VGND VGND VPWR
+ VPWR _21660_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20611_ _22434_/A VGND VGND VPWR VPWR _20611_/X sky130_fd_sc_hd__buf_2
XFILLER_162_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21591_ _33000_/Q _32936_/Q _32872_/Q _32808_/Q _21589_/X _21590_/X VGND VGND VPWR
+ VPWR _21591_/X sky130_fd_sc_hd__mux4_1
X_33577_ _34281_/CLK _33577_/D VGND VGND VPWR VPWR _33577_/Q sky130_fd_sc_hd__dfxtp_1
X_30789_ _23220_/X _35623_/Q _30797_/S VGND VGND VPWR VPWR _30790_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20542_ _20538_/X _20541_/X _20167_/A VGND VGND VPWR VPWR _20543_/D sky130_fd_sc_hd__o21ba_1
X_23330_ input54/X VGND VGND VPWR VPWR _23330_/X sky130_fd_sc_hd__buf_4
XFILLER_178_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35316_ _35574_/CLK _35316_/D VGND VGND VPWR VPWR _35316_/Q sky130_fd_sc_hd__dfxtp_1
X_32528_ _34317_/CLK _32528_/D VGND VGND VPWR VPWR _32528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20473_ _33226_/Q _32586_/Q _35978_/Q _35914_/Q _18375_/X _18376_/X VGND VGND VPWR
+ VPWR _20473_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35247_ _35757_/CLK _35247_/D VGND VGND VPWR VPWR _35247_/Q sky130_fd_sc_hd__dfxtp_1
X_23261_ input31/X VGND VGND VPWR VPWR _23261_/X sky130_fd_sc_hd__clkbuf_4
X_32459_ _35339_/CLK _32459_/D VGND VGND VPWR VPWR _32459_/Q sky130_fd_sc_hd__dfxtp_1
X_25000_ _25000_/A VGND VGND VPWR VPWR _32976_/D sky130_fd_sc_hd__clkbuf_1
X_22212_ _34553_/Q _32441_/Q _34425_/Q _34361_/Q _22178_/X _22179_/X VGND VGND VPWR
+ VPWR _22212_/X sky130_fd_sc_hd__mux4_1
X_23192_ _23192_/A VGND VGND VPWR VPWR _32178_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35178_ _36011_/CLK _35178_/D VGND VGND VPWR VPWR _35178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22143_ _35063_/Q _34999_/Q _34935_/Q _34871_/Q _22109_/X _22110_/X VGND VGND VPWR
+ VPWR _22143_/X sky130_fd_sc_hd__mux4_1
X_34129_ _34260_/CLK _34129_/D VGND VGND VPWR VPWR _34129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26951_ _26950_/X _33847_/Q _26975_/S VGND VGND VPWR VPWR _26952_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22074_ _34294_/Q _34230_/Q _34166_/Q _34102_/Q _22042_/X _22043_/X VGND VGND VPWR
+ VPWR _22074_/X sky130_fd_sc_hd__mux4_1
XTAP_6739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21025_ _33240_/Q _36120_/Q _33112_/Q _33048_/Q _20952_/X _20953_/X VGND VGND VPWR
+ VPWR _21025_/X sky130_fd_sc_hd__mux4_1
X_25902_ _25902_/A VGND VGND VPWR VPWR _33370_/D sky130_fd_sc_hd__clkbuf_1
X_29670_ _35093_/Q _29073_/X _29674_/S VGND VGND VPWR VPWR _29671_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26882_ _26881_/X _33825_/Q _26882_/S VGND VGND VPWR VPWR _26883_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28621_ _26987_/X _34627_/Q _28633_/S VGND VGND VPWR VPWR _28622_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25833_ _25128_/X _33338_/Q _25843_/S VGND VGND VPWR VPWR _25834_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_417_CLK clkbuf_6_35__f_CLK/X VGND VGND VPWR VPWR _34932_/CLK sky130_fd_sc_hd__clkbuf_16
X_28552_ _26884_/X _34594_/Q _28570_/S VGND VGND VPWR VPWR _28553_/A sky130_fd_sc_hd__mux2_1
X_25764_ _25026_/X _33305_/Q _25780_/S VGND VGND VPWR VPWR _25765_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22976_ input25/X VGND VGND VPWR VPWR _22976_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_210_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27503_ _26934_/X _34098_/Q _27509_/S VGND VGND VPWR VPWR _27504_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24715_ _23074_/X _32845_/Q _24715_/S VGND VGND VPWR VPWR _24716_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28483_ _28483_/A VGND VGND VPWR VPWR _34561_/D sky130_fd_sc_hd__clkbuf_1
X_21927_ _21754_/X _21925_/X _21926_/X _21759_/X VGND VGND VPWR VPWR _21927_/X sky130_fd_sc_hd__a22o_1
XFILLER_76_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25695_ _25695_/A VGND VGND VPWR VPWR _33273_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27434_ _26832_/X _34065_/Q _27446_/S VGND VGND VPWR VPWR _27435_/A sky130_fd_sc_hd__mux2_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24646_ _24715_/S VGND VGND VPWR VPWR _24665_/S sky130_fd_sc_hd__buf_6
XFILLER_163_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21858_ _21749_/X _21856_/X _21857_/X _21752_/X VGND VGND VPWR VPWR _21858_/X sky130_fd_sc_hd__a22o_1
XFILLER_208_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20809_ _33490_/Q _33426_/Q _33362_/Q _33298_/Q _20598_/X _20599_/X VGND VGND VPWR
+ VPWR _20809_/X sky130_fd_sc_hd__mux4_1
X_27365_ _27365_/A VGND VGND VPWR VPWR _34032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24577_ _23074_/X _32781_/Q _24577_/S VGND VGND VPWR VPWR _24578_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21789_ _34541_/Q _32429_/Q _34413_/Q _34349_/Q _21472_/X _21473_/X VGND VGND VPWR
+ VPWR _21789_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29104_ input9/X VGND VGND VPWR VPWR _29104_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_106_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26316_ _25044_/X _33567_/Q _26320_/S VGND VGND VPWR VPWR _26317_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23528_ _23028_/X _32318_/Q _23530_/S VGND VGND VPWR VPWR _23529_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27296_ _27296_/A VGND VGND VPWR VPWR _33999_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29035_ _29035_/A VGND VGND VPWR VPWR _34823_/D sky130_fd_sc_hd__clkbuf_1
X_26247_ _26247_/A VGND VGND VPWR VPWR _33534_/D sky130_fd_sc_hd__clkbuf_1
X_23459_ _22926_/X _32285_/Q _23467_/S VGND VGND VPWR VPWR _23460_/A sky130_fd_sc_hd__mux2_1
X_16000_ _33486_/Q _33422_/Q _33358_/Q _33294_/Q _15998_/X _15999_/X VGND VGND VPWR
+ VPWR _16000_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26178_ _26178_/A VGND VGND VPWR VPWR _33501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25129_ _25128_/X _33018_/Q _25144_/S VGND VGND VPWR VPWR _25130_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29937_ _29937_/A VGND VGND VPWR VPWR _35219_/D sky130_fd_sc_hd__clkbuf_1
X_17951_ _17769_/X _17949_/X _17950_/X _17773_/X VGND VGND VPWR VPWR _17951_/X sky130_fd_sc_hd__a22o_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16902_ _16896_/X _16901_/X _16794_/X VGND VGND VPWR VPWR _16910_/C sky130_fd_sc_hd__o21ba_1
XFILLER_239_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17882_ _33025_/Q _32961_/Q _32897_/Q _32833_/Q _17695_/X _17696_/X VGND VGND VPWR
+ VPWR _17882_/X sky130_fd_sc_hd__mux4_1
X_29868_ _35187_/Q _29166_/X _29872_/S VGND VGND VPWR VPWR _29869_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19621_ _19617_/X _19620_/X _19447_/X VGND VGND VPWR VPWR _19629_/C sky130_fd_sc_hd__o21ba_1
XFILLER_4_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28819_ _26881_/X _34721_/Q _28819_/S VGND VGND VPWR VPWR _28820_/A sky130_fd_sc_hd__mux2_1
X_16833_ _34787_/Q _34723_/Q _34659_/Q _34595_/Q _16582_/X _16583_/X VGND VGND VPWR
+ VPWR _16833_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29799_ _35154_/Q _29064_/X _29809_/S VGND VGND VPWR VPWR _29800_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_408_CLK clkbuf_6_33__f_CLK/X VGND VGND VPWR VPWR _35179_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31830_ _31830_/A VGND VGND VPWR VPWR _36116_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19552_ _35567_/Q _35503_/Q _35439_/Q _35375_/Q _19550_/X _19551_/X VGND VGND VPWR
+ VPWR _19552_/X sky130_fd_sc_hd__mux4_1
X_16764_ _16760_/X _16763_/X _16455_/X VGND VGND VPWR VPWR _16765_/D sky130_fd_sc_hd__o21ba_1
XFILLER_111_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18503_ _18499_/X _18502_/X _18400_/X VGND VGND VPWR VPWR _18504_/D sky130_fd_sc_hd__o21ba_1
XFILLER_19_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31761_ _36084_/Q input32/X _31763_/S VGND VGND VPWR VPWR _31762_/A sky130_fd_sc_hd__mux2_1
X_19483_ _33197_/Q _32557_/Q _35949_/Q _35885_/Q _19374_/X _19375_/X VGND VGND VPWR
+ VPWR _19483_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16695_ _33760_/Q _33696_/Q _33632_/Q _33568_/Q _16490_/X _16491_/X VGND VGND VPWR
+ VPWR _16695_/X sky130_fd_sc_hd__mux4_1
XFILLER_206_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30712_ _30712_/A VGND VGND VPWR VPWR _35586_/D sky130_fd_sc_hd__clkbuf_1
X_33500_ _34074_/CLK _33500_/D VGND VGND VPWR VPWR _33500_/Q sky130_fd_sc_hd__dfxtp_1
X_18434_ _18434_/A _18434_/B _18434_/C _18434_/D VGND VGND VPWR VPWR _18435_/A sky130_fd_sc_hd__or4_4
X_31692_ _36051_/Q input56/X _31700_/S VGND VGND VPWR VPWR _31693_/A sky130_fd_sc_hd__mux2_1
X_34480_ _35760_/CLK _34480_/D VGND VGND VPWR VPWR _34480_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_871 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33431_ _34001_/CLK _33431_/D VGND VGND VPWR VPWR _33431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18365_ _20232_/A VGND VGND VPWR VPWR _18365_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30643_ _30733_/S VGND VGND VPWR VPWR _30662_/S sky130_fd_sc_hd__buf_4
XFILLER_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _35761_/Q _35121_/Q _34481_/Q _33841_/Q _17140_/X _17141_/X VGND VGND VPWR
+ VPWR _17316_/X sky130_fd_sc_hd__mux4_1
X_33362_ _33940_/CLK _33362_/D VGND VGND VPWR VPWR _33362_/Q sky130_fd_sc_hd__dfxtp_1
X_36150_ _36150_/CLK _36150_/D VGND VGND VPWR VPWR _36150_/Q sky130_fd_sc_hd__dfxtp_1
X_18296_ _20069_/A VGND VGND VPWR VPWR _20160_/A sky130_fd_sc_hd__buf_12
X_30574_ _23307_/X _35521_/Q _30590_/S VGND VGND VPWR VPWR _30575_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35101_ _35933_/CLK _35101_/D VGND VGND VPWR VPWR _35101_/Q sky130_fd_sc_hd__dfxtp_1
X_32313_ _35320_/CLK _32313_/D VGND VGND VPWR VPWR _32313_/Q sky130_fd_sc_hd__dfxtp_1
X_17247_ _35823_/Q _32200_/Q _35695_/Q _35631_/Q _16960_/X _16961_/X VGND VGND VPWR
+ VPWR _17247_/X sky130_fd_sc_hd__mux4_1
X_33293_ _34316_/CLK _33293_/D VGND VGND VPWR VPWR _33293_/Q sky130_fd_sc_hd__dfxtp_1
X_36081_ _36081_/CLK _36081_/D VGND VGND VPWR VPWR _36081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35032_ _35098_/CLK _35032_/D VGND VGND VPWR VPWR _35032_/Q sky130_fd_sc_hd__dfxtp_1
X_32244_ _34228_/CLK _32244_/D VGND VGND VPWR VPWR _32244_/Q sky130_fd_sc_hd__dfxtp_1
X_17178_ _17174_/X _17177_/X _17136_/X _17137_/X VGND VGND VPWR VPWR _17193_/B sky130_fd_sc_hd__o211a_1
XFILLER_127_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16129_ _16074_/X _16127_/X _16128_/X _16084_/X VGND VGND VPWR VPWR _16129_/X sky130_fd_sc_hd__a22o_1
XFILLER_6_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32175_ _34271_/CLK _32175_/D VGND VGND VPWR VPWR _32175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31126_ _35783_/Q _29228_/X _31130_/S VGND VGND VPWR VPWR _31127_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35934_ _35935_/CLK _35934_/D VGND VGND VPWR VPWR _35934_/Q sky130_fd_sc_hd__dfxtp_1
X_31057_ _35750_/Q _29126_/X _31067_/S VGND VGND VPWR VPWR _31058_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30008_ _30008_/A VGND VGND VPWR VPWR _35253_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19819_ _34295_/Q _34231_/Q _34167_/Q _34103_/Q _19742_/X _19743_/X VGND VGND VPWR
+ VPWR _19819_/X sky130_fd_sc_hd__mux4_1
X_35865_ _35931_/CLK _35865_/D VGND VGND VPWR VPWR _35865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34816_ _34816_/CLK _34816_/D VGND VGND VPWR VPWR _34816_/Q sky130_fd_sc_hd__dfxtp_1
X_22830_ _35788_/Q _35148_/Q _34508_/Q _33868_/Q _20708_/X _20709_/X VGND VGND VPWR
+ VPWR _22830_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35796_ _35797_/CLK _35796_/D VGND VGND VPWR VPWR _35796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22761_ _22757_/X _22760_/X _22434_/A VGND VGND VPWR VPWR _22783_/A sky130_fd_sc_hd__o21ba_1
X_34747_ _35707_/CLK _34747_/D VGND VGND VPWR VPWR _34747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31959_ _35036_/CLK _31959_/D VGND VGND VPWR VPWR _31959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24500_ _22960_/X _32744_/Q _24506_/S VGND VGND VPWR VPWR _24501_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21712_ _35307_/Q _35243_/Q _35179_/Q _32299_/Q _21606_/X _21607_/X VGND VGND VPWR
+ VPWR _21712_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25480_ _33173_/Q _24267_/X _25484_/S VGND VGND VPWR VPWR _25481_/A sky130_fd_sc_hd__mux2_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22692_ _22688_/X _22691_/X _22467_/X VGND VGND VPWR VPWR _22693_/D sky130_fd_sc_hd__o21ba_1
XFILLER_240_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34678_ _34745_/CLK _34678_/D VGND VGND VPWR VPWR _34678_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24431_ input57/X VGND VGND VPWR VPWR _24431_/X sky130_fd_sc_hd__clkbuf_4
X_21643_ _35049_/Q _34985_/Q _34921_/Q _34857_/Q _21403_/X _21404_/X VGND VGND VPWR
+ VPWR _21643_/X sky130_fd_sc_hd__mux4_1
X_33629_ _34142_/CLK _33629_/D VGND VGND VPWR VPWR _33629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27150_ _27011_/X _33931_/Q _27154_/S VGND VGND VPWR VPWR _27151_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24362_ _24362_/A VGND VGND VPWR VPWR _32691_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_30 _32116_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21574_ _21401_/X _21572_/X _21573_/X _21406_/X VGND VGND VPWR VPWR _21574_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_835 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_41 _32118_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 _32126_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26101_ _25125_/X _33465_/Q _26113_/S VGND VGND VPWR VPWR _26102_/A sky130_fd_sc_hd__mux2_1
X_23313_ input49/X VGND VGND VPWR VPWR _23313_/X sky130_fd_sc_hd__buf_4
XANTENNA_63 _32126_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20525_ _32524_/Q _32396_/Q _32076_/Q _36044_/Q _20282_/X _19307_/A VGND VGND VPWR
+ VPWR _20525_/X sky130_fd_sc_hd__mux4_1
X_27081_ _26909_/X _33898_/Q _27083_/S VGND VGND VPWR VPWR _27082_/A sky130_fd_sc_hd__mux2_1
XANTENNA_74 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24293_ _32669_/Q _24292_/X _24305_/S VGND VGND VPWR VPWR _24294_/A sky130_fd_sc_hd__mux2_1
XANTENNA_85 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26032_ _25022_/X _33432_/Q _26050_/S VGND VGND VPWR VPWR _26033_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20456_ _34314_/Q _34250_/Q _34186_/Q _34122_/Q _18345_/X _18346_/X VGND VGND VPWR
+ VPWR _20456_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23244_ input26/X VGND VGND VPWR VPWR _23244_/X sky130_fd_sc_hd__buf_4
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20387_ _35335_/Q _35271_/Q _35207_/Q _32327_/Q _18388_/X _18390_/X VGND VGND VPWR
+ VPWR _20387_/X sky130_fd_sc_hd__mux4_1
X_23175_ input15/X VGND VGND VPWR VPWR _23175_/X sky130_fd_sc_hd__buf_4
XFILLER_238_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22126_ _33271_/Q _36151_/Q _33143_/Q _33079_/Q _22011_/X _22012_/X VGND VGND VPWR
+ VPWR _22126_/X sky130_fd_sc_hd__mux4_1
X_27983_ _27983_/A VGND VGND VPWR VPWR _34324_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_1309 _17061_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput170 _36198_/Q VGND VGND VPWR VPWR D2[24] sky130_fd_sc_hd__buf_2
XFILLER_82_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput181 _36208_/Q VGND VGND VPWR VPWR D2[34] sky130_fd_sc_hd__buf_2
XFILLER_153_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput192 _36218_/Q VGND VGND VPWR VPWR D2[44] sky130_fd_sc_hd__buf_2
XTAP_5802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29722_ _29722_/A VGND VGND VPWR VPWR _35117_/D sky130_fd_sc_hd__clkbuf_1
X_26934_ input30/X VGND VGND VPWR VPWR _26934_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22057_ _35829_/Q _32207_/Q _35701_/Q _35637_/Q _21913_/X _21914_/X VGND VGND VPWR
+ VPWR _22057_/X sky130_fd_sc_hd__mux4_1
XFILLER_248_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21008_ _34519_/Q _32407_/Q _34391_/Q _34327_/Q _20766_/X _20767_/X VGND VGND VPWR
+ VPWR _21008_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29653_ _29653_/A VGND VGND VPWR VPWR _35085_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26865_ _26865_/A VGND VGND VPWR VPWR _33819_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28604_ _26962_/X _34619_/Q _28612_/S VGND VGND VPWR VPWR _28605_/A sky130_fd_sc_hd__mux2_1
X_25816_ _25103_/X _33330_/Q _25822_/S VGND VGND VPWR VPWR _25817_/A sky130_fd_sc_hd__mux2_1
X_29584_ _35052_/Q _29144_/X _29602_/S VGND VGND VPWR VPWR _29585_/A sky130_fd_sc_hd__mux2_1
X_26796_ _26796_/A VGND VGND VPWR VPWR _33793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28535_ _26860_/X _34586_/Q _28549_/S VGND VGND VPWR VPWR _28536_/A sky130_fd_sc_hd__mux2_1
X_25747_ _25001_/X _33297_/Q _25759_/S VGND VGND VPWR VPWR _25748_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1096 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22959_ _22959_/A VGND VGND VPWR VPWR _32039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28466_ _28466_/A VGND VGND VPWR VPWR _34553_/D sky130_fd_sc_hd__clkbuf_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16480_ _34777_/Q _34713_/Q _34649_/Q _34585_/Q _16229_/X _16230_/X VGND VGND VPWR
+ VPWR _16480_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25678_ _25678_/A VGND VGND VPWR VPWR _33265_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27417_ _27417_/A VGND VGND VPWR VPWR _34057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24629_ _24629_/A VGND VGND VPWR VPWR _32803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28397_ _28397_/A VGND VGND VPWR VPWR _34520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18150_ _35081_/Q _35017_/Q _34953_/Q _34889_/Q _17862_/X _17863_/X VGND VGND VPWR
+ VPWR _18150_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27348_ _27348_/A VGND VGND VPWR VPWR _34024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17101_ _33003_/Q _32939_/Q _32875_/Q _32811_/Q _16989_/X _16990_/X VGND VGND VPWR
+ VPWR _17101_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18081_ _15977_/X _18079_/X _18080_/X _15987_/X VGND VGND VPWR VPWR _18081_/X sky130_fd_sc_hd__a22o_1
XFILLER_200_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27279_ _27002_/X _33992_/Q _27281_/S VGND VGND VPWR VPWR _27280_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29018_ _29018_/A VGND VGND VPWR VPWR _34815_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17032_ _35817_/Q _32194_/Q _35689_/Q _35625_/Q _16960_/X _16961_/X VGND VGND VPWR
+ VPWR _17032_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30290_ _35387_/Q _29191_/X _30298_/S VGND VGND VPWR VPWR _30291_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1086 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18983_ _33183_/Q _32543_/Q _35935_/Q _35871_/Q _18668_/X _18669_/X VGND VGND VPWR
+ VPWR _18983_/X sky130_fd_sc_hd__mux4_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _35074_/Q _35010_/Q _34946_/Q _34882_/Q _17862_/X _17863_/X VGND VGND VPWR
+ VPWR _17934_/X sky130_fd_sc_hd__mux4_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33980_ _34171_/CLK _33980_/D VGND VGND VPWR VPWR _33980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32931_ _32994_/CLK _32931_/D VGND VGND VPWR VPWR _32931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17865_ _17865_/A VGND VGND VPWR VPWR _17865_/X sky130_fd_sc_hd__buf_4
XFILLER_227_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19604_ _19502_/X _19602_/X _19603_/X _19505_/X VGND VGND VPWR VPWR _19604_/X sky130_fd_sc_hd__a22o_1
XFILLER_226_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35650_ _35715_/CLK _35650_/D VGND VGND VPWR VPWR _35650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16816_ _34019_/Q _33955_/Q _33891_/Q _32163_/Q _16667_/X _16668_/X VGND VGND VPWR
+ VPWR _16816_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32862_ _35481_/CLK _32862_/D VGND VGND VPWR VPWR _32862_/Q sky130_fd_sc_hd__dfxtp_1
X_17796_ _17796_/A VGND VGND VPWR VPWR _17796_/X sky130_fd_sc_hd__buf_4
XFILLER_4_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1074 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34601_ _34794_/CLK _34601_/D VGND VGND VPWR VPWR _34601_/Q sky130_fd_sc_hd__dfxtp_1
X_31813_ _36109_/Q input60/X _31813_/S VGND VGND VPWR VPWR _31814_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19535_ _19495_/X _19533_/X _19534_/X _19500_/X VGND VGND VPWR VPWR _19535_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35581_ _35581_/CLK _35581_/D VGND VGND VPWR VPWR _35581_/Q sky130_fd_sc_hd__dfxtp_1
X_16747_ _32481_/Q _32353_/Q _32033_/Q _36001_/Q _16570_/X _16711_/X VGND VGND VPWR
+ VPWR _16747_/X sky130_fd_sc_hd__mux4_1
X_32793_ _36119_/CLK _32793_/D VGND VGND VPWR VPWR _32793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34532_ _35042_/CLK _34532_/D VGND VGND VPWR VPWR _34532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16678_ _16674_/X _16677_/X _16430_/X _16431_/X VGND VGND VPWR VPWR _16693_/B sky130_fd_sc_hd__o211a_1
X_31744_ _31813_/S VGND VGND VPWR VPWR _31763_/S sky130_fd_sc_hd__buf_6
X_19466_ _34285_/Q _34221_/Q _34157_/Q _34093_/Q _19389_/X _19390_/X VGND VGND VPWR
+ VPWR _19466_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18417_ _32975_/Q _32911_/Q _32847_/Q _32783_/Q _18333_/X _18335_/X VGND VGND VPWR
+ VPWR _18417_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34463_ _35743_/CLK _34463_/D VGND VGND VPWR VPWR _34463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31675_ _31675_/A VGND VGND VPWR VPWR _36043_/D sky130_fd_sc_hd__clkbuf_1
X_19397_ _32747_/Q _32683_/Q _32619_/Q _36075_/Q _19219_/X _19356_/X VGND VGND VPWR
+ VPWR _19397_/X sky130_fd_sc_hd__mux4_1
XFILLER_188_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36202_ _36202_/CLK _36202_/D VGND VGND VPWR VPWR _36202_/Q sky130_fd_sc_hd__dfxtp_1
X_33414_ _34306_/CLK _33414_/D VGND VGND VPWR VPWR _33414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18348_ _20278_/A VGND VGND VPWR VPWR _20294_/A sky130_fd_sc_hd__buf_12
XFILLER_124_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30626_ _30626_/A VGND VGND VPWR VPWR _35545_/D sky130_fd_sc_hd__clkbuf_1
X_34394_ _34970_/CLK _34394_/D VGND VGND VPWR VPWR _34394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36133_ _36134_/CLK _36133_/D VGND VGND VPWR VPWR _36133_/Q sky130_fd_sc_hd__dfxtp_1
X_33345_ _34305_/CLK _33345_/D VGND VGND VPWR VPWR _33345_/Q sky130_fd_sc_hd__dfxtp_1
X_18279_ _18357_/A VGND VGND VPWR VPWR _20202_/A sky130_fd_sc_hd__buf_12
X_30557_ _23280_/X _35513_/Q _30569_/S VGND VGND VPWR VPWR _30558_/A sky130_fd_sc_hd__mux2_1
X_20310_ _20208_/X _20308_/X _20309_/X _20211_/X VGND VGND VPWR VPWR _20310_/X sky130_fd_sc_hd__a22o_1
XFILLER_198_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21290_ _35039_/Q _34975_/Q _34911_/Q _34847_/Q _21050_/X _21051_/X VGND VGND VPWR
+ VPWR _21290_/X sky130_fd_sc_hd__mux4_1
Xinput50 DW[54] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_16
X_36064_ _36067_/CLK _36064_/D VGND VGND VPWR VPWR _36064_/Q sky130_fd_sc_hd__dfxtp_1
X_33276_ _36156_/CLK _33276_/D VGND VGND VPWR VPWR _33276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput61 DW[6] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__buf_8
X_30488_ _23117_/X _35480_/Q _30506_/S VGND VGND VPWR VPWR _30489_/A sky130_fd_sc_hd__mux2_1
Xinput72 R2[1] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput83 RW[0] VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__buf_4
X_35015_ _35781_/CLK _35015_/D VGND VGND VPWR VPWR _35015_/Q sky130_fd_sc_hd__dfxtp_1
X_20241_ _20201_/X _20239_/X _20240_/X _20206_/X VGND VGND VPWR VPWR _20241_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32227_ _35848_/CLK _32227_/D VGND VGND VPWR VPWR _32227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20172_ _34305_/Q _34241_/Q _34177_/Q _34113_/Q _20095_/X _20096_/X VGND VGND VPWR
+ VPWR _20172_/X sky130_fd_sc_hd__mux4_1
X_32158_ _36200_/CLK _32158_/D VGND VGND VPWR VPWR _32158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31109_ _35775_/Q _29203_/X _31109_/S VGND VGND VPWR VPWR _31110_/A sky130_fd_sc_hd__mux2_1
X_24980_ _24980_/A VGND VGND VPWR VPWR _32969_/D sky130_fd_sc_hd__clkbuf_1
X_32089_ _35040_/CLK _32089_/D VGND VGND VPWR VPWR _32089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35917_ _35917_/CLK _35917_/D VGND VGND VPWR VPWR _35917_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23931_ _23016_/X _32506_/Q _23941_/S VGND VGND VPWR VPWR _23932_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26650_ _25137_/X _33725_/Q _26654_/S VGND VGND VPWR VPWR _26651_/A sky130_fd_sc_hd__mux2_1
XTAP_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35848_ _35848_/CLK _35848_/D VGND VGND VPWR VPWR _35848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23862_ _22914_/X _32473_/Q _23878_/S VGND VGND VPWR VPWR _23863_/A sky130_fd_sc_hd__mux2_1
XTAP_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25601_ _25601_/A VGND VGND VPWR VPWR _31140_/B sky130_fd_sc_hd__buf_8
XFILLER_84_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22813_ _22813_/A _22813_/B _22813_/C _22813_/D VGND VGND VPWR VPWR _22814_/A sky130_fd_sc_hd__or4_4
XANTENNA_707 _22532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26581_ _25035_/X _33692_/Q _26591_/S VGND VGND VPWR VPWR _26582_/A sky130_fd_sc_hd__mux2_1
X_35779_ _35779_/CLK _35779_/D VGND VGND VPWR VPWR _35779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23793_ _23013_/X _32441_/Q _23805_/S VGND VGND VPWR VPWR _23794_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_718 _22453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_729 _20940_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28320_ _28320_/A VGND VGND VPWR VPWR _34484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25532_ _25532_/A VGND VGND VPWR VPWR _33197_/D sky130_fd_sc_hd__clkbuf_1
X_22744_ _20597_/X _22742_/X _22743_/X _20603_/X VGND VGND VPWR VPWR _22744_/X sky130_fd_sc_hd__a22o_1
XFILLER_197_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28251_ _28251_/A VGND VGND VPWR VPWR _34451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1029 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25463_ _25463_/A VGND VGND VPWR VPWR _30600_/B sky130_fd_sc_hd__buf_6
XFILLER_240_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22675_ _32519_/Q _32391_/Q _32071_/Q _36039_/Q _22582_/X _22370_/X VGND VGND VPWR
+ VPWR _22675_/X sky130_fd_sc_hd__mux4_1
XFILLER_198_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27202_ _26888_/X _33955_/Q _27218_/S VGND VGND VPWR VPWR _27203_/A sky130_fd_sc_hd__mux2_1
X_24414_ _32708_/Q _24413_/X _24429_/S VGND VGND VPWR VPWR _24415_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28182_ _26937_/X _34419_/Q _28186_/S VGND VGND VPWR VPWR _28183_/A sky130_fd_sc_hd__mux2_1
X_21626_ _33257_/Q _36137_/Q _33129_/Q _33065_/Q _21305_/X _21306_/X VGND VGND VPWR
+ VPWR _21626_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25394_ _25091_/X _33134_/Q _25408_/S VGND VGND VPWR VPWR _25395_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27133_ _27133_/A VGND VGND VPWR VPWR _33922_/D sky130_fd_sc_hd__clkbuf_1
X_24345_ input26/X VGND VGND VPWR VPWR _24345_/X sky130_fd_sc_hd__clkbuf_8
X_21557_ _32999_/Q _32935_/Q _32871_/Q _32807_/Q _21236_/X _21237_/X VGND VGND VPWR
+ VPWR _21557_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20508_ _18344_/X _20506_/X _20507_/X _18354_/X VGND VGND VPWR VPWR _20508_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27064_ _27154_/S VGND VGND VPWR VPWR _27083_/S sky130_fd_sc_hd__buf_4
X_24276_ input2/X VGND VGND VPWR VPWR _24276_/X sky130_fd_sc_hd__buf_4
X_21488_ _33253_/Q _36133_/Q _33125_/Q _33061_/Q _21305_/X _21306_/X VGND VGND VPWR
+ VPWR _21488_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26015_ _24998_/X _33424_/Q _26029_/S VGND VGND VPWR VPWR _26016_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23227_ _23227_/A VGND VGND VPWR VPWR _32193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20439_ _35849_/Q _32229_/Q _35721_/Q _35657_/Q _18289_/X _18291_/X VGND VGND VPWR
+ VPWR _20439_/X sky130_fd_sc_hd__mux4_1
XTAP_7012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23158_ _23158_/A VGND VGND VPWR VPWR _29924_/A sky130_fd_sc_hd__buf_6
XTAP_7056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1106 _17471_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1117 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22109_ _22462_/A VGND VGND VPWR VPWR _22109_/X sky130_fd_sc_hd__buf_4
XFILLER_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1128 _31996_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15980_ _17902_/A VGND VGND VPWR VPWR _15980_/X sky130_fd_sc_hd__buf_8
XTAP_6355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23089_ _23089_/A VGND VGND VPWR VPWR _32142_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_1139 _20134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27966_ _34317_/Q _24440_/X _27966_/S VGND VGND VPWR VPWR _27967_/A sky130_fd_sc_hd__mux2_1
XTAP_6366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29705_ _29705_/A VGND VGND VPWR VPWR _35109_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26917_ _26915_/X _33836_/Q _26944_/S VGND VGND VPWR VPWR _26918_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27897_ _27966_/S VGND VGND VPWR VPWR _27916_/S sky130_fd_sc_hd__buf_6
XFILLER_212_1158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29636_ _35077_/Q _29222_/X _29644_/S VGND VGND VPWR VPWR _29637_/A sky130_fd_sc_hd__mux2_1
XTAP_5698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17650_ _17650_/A _17650_/B _17650_/C _17650_/D VGND VGND VPWR VPWR _17651_/A sky130_fd_sc_hd__or4_4
XFILLER_208_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26848_ _26847_/X _33814_/Q _26851_/S VGND VGND VPWR VPWR _26849_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16601_ _33245_/Q _36125_/Q _33117_/Q _33053_/Q _16352_/X _16353_/X VGND VGND VPWR
+ VPWR _16601_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17581_ _35064_/Q _35000_/Q _34936_/Q _34872_/Q _17509_/X _17510_/X VGND VGND VPWR
+ VPWR _17581_/X sky130_fd_sc_hd__mux4_1
X_26779_ _26779_/A VGND VGND VPWR VPWR _33785_/D sky130_fd_sc_hd__clkbuf_1
X_29567_ _35044_/Q _29120_/X _29581_/S VGND VGND VPWR VPWR _29568_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16532_ _16496_/X _16530_/X _16531_/X _16499_/X VGND VGND VPWR VPWR _16532_/X sky130_fd_sc_hd__a22o_1
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19320_ _20146_/A VGND VGND VPWR VPWR _19320_/X sky130_fd_sc_hd__buf_6
XFILLER_186_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28518_ _26835_/X _34578_/Q _28528_/S VGND VGND VPWR VPWR _28519_/A sky130_fd_sc_hd__mux2_1
X_29498_ _29498_/A VGND VGND VPWR VPWR _35011_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16463_ _34009_/Q _33945_/Q _33881_/Q _32153_/Q _16314_/X _16315_/X VGND VGND VPWR
+ VPWR _16463_/X sky130_fd_sc_hd__mux4_1
X_19251_ _19149_/X _19249_/X _19250_/X _19152_/X VGND VGND VPWR VPWR _19251_/X sky130_fd_sc_hd__a22o_1
XFILLER_204_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28449_ _28449_/A VGND VGND VPWR VPWR _34545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18202_ _35595_/Q _35531_/Q _35467_/Q _35403_/Q _17956_/X _17957_/X VGND VGND VPWR
+ VPWR _18202_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31460_ _23199_/X _35941_/Q _31472_/S VGND VGND VPWR VPWR _31461_/A sky130_fd_sc_hd__mux2_1
X_19182_ _19142_/X _19180_/X _19181_/X _19147_/X VGND VGND VPWR VPWR _19182_/X sky130_fd_sc_hd__a22o_1
XPHY_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16394_ _32471_/Q _32343_/Q _32023_/Q _35991_/Q _16217_/X _16358_/X VGND VGND VPWR
+ VPWR _16394_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18133_ _33289_/Q _36169_/Q _33161_/Q _33097_/Q _16028_/X _17157_/A VGND VGND VPWR
+ VPWR _18133_/X sky130_fd_sc_hd__mux4_1
X_30411_ _23264_/X _35444_/Q _30413_/S VGND VGND VPWR VPWR _30412_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_991 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31391_ _31391_/A VGND VGND VPWR VPWR _35908_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1036 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18064_ _18064_/A VGND VGND VPWR VPWR _32006_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_184_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30342_ _23102_/X _35411_/Q _30350_/S VGND VGND VPWR VPWR _30343_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33130_ _36137_/CLK _33130_/D VGND VGND VPWR VPWR _33130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17015_ _17015_/A VGND VGND VPWR VPWR _31976_/D sky130_fd_sc_hd__clkbuf_1
X_33061_ _36134_/CLK _33061_/D VGND VGND VPWR VPWR _33061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30273_ _35379_/Q _29166_/X _30277_/S VGND VGND VPWR VPWR _30274_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32012_ _36194_/CLK _32012_/D VGND VGND VPWR VPWR _32012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18966_ _33503_/Q _33439_/Q _33375_/Q _33311_/Q _18717_/X _18718_/X VGND VGND VPWR
+ VPWR _18966_/X sky130_fd_sc_hd__mux4_1
XFILLER_26_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17917_ _32514_/Q _32386_/Q _32066_/Q _36034_/Q _17629_/X _17770_/X VGND VGND VPWR
+ VPWR _17917_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33963_ _36136_/CLK _33963_/D VGND VGND VPWR VPWR _33963_/Q sky130_fd_sc_hd__dfxtp_1
X_18897_ _34013_/Q _33949_/Q _33885_/Q _32157_/Q _18614_/X _18615_/X VGND VGND VPWR
+ VPWR _18897_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35702_ _35831_/CLK _35702_/D VGND VGND VPWR VPWR _35702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32914_ _32978_/CLK _32914_/D VGND VGND VPWR VPWR _32914_/Q sky130_fd_sc_hd__dfxtp_1
X_17848_ _35776_/Q _35136_/Q _34496_/Q _33856_/Q _17846_/X _17847_/X VGND VGND VPWR
+ VPWR _17848_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33894_ _34087_/CLK _33894_/D VGND VGND VPWR VPWR _33894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35633_ _35954_/CLK _35633_/D VGND VGND VPWR VPWR _35633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32845_ _35919_/CLK _32845_/D VGND VGND VPWR VPWR _32845_/Q sky130_fd_sc_hd__dfxtp_1
X_17779_ _35582_/Q _35518_/Q _35454_/Q _35390_/Q _17603_/X _17604_/X VGND VGND VPWR
+ VPWR _17779_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19518_ _35566_/Q _35502_/Q _35438_/Q _35374_/Q _19197_/X _19198_/X VGND VGND VPWR
+ VPWR _19518_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35564_ _35564_/CLK _35564_/D VGND VGND VPWR VPWR _35564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32776_ _36169_/CLK _32776_/D VGND VGND VPWR VPWR _32776_/Q sky130_fd_sc_hd__dfxtp_1
X_20790_ _20644_/X _20788_/X _20789_/X _20654_/X VGND VGND VPWR VPWR _20790_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34515_ _34967_/CLK _34515_/D VGND VGND VPWR VPWR _34515_/Q sky130_fd_sc_hd__dfxtp_1
X_19449_ _19449_/A VGND VGND VPWR VPWR _19449_/X sky130_fd_sc_hd__clkbuf_4
X_31727_ _31727_/A VGND VGND VPWR VPWR _36067_/D sky130_fd_sc_hd__clkbuf_1
X_35495_ _35750_/CLK _35495_/D VGND VGND VPWR VPWR _35495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_1160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22460_ _22460_/A VGND VGND VPWR VPWR _22460_/X sky130_fd_sc_hd__buf_4
X_34446_ _35728_/CLK _34446_/D VGND VGND VPWR VPWR _34446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31658_ _36035_/Q input49/X _31670_/S VGND VGND VPWR VPWR _31659_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21411_ _21411_/A VGND VGND VPWR VPWR _36194_/D sky130_fd_sc_hd__clkbuf_1
X_30609_ _30609_/A VGND VGND VPWR VPWR _35537_/D sky130_fd_sc_hd__clkbuf_1
X_34377_ _35337_/CLK _34377_/D VGND VGND VPWR VPWR _34377_/Q sky130_fd_sc_hd__dfxtp_1
X_22391_ _22387_/X _22390_/X _22114_/X VGND VGND VPWR VPWR _22392_/D sky130_fd_sc_hd__o21ba_1
X_31589_ _36002_/Q input13/X _31607_/S VGND VGND VPWR VPWR _31590_/A sky130_fd_sc_hd__mux2_1
X_36116_ _36116_/CLK _36116_/D VGND VGND VPWR VPWR _36116_/Q sky130_fd_sc_hd__dfxtp_1
X_24130_ _24130_/A VGND VGND VPWR VPWR _32599_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21342_ _21096_/X _21340_/X _21341_/X _21099_/X VGND VGND VPWR VPWR _21342_/X sky130_fd_sc_hd__a22o_1
XFILLER_15_1480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33328_ _33520_/CLK _33328_/D VGND VGND VPWR VPWR _33328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36047_ _36048_/CLK _36047_/D VGND VGND VPWR VPWR _36047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24061_ _23007_/X _32567_/Q _24077_/S VGND VGND VPWR VPWR _24062_/A sky130_fd_sc_hd__mux2_1
X_33259_ _34283_/CLK _33259_/D VGND VGND VPWR VPWR _33259_/Q sky130_fd_sc_hd__dfxtp_1
X_21273_ _33247_/Q _36127_/Q _33119_/Q _33055_/Q _20952_/X _20953_/X VGND VGND VPWR
+ VPWR _21273_/X sky130_fd_sc_hd__mux4_1
X_23012_ _23012_/A VGND VGND VPWR VPWR _32056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20224_ _35586_/Q _35522_/Q _35458_/Q _35394_/Q _19903_/X _19904_/X VGND VGND VPWR
+ VPWR _20224_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27820_ _27820_/A VGND VGND VPWR VPWR _34247_/D sky130_fd_sc_hd__clkbuf_1
X_20155_ _20155_/A VGND VGND VPWR VPWR _20155_/X sky130_fd_sc_hd__buf_4
XFILLER_131_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24963_ _23038_/X _32961_/Q _24979_/S VGND VGND VPWR VPWR _24964_/A sky130_fd_sc_hd__mux2_1
X_20086_ _35326_/Q _35262_/Q _35198_/Q _32318_/Q _20012_/X _20013_/X VGND VGND VPWR
+ VPWR _20086_/X sky130_fd_sc_hd__mux4_1
XTAP_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27751_ _27751_/A VGND VGND VPWR VPWR _34214_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26702_ _33749_/Q _24267_/X _26706_/S VGND VGND VPWR VPWR _26703_/A sky130_fd_sc_hd__mux2_1
XTAP_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23914_ _22991_/X _32498_/Q _23920_/S VGND VGND VPWR VPWR _23915_/A sky130_fd_sc_hd__mux2_1
X_27682_ _34182_/Q _24419_/X _27688_/S VGND VGND VPWR VPWR _27683_/A sky130_fd_sc_hd__mux2_1
XTAP_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24894_ _24894_/A VGND VGND VPWR VPWR _32928_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29421_ _23139_/X _34975_/Q _29425_/S VGND VGND VPWR VPWR _29422_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26633_ _25112_/X _33717_/Q _26633_/S VGND VGND VPWR VPWR _26634_/A sky130_fd_sc_hd__mux2_1
X_23845_ _22889_/X _32465_/Q _23857_/S VGND VGND VPWR VPWR _23846_/A sky130_fd_sc_hd__mux2_1
XTAP_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_504 _17825_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_515 _17938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_526 _18033_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_537 _20096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26564_ _25010_/X _33684_/Q _26570_/S VGND VGND VPWR VPWR _26565_/A sky130_fd_sc_hd__mux2_1
X_29352_ _29352_/A VGND VGND VPWR VPWR _34942_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23776_ _22988_/X _32433_/Q _23784_/S VGND VGND VPWR VPWR _23777_/A sky130_fd_sc_hd__mux2_1
XANTENNA_548 _20162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_559 _20158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20988_ _34007_/Q _33943_/Q _33879_/Q _32151_/Q _20914_/X _20915_/X VGND VGND VPWR
+ VPWR _20988_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25515_ _25515_/A VGND VGND VPWR VPWR _33189_/D sky130_fd_sc_hd__clkbuf_1
X_28303_ _34476_/Q _24338_/X _28321_/S VGND VGND VPWR VPWR _28304_/A sky130_fd_sc_hd__mux2_1
X_22727_ _22501_/X _22725_/X _22726_/X _22506_/X VGND VGND VPWR VPWR _22727_/X sky130_fd_sc_hd__a22o_1
X_29283_ _29283_/A VGND VGND VPWR VPWR _34909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26495_ _25109_/X _33652_/Q _26497_/S VGND VGND VPWR VPWR _26496_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28234_ _27014_/X _34444_/Q _28236_/S VGND VGND VPWR VPWR _28235_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25446_ _25168_/X _33159_/Q _25450_/S VGND VGND VPWR VPWR _25447_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22658_ _22455_/X _22656_/X _22657_/X _22458_/X VGND VGND VPWR VPWR _22658_/X sky130_fd_sc_hd__a22o_1
XFILLER_199_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28165_ _26912_/X _34411_/Q _28165_/S VGND VGND VPWR VPWR _28166_/A sky130_fd_sc_hd__mux2_1
X_21609_ _21396_/X _21605_/X _21608_/X _21399_/X VGND VGND VPWR VPWR _21609_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25377_ _25066_/X _33126_/Q _25387_/S VGND VGND VPWR VPWR _25378_/A sky130_fd_sc_hd__mux2_1
X_22589_ _22300_/X _22587_/X _22588_/X _22303_/X VGND VGND VPWR VPWR _22589_/X sky130_fd_sc_hd__a22o_1
XFILLER_194_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27116_ _27116_/A VGND VGND VPWR VPWR _33914_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24328_ _24328_/A VGND VGND VPWR VPWR _32680_/D sky130_fd_sc_hd__clkbuf_1
X_28096_ _28096_/A VGND VGND VPWR VPWR _34378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27047_ _27047_/A VGND VGND VPWR VPWR _33881_/D sky130_fd_sc_hd__clkbuf_1
X_24259_ _32658_/Q _24258_/X _24274_/S VGND VGND VPWR VPWR _24260_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18820_ _19173_/A VGND VGND VPWR VPWR _18820_/X sky130_fd_sc_hd__buf_4
XTAP_6130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28998_ _28998_/A VGND VGND VPWR VPWR _29017_/S sky130_fd_sc_hd__buf_4
XFILLER_62_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18751_ _19457_/A VGND VGND VPWR VPWR _18751_/X sky130_fd_sc_hd__buf_4
X_27949_ _27949_/A VGND VGND VPWR VPWR _34308_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17702_ _35772_/Q _35132_/Q _34492_/Q _33852_/Q _17493_/X _17494_/X VGND VGND VPWR
+ VPWR _17702_/X sky130_fd_sc_hd__mux4_1
XFILLER_237_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18682_ _33751_/Q _33687_/Q _33623_/Q _33559_/Q _18437_/X _18438_/X VGND VGND VPWR
+ VPWR _18682_/X sky130_fd_sc_hd__mux4_1
XTAP_5484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30960_ _35704_/Q _29182_/X _30974_/S VGND VGND VPWR VPWR _30961_/A sky130_fd_sc_hd__mux2_1
XTAP_5495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29619_ _35069_/Q _29197_/X _29623_/S VGND VGND VPWR VPWR _29620_/A sky130_fd_sc_hd__mux2_1
X_17633_ _17628_/X _17632_/X _17489_/X _17490_/X VGND VGND VPWR VPWR _17650_/B sky130_fd_sc_hd__o211a_1
XFILLER_236_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30891_ _30891_/A VGND VGND VPWR VPWR _35671_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32630_ _36086_/CLK _32630_/D VGND VGND VPWR VPWR _32630_/Q sky130_fd_sc_hd__dfxtp_1
X_17564_ _32504_/Q _32376_/Q _32056_/Q _36024_/Q _17276_/X _17417_/X VGND VGND VPWR
+ VPWR _17564_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19303_ _19299_/X _19300_/X _19301_/X _19302_/X VGND VGND VPWR VPWR _19303_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16515_ _16511_/X _16514_/X _16441_/X VGND VGND VPWR VPWR _16525_/C sky130_fd_sc_hd__o21ba_1
XFILLER_56_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32561_ _35889_/CLK _32561_/D VGND VGND VPWR VPWR _32561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17495_ _35766_/Q _35126_/Q _34486_/Q _33846_/Q _17493_/X _17494_/X VGND VGND VPWR
+ VPWR _17495_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34300_ _36157_/CLK _34300_/D VGND VGND VPWR VPWR _34300_/Q sky130_fd_sc_hd__dfxtp_1
X_31512_ _23297_/X _35966_/Q _31514_/S VGND VGND VPWR VPWR _31513_/A sky130_fd_sc_hd__mux2_1
X_19234_ _19230_/X _19233_/X _19094_/X VGND VGND VPWR VPWR _19244_/C sky130_fd_sc_hd__o21ba_1
X_35280_ _35280_/CLK _35280_/D VGND VGND VPWR VPWR _35280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16446_ _17152_/A VGND VGND VPWR VPWR _16446_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_220_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32492_ _36013_/CLK _32492_/D VGND VGND VPWR VPWR _32492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34231_ _34295_/CLK _34231_/D VGND VGND VPWR VPWR _34231_/Q sky130_fd_sc_hd__dfxtp_1
X_16377_ _35030_/Q _34966_/Q _34902_/Q _34838_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _16377_/X sky130_fd_sc_hd__mux4_1
X_19165_ _35556_/Q _35492_/Q _35428_/Q _35364_/Q _18844_/X _18845_/X VGND VGND VPWR
+ VPWR _19165_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31443_ _23133_/X _35933_/Q _31451_/S VGND VGND VPWR VPWR _31444_/A sky130_fd_sc_hd__mux2_1
X_18116_ _34824_/Q _34760_/Q _34696_/Q _34632_/Q _17994_/X _17995_/X VGND VGND VPWR
+ VPWR _18116_/X sky130_fd_sc_hd__mux4_1
X_31374_ _31374_/A VGND VGND VPWR VPWR _35900_/D sky130_fd_sc_hd__clkbuf_1
X_34162_ _35765_/CLK _34162_/D VGND VGND VPWR VPWR _34162_/Q sky130_fd_sc_hd__dfxtp_1
X_19096_ _19449_/A VGND VGND VPWR VPWR _19096_/X sky130_fd_sc_hd__buf_4
XFILLER_117_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30325_ _35404_/Q _29243_/X _30327_/S VGND VGND VPWR VPWR _30326_/A sky130_fd_sc_hd__mux2_1
X_33113_ _36059_/CLK _33113_/D VGND VGND VPWR VPWR _33113_/Q sky130_fd_sc_hd__dfxtp_1
X_18047_ _17769_/X _18045_/X _18046_/X _17773_/X VGND VGND VPWR VPWR _18047_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34093_ _35252_/CLK _34093_/D VGND VGND VPWR VPWR _34093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33044_ _36117_/CLK _33044_/D VGND VGND VPWR VPWR _33044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30256_ _35371_/Q _29141_/X _30256_/S VGND VGND VPWR VPWR _30257_/A sky130_fd_sc_hd__mux2_1
X_30187_ _30187_/A VGND VGND VPWR VPWR _35338_/D sky130_fd_sc_hd__clkbuf_1
X_19998_ _19716_/X _19994_/X _19997_/X _19720_/X VGND VGND VPWR VPWR _19998_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18949_ _20165_/A VGND VGND VPWR VPWR _18949_/X sky130_fd_sc_hd__clkbuf_4
X_34995_ _34997_/CLK _34995_/D VGND VGND VPWR VPWR _34995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21960_ _22313_/A VGND VGND VPWR VPWR _21960_/X sky130_fd_sc_hd__buf_4
XFILLER_80_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33946_ _33946_/CLK _33946_/D VGND VGND VPWR VPWR _33946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20911_ _34261_/Q _34197_/Q _34133_/Q _34069_/Q _20605_/X _20607_/X VGND VGND VPWR
+ VPWR _20911_/X sky130_fd_sc_hd__mux4_1
X_33877_ _35280_/CLK _33877_/D VGND VGND VPWR VPWR _33877_/Q sky130_fd_sc_hd__dfxtp_1
X_21891_ _35312_/Q _35248_/Q _35184_/Q _32304_/Q _21606_/X _21607_/X VGND VGND VPWR
+ VPWR _21891_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35616_ _35809_/CLK _35616_/D VGND VGND VPWR VPWR _35616_/Q sky130_fd_sc_hd__dfxtp_1
X_23630_ _32365_/Q _23241_/X _23646_/S VGND VGND VPWR VPWR _23631_/A sky130_fd_sc_hd__mux2_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20842_ _20736_/X _20840_/X _20841_/X _20741_/X VGND VGND VPWR VPWR _20842_/X sky130_fd_sc_hd__a22o_1
XFILLER_214_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32828_ _36029_/CLK _32828_/D VGND VGND VPWR VPWR _32828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23561_ input83/X _23561_/B VGND VGND VPWR VPWR _31680_/B sky130_fd_sc_hd__nand2_8
X_35547_ _35933_/CLK _35547_/D VGND VGND VPWR VPWR _35547_/Q sky130_fd_sc_hd__dfxtp_1
X_20773_ _20773_/A VGND VGND VPWR VPWR _36176_/D sky130_fd_sc_hd__clkbuf_1
X_32759_ _36088_/CLK _32759_/D VGND VGND VPWR VPWR _32759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25300_ _25153_/X _33090_/Q _25314_/S VGND VGND VPWR VPWR _25301_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22512_ _22508_/X _22509_/X _22510_/X _22511_/X VGND VGND VPWR VPWR _22512_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26280_ _26412_/S VGND VGND VPWR VPWR _26299_/S sky130_fd_sc_hd__buf_4
XFILLER_50_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35478_ _35927_/CLK _35478_/D VGND VGND VPWR VPWR _35478_/Q sky130_fd_sc_hd__dfxtp_1
X_23492_ _23492_/A VGND VGND VPWR VPWR _32300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25231_ _25231_/A VGND VGND VPWR VPWR _33057_/D sky130_fd_sc_hd__clkbuf_1
X_22443_ _22443_/A VGND VGND VPWR VPWR _22443_/X sky130_fd_sc_hd__buf_4
X_34429_ _35581_/CLK _34429_/D VGND VGND VPWR VPWR _34429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25162_ input51/X VGND VGND VPWR VPWR _25162_/X sky130_fd_sc_hd__clkbuf_4
X_22374_ _22369_/X _22371_/X _22372_/X _22373_/X VGND VGND VPWR VPWR _22374_/X sky130_fd_sc_hd__a22o_1
XFILLER_159_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24113_ _22883_/X _32591_/Q _24129_/S VGND VGND VPWR VPWR _24114_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_1034 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21325_ _21319_/X _21324_/X _21041_/X VGND VGND VPWR VPWR _21333_/C sky130_fd_sc_hd__o21ba_1
X_25093_ _25093_/A VGND VGND VPWR VPWR _33006_/D sky130_fd_sc_hd__clkbuf_1
X_29970_ _35235_/Q _29117_/X _29986_/S VGND VGND VPWR VPWR _29971_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28921_ _34769_/Q _24255_/X _28933_/S VGND VGND VPWR VPWR _28922_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24044_ _22982_/X _32559_/Q _24056_/S VGND VGND VPWR VPWR _24045_/A sky130_fd_sc_hd__mux2_1
X_21256_ _21043_/X _21252_/X _21255_/X _21046_/X VGND VGND VPWR VPWR _21256_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_6_47__f_CLK clkbuf_5_23_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_47__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_20207_ _20201_/X _20204_/X _20205_/X _20206_/X VGND VGND VPWR VPWR _20207_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28852_ _28852_/A VGND VGND VPWR VPWR _34736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21187_ _34524_/Q _32412_/Q _34396_/Q _34332_/Q _21119_/X _21120_/X VGND VGND VPWR
+ VPWR _21187_/X sky130_fd_sc_hd__mux4_1
X_27803_ _27803_/A VGND VGND VPWR VPWR _34239_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20138_ _20061_/X _20136_/X _20137_/X _20067_/X VGND VGND VPWR VPWR _20138_/X sky130_fd_sc_hd__a22o_1
X_25995_ _25168_/X _33415_/Q _25999_/S VGND VGND VPWR VPWR _25996_/A sky130_fd_sc_hd__mux2_1
X_28783_ _28783_/A VGND VGND VPWR VPWR _34703_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20069_ _20069_/A VGND VGND VPWR VPWR _20069_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24946_ _23013_/X _32953_/Q _24958_/S VGND VGND VPWR VPWR _24947_/A sky130_fd_sc_hd__mux2_1
X_27734_ _27734_/A VGND VGND VPWR VPWR _34206_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27665_ _34174_/Q _24394_/X _27667_/S VGND VGND VPWR VPWR _27666_/A sky130_fd_sc_hd__mux2_1
X_24877_ _22910_/X _32920_/Q _24895_/S VGND VGND VPWR VPWR _24878_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_301 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_312 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29404_ _23114_/X _34967_/Q _29404_/S VGND VGND VPWR VPWR _29405_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23828_ _23065_/X _32458_/Q _23834_/S VGND VGND VPWR VPWR _23829_/A sky130_fd_sc_hd__mux2_1
XANTENNA_323 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26616_ _26616_/A VGND VGND VPWR VPWR _33708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_334 _32141_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27596_ _34141_/Q _24292_/X _27604_/S VGND VGND VPWR VPWR _27597_/A sky130_fd_sc_hd__mux2_1
XTAP_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_345 _36205_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_356 _36207_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_367 _36207_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26547_ _25186_/X _33677_/Q _26547_/S VGND VGND VPWR VPWR _26548_/A sky130_fd_sc_hd__mux2_1
X_29335_ _23270_/X _34934_/Q _29353_/S VGND VGND VPWR VPWR _29336_/A sky130_fd_sc_hd__mux2_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_378 _36208_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23759_ _22963_/X _32425_/Q _23763_/S VGND VGND VPWR VPWR _23760_/A sky130_fd_sc_hd__mux2_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_389 _36209_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _17712_/A VGND VGND VPWR VPWR _16300_/X sky130_fd_sc_hd__buf_6
XFILLER_13_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17280_ _17275_/X _17279_/X _17136_/X _17137_/X VGND VGND VPWR VPWR _17297_/B sky130_fd_sc_hd__o211a_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29266_ _29266_/A VGND VGND VPWR VPWR _34901_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26478_ _26547_/S VGND VGND VPWR VPWR _26497_/S sky130_fd_sc_hd__buf_6
XFILLER_158_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16231_ _34770_/Q _34706_/Q _34642_/Q _34578_/Q _16229_/X _16230_/X VGND VGND VPWR
+ VPWR _16231_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28217_ _28217_/A VGND VGND VPWR VPWR _34435_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25429_ _25143_/X _33151_/Q _25429_/S VGND VGND VPWR VPWR _25430_/A sky130_fd_sc_hd__mux2_1
X_29197_ input42/X VGND VGND VPWR VPWR _29197_/X sky130_fd_sc_hd__clkbuf_4
X_16162_ _16158_/X _16161_/X _16071_/X VGND VGND VPWR VPWR _16172_/C sky130_fd_sc_hd__o21ba_1
X_28148_ _28148_/A VGND VGND VPWR VPWR _34402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28079_ _26984_/X _34370_/Q _28093_/S VGND VGND VPWR VPWR _28080_/A sky130_fd_sc_hd__mux2_1
X_16093_ _17770_/A VGND VGND VPWR VPWR _17157_/A sky130_fd_sc_hd__buf_12
XFILLER_5_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30110_ _30110_/A VGND VGND VPWR VPWR _35301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19921_ _33530_/Q _33466_/Q _33402_/Q _33338_/Q _19776_/X _19777_/X VGND VGND VPWR
+ VPWR _19921_/X sky130_fd_sc_hd__mux4_1
X_31090_ _31138_/S VGND VGND VPWR VPWR _31109_/S sky130_fd_sc_hd__buf_4
XFILLER_29_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30041_ _35269_/Q _29222_/X _30049_/S VGND VGND VPWR VPWR _30042_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19852_ _34296_/Q _34232_/Q _34168_/Q _34104_/Q _19742_/X _19743_/X VGND VGND VPWR
+ VPWR _19852_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_917 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_150_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _35787_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18803_ _33242_/Q _36122_/Q _33114_/Q _33050_/Q _18652_/X _18653_/X VGND VGND VPWR
+ VPWR _18803_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_1389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19783_ _32758_/Q _32694_/Q _32630_/Q _36086_/Q _19572_/X _19709_/X VGND VGND VPWR
+ VPWR _19783_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16995_ _35816_/Q _32192_/Q _35688_/Q _35624_/Q _16960_/X _16961_/X VGND VGND VPWR
+ VPWR _16995_/X sky130_fd_sc_hd__mux4_1
X_33800_ _34312_/CLK _33800_/D VGND VGND VPWR VPWR _33800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18734_ _20294_/A VGND VGND VPWR VPWR _18734_/X sky130_fd_sc_hd__buf_6
XTAP_5270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34780_ _35098_/CLK _34780_/D VGND VGND VPWR VPWR _34780_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31992_ _36200_/CLK _31992_/D VGND VGND VPWR VPWR _31992_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33731_ _33795_/CLK _33731_/D VGND VGND VPWR VPWR _33731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18665_ _35734_/Q _35094_/Q _34454_/Q _33814_/Q _18349_/X _18351_/X VGND VGND VPWR
+ VPWR _18665_/X sky130_fd_sc_hd__mux4_1
X_30943_ _35696_/Q _29157_/X _30953_/S VGND VGND VPWR VPWR _30944_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17616_ _17616_/A _17616_/B _17616_/C _17616_/D VGND VGND VPWR VPWR _17617_/A sky130_fd_sc_hd__or4_1
X_33662_ _34303_/CLK _33662_/D VGND VGND VPWR VPWR _33662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30874_ _35663_/Q _29055_/X _30890_/S VGND VGND VPWR VPWR _30875_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18596_ _20165_/A VGND VGND VPWR VPWR _18596_/X sky130_fd_sc_hd__buf_4
XTAP_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35401_ _35977_/CLK _35401_/D VGND VGND VPWR VPWR _35401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32613_ _36069_/CLK _32613_/D VGND VGND VPWR VPWR _32613_/Q sky130_fd_sc_hd__dfxtp_1
X_17547_ _17547_/A VGND VGND VPWR VPWR _31991_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_233_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33593_ _34298_/CLK _33593_/D VGND VGND VPWR VPWR _33593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_890 _25458_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35332_ _35332_/CLK _35332_/D VGND VGND VPWR VPWR _35332_/Q sky130_fd_sc_hd__dfxtp_1
X_32544_ _35938_/CLK _32544_/D VGND VGND VPWR VPWR _32544_/Q sky130_fd_sc_hd__dfxtp_1
X_17478_ _33526_/Q _33462_/Q _33398_/Q _33334_/Q _17476_/X _17477_/X VGND VGND VPWR
+ VPWR _17478_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19217_ _19149_/X _19215_/X _19216_/X _19152_/X VGND VGND VPWR VPWR _19217_/X sky130_fd_sc_hd__a22o_1
X_35263_ _35581_/CLK _35263_/D VGND VGND VPWR VPWR _35263_/Q sky130_fd_sc_hd__dfxtp_1
X_16429_ _16357_/X _16427_/X _16428_/X _16361_/X VGND VGND VPWR VPWR _16429_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32475_ _35995_/CLK _32475_/D VGND VGND VPWR VPWR _32475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34214_ _34277_/CLK _34214_/D VGND VGND VPWR VPWR _34214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31426_ _23108_/X _35925_/Q _31430_/S VGND VGND VPWR VPWR _31427_/A sky130_fd_sc_hd__mux2_1
X_19148_ _19142_/X _19145_/X _19146_/X _19147_/X VGND VGND VPWR VPWR _19148_/X sky130_fd_sc_hd__a22o_1
X_35194_ _35386_/CLK _35194_/D VGND VGND VPWR VPWR _35194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_955 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34145_ _34145_/CLK _34145_/D VGND VGND VPWR VPWR _34145_/Q sky130_fd_sc_hd__dfxtp_1
X_19079_ _19002_/X _19077_/X _19078_/X _19008_/X VGND VGND VPWR VPWR _19079_/X sky130_fd_sc_hd__a22o_1
X_31357_ _31357_/A VGND VGND VPWR VPWR _35892_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21110_ _35738_/Q _35098_/Q _34458_/Q _33818_/Q _21034_/X _21035_/X VGND VGND VPWR
+ VPWR _21110_/X sky130_fd_sc_hd__mux4_1
X_30308_ _30308_/A VGND VGND VPWR VPWR _35395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22090_ _22443_/A VGND VGND VPWR VPWR _22090_/X sky130_fd_sc_hd__clkbuf_4
X_34076_ _34080_/CLK _34076_/D VGND VGND VPWR VPWR _34076_/Q sky130_fd_sc_hd__dfxtp_1
X_31288_ _31288_/A VGND VGND VPWR VPWR _35859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33027_ _36100_/CLK _33027_/D VGND VGND VPWR VPWR _33027_/Q sky130_fd_sc_hd__dfxtp_1
X_21041_ _22453_/A VGND VGND VPWR VPWR _21041_/X sky130_fd_sc_hd__buf_2
XFILLER_82_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_141_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _35532_/CLK sky130_fd_sc_hd__clkbuf_16
X_30239_ _30239_/A VGND VGND VPWR VPWR _35362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24800_ _22997_/X _32884_/Q _24802_/S VGND VGND VPWR VPWR _24801_/A sky130_fd_sc_hd__mux2_1
X_25780_ _25050_/X _33313_/Q _25780_/S VGND VGND VPWR VPWR _25781_/A sky130_fd_sc_hd__mux2_1
X_34978_ _35042_/CLK _34978_/D VGND VGND VPWR VPWR _34978_/Q sky130_fd_sc_hd__dfxtp_1
X_22992_ _22991_/X _32050_/Q _23001_/S VGND VGND VPWR VPWR _22993_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24731_ _22895_/X _32851_/Q _24739_/S VGND VGND VPWR VPWR _24732_/A sky130_fd_sc_hd__mux2_1
X_33929_ _34817_/CLK _33929_/D VGND VGND VPWR VPWR _33929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21943_ _22430_/A VGND VGND VPWR VPWR _21943_/X sky130_fd_sc_hd__clkbuf_4
X_27450_ _27450_/A VGND VGND VPWR VPWR _34072_/D sky130_fd_sc_hd__clkbuf_1
X_24662_ _24662_/A VGND VGND VPWR VPWR _32819_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21874_ _33264_/Q _36144_/Q _33136_/Q _33072_/Q _21658_/X _21659_/X VGND VGND VPWR
+ VPWR _21874_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26401_ _26401_/A VGND VGND VPWR VPWR _33607_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23613_ _32357_/Q _23199_/X _23625_/S VGND VGND VPWR VPWR _23614_/A sky130_fd_sc_hd__mux2_1
X_20825_ _35538_/Q _35474_/Q _35410_/Q _35346_/Q _20791_/X _20792_/X VGND VGND VPWR
+ VPWR _20825_/X sky130_fd_sc_hd__mux4_1
X_27381_ _34040_/Q _24376_/X _27395_/S VGND VGND VPWR VPWR _27382_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24593_ _24593_/A VGND VGND VPWR VPWR _32786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1022 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26332_ _26332_/A VGND VGND VPWR VPWR _33574_/D sky130_fd_sc_hd__clkbuf_1
X_29120_ input15/X VGND VGND VPWR VPWR _29120_/X sky130_fd_sc_hd__clkbuf_4
X_23544_ _23544_/A VGND VGND VPWR VPWR _32325_/D sky130_fd_sc_hd__clkbuf_1
X_20756_ _35792_/Q _32166_/Q _35664_/Q _35600_/Q _20645_/X _20646_/X VGND VGND VPWR
+ VPWR _20756_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29051_ _31275_/A _30059_/A VGND VGND VPWR VPWR _29247_/S sky130_fd_sc_hd__nor2_8
X_26263_ _25165_/X _33542_/Q _26269_/S VGND VGND VPWR VPWR _26264_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23475_ _23475_/A VGND VGND VPWR VPWR _32292_/D sky130_fd_sc_hd__clkbuf_1
X_20687_ _21754_/A VGND VGND VPWR VPWR _20687_/X sky130_fd_sc_hd__clkbuf_4
X_25214_ _25026_/X _33049_/Q _25230_/S VGND VGND VPWR VPWR _25215_/A sky130_fd_sc_hd__mux2_1
X_28002_ _28002_/A VGND VGND VPWR VPWR _34333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22426_ _33792_/Q _33728_/Q _33664_/Q _33600_/Q _22149_/X _22150_/X VGND VGND VPWR
+ VPWR _22426_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26194_ _25063_/X _33509_/Q _26206_/S VGND VGND VPWR VPWR _26195_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25145_ _25145_/A VGND VGND VPWR VPWR _33023_/D sky130_fd_sc_hd__clkbuf_1
X_22357_ _33534_/Q _33470_/Q _33406_/Q _33342_/Q _22076_/X _22077_/X VGND VGND VPWR
+ VPWR _22357_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_380_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _35760_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_152_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21308_ _22506_/A VGND VGND VPWR VPWR _21308_/X sky130_fd_sc_hd__clkbuf_4
X_29953_ _35227_/Q _29092_/X _29965_/S VGND VGND VPWR VPWR _29954_/A sky130_fd_sc_hd__mux2_1
X_25076_ _25075_/X _33001_/Q _25082_/S VGND VGND VPWR VPWR _25077_/A sky130_fd_sc_hd__mux2_1
X_22288_ _34044_/Q _33980_/Q _33916_/Q _32252_/Q _21973_/X _21974_/X VGND VGND VPWR
+ VPWR _22288_/X sky130_fd_sc_hd__mux4_1
X_28904_ _28904_/A VGND VGND VPWR VPWR _34761_/D sky130_fd_sc_hd__clkbuf_1
X_24027_ _22957_/X _32551_/Q _24035_/S VGND VGND VPWR VPWR _24028_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_132_CLK clkbuf_6_23__f_CLK/X VGND VGND VPWR VPWR _35021_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_215_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21239_ _20957_/X _21235_/X _21238_/X _20961_/X VGND VGND VPWR VPWR _21239_/X sky130_fd_sc_hd__a22o_1
X_29884_ _29884_/A VGND VGND VPWR VPWR _35194_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28835_ _28835_/A VGND VGND VPWR VPWR _34728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28766_ _27002_/X _34696_/Q _28768_/S VGND VGND VPWR VPWR _28767_/A sky130_fd_sc_hd__mux2_1
X_16780_ _32482_/Q _32354_/Q _32034_/Q _36002_/Q _16570_/X _16711_/X VGND VGND VPWR
+ VPWR _16780_/X sky130_fd_sc_hd__mux4_1
X_25978_ _25143_/X _33407_/Q _25978_/S VGND VGND VPWR VPWR _25979_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27717_ _27717_/A VGND VGND VPWR VPWR _34198_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_1459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24929_ _22988_/X _32945_/Q _24937_/S VGND VGND VPWR VPWR _24930_/A sky130_fd_sc_hd__mux2_1
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28697_ _26900_/X _34663_/Q _28705_/S VGND VGND VPWR VPWR _28698_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18450_ _33232_/Q _36112_/Q _33104_/Q _33040_/Q _18320_/X _18321_/X VGND VGND VPWR
+ VPWR _18450_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27648_ _27696_/S VGND VGND VPWR VPWR _27667_/S sky130_fd_sc_hd__buf_4
XFILLER_61_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_131 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_142 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _33780_/Q _33716_/Q _33652_/Q _33588_/Q _17196_/X _17197_/X VGND VGND VPWR
+ VPWR _17401_/X sky130_fd_sc_hd__mux4_1
XANTENNA_153 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18381_ _19307_/A VGND VGND VPWR VPWR _18381_/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_199_CLK clkbuf_6_51__f_CLK/X VGND VGND VPWR VPWR _35968_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_164 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27579_ _34133_/Q _24267_/X _27583_/S VGND VGND VPWR VPWR _27580_/A sky130_fd_sc_hd__mux2_1
XANTENNA_175 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29318_ _23244_/X _34926_/Q _29332_/S VGND VGND VPWR VPWR _29319_/A sky130_fd_sc_hd__mux2_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17332_ _34290_/Q _34226_/Q _34162_/Q _34098_/Q _17089_/X _17090_/X VGND VGND VPWR
+ VPWR _17332_/X sky130_fd_sc_hd__mux4_1
X_30590_ _23333_/X _35529_/Q _30590_/S VGND VGND VPWR VPWR _30591_/A sky130_fd_sc_hd__mux2_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29249_ _29384_/A _31410_/B VGND VGND VPWR VPWR _29382_/S sky130_fd_sc_hd__nand2_8
XFILLER_144_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17263_ _17263_/A _17263_/B _17263_/C _17263_/D VGND VGND VPWR VPWR _17264_/A sky130_fd_sc_hd__or4_4
XFILLER_35_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19002_ _20201_/A VGND VGND VPWR VPWR _19002_/X sky130_fd_sc_hd__clkbuf_4
X_16214_ _32722_/Q _32658_/Q _32594_/Q _36050_/Q _16213_/X _17713_/A VGND VGND VPWR
+ VPWR _16214_/X sky130_fd_sc_hd__mux4_1
X_32260_ _34243_/CLK _32260_/D VGND VGND VPWR VPWR _32260_/Q sky130_fd_sc_hd__dfxtp_1
X_17194_ _17194_/A VGND VGND VPWR VPWR _31981_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16145_ _34000_/Q _33936_/Q _33872_/Q _32144_/Q _16108_/X _16109_/X VGND VGND VPWR
+ VPWR _16145_/X sky130_fd_sc_hd__mux4_1
X_31211_ _35823_/Q input27/X _31223_/S VGND VGND VPWR VPWR _31212_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32191_ _35815_/CLK _32191_/D VGND VGND VPWR VPWR _32191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_371_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _33007_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_192_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16076_ _17932_/A VGND VGND VPWR VPWR _16076_/X sky130_fd_sc_hd__buf_4
X_31142_ _35790_/Q input1/X _31160_/S VGND VGND VPWR VPWR _31143_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19904_ _20257_/A VGND VGND VPWR VPWR _19904_/X sky130_fd_sc_hd__buf_4
XFILLER_142_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31073_ _31073_/A VGND VGND VPWR VPWR _35757_/D sky130_fd_sc_hd__clkbuf_1
X_35950_ _35950_/CLK _35950_/D VGND VGND VPWR VPWR _35950_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_123_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _33940_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_233_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_30__f_CLK clkbuf_5_15_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_30__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30024_ _35261_/Q _29197_/X _30028_/S VGND VGND VPWR VPWR _30025_/A sky130_fd_sc_hd__mux2_1
X_34901_ _36196_/CLK _34901_/D VGND VGND VPWR VPWR _34901_/Q sky130_fd_sc_hd__dfxtp_1
X_19835_ _35575_/Q _35511_/Q _35447_/Q _35383_/Q _19550_/X _19551_/X VGND VGND VPWR
+ VPWR _19835_/X sky130_fd_sc_hd__mux4_1
X_35881_ _35947_/CLK _35881_/D VGND VGND VPWR VPWR _35881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34832_ _35281_/CLK _34832_/D VGND VGND VPWR VPWR _34832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19766_ _19449_/X _19764_/X _19765_/X _19452_/X VGND VGND VPWR VPWR _19766_/X sky130_fd_sc_hd__a22o_1
X_16978_ _33768_/Q _33704_/Q _33640_/Q _33576_/Q _16843_/X _16844_/X VGND VGND VPWR
+ VPWR _16978_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput4 DW[12] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__buf_8
X_18717_ _20095_/A VGND VGND VPWR VPWR _18717_/X sky130_fd_sc_hd__buf_4
X_34763_ _35339_/CLK _34763_/D VGND VGND VPWR VPWR _34763_/Q sky130_fd_sc_hd__dfxtp_1
X_31975_ _35034_/CLK _31975_/D VGND VGND VPWR VPWR _31975_/Q sky130_fd_sc_hd__dfxtp_1
X_19697_ _19454_/X _19695_/X _19696_/X _19459_/X VGND VGND VPWR VPWR _19697_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33714_ _33779_/CLK _33714_/D VGND VGND VPWR VPWR _33714_/Q sky130_fd_sc_hd__dfxtp_1
X_18648_ _18644_/X _18647_/X _18311_/X VGND VGND VPWR VPWR _18680_/A sky130_fd_sc_hd__o21ba_2
X_30926_ _35688_/Q _29132_/X _30932_/S VGND VGND VPWR VPWR _30927_/A sky130_fd_sc_hd__mux2_1
X_34694_ _35334_/CLK _34694_/D VGND VGND VPWR VPWR _34694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33645_ _34283_/CLK _33645_/D VGND VGND VPWR VPWR _33645_/Q sky130_fd_sc_hd__dfxtp_1
X_30857_ _30857_/A VGND VGND VPWR VPWR _35655_/D sky130_fd_sc_hd__clkbuf_1
X_18579_ _32724_/Q _32660_/Q _32596_/Q _36052_/Q _18513_/X _20013_/A VGND VGND VPWR
+ VPWR _18579_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20610_ input75/X input76/X VGND VGND VPWR VPWR _22434_/A sky130_fd_sc_hd__or2b_4
XFILLER_36_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33576_ _34870_/CLK _33576_/D VGND VGND VPWR VPWR _33576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21590_ _22430_/A VGND VGND VPWR VPWR _21590_/X sky130_fd_sc_hd__buf_6
XFILLER_240_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30788_ _30788_/A VGND VGND VPWR VPWR _35622_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35315_ _35315_/CLK _35315_/D VGND VGND VPWR VPWR _35315_/Q sky130_fd_sc_hd__dfxtp_1
X_20541_ _18356_/X _20539_/X _20540_/X _18368_/X VGND VGND VPWR VPWR _20541_/X sky130_fd_sc_hd__a22o_1
X_32527_ _35919_/CLK _32527_/D VGND VGND VPWR VPWR _32527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35246_ _35500_/CLK _35246_/D VGND VGND VPWR VPWR _35246_/Q sky130_fd_sc_hd__dfxtp_1
X_23260_ _23260_/A VGND VGND VPWR VPWR _32204_/D sky130_fd_sc_hd__clkbuf_1
X_32458_ _35147_/CLK _32458_/D VGND VGND VPWR VPWR _32458_/Q sky130_fd_sc_hd__dfxtp_1
X_20472_ _35594_/Q _35530_/Q _35466_/Q _35402_/Q _20256_/X _20257_/X VGND VGND VPWR
+ VPWR _20472_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22211_ _22102_/X _22209_/X _22210_/X _22105_/X VGND VGND VPWR VPWR _22211_/X sky130_fd_sc_hd__a22o_1
X_31409_ _31409_/A VGND VGND VPWR VPWR _35917_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_774 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35177_ _35179_/CLK _35177_/D VGND VGND VPWR VPWR _35177_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_362_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _34288_/CLK sky130_fd_sc_hd__clkbuf_16
X_23191_ _32178_/Q _23127_/X _23206_/S VGND VGND VPWR VPWR _23192_/A sky130_fd_sc_hd__mux2_1
X_32389_ _36037_/CLK _32389_/D VGND VGND VPWR VPWR _32389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34128_ _34259_/CLK _34128_/D VGND VGND VPWR VPWR _34128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22142_ _34551_/Q _32439_/Q _34423_/Q _34359_/Q _21825_/X _21826_/X VGND VGND VPWR
+ VPWR _22142_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34059_ _35273_/CLK _34059_/D VGND VGND VPWR VPWR _34059_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_114_CLK clkbuf_6_20__f_CLK/X VGND VGND VPWR VPWR _36211_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_173_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22073_ _33782_/Q _33718_/Q _33654_/Q _33590_/Q _21796_/X _21797_/X VGND VGND VPWR
+ VPWR _22073_/X sky130_fd_sc_hd__mux4_1
X_26950_ input36/X VGND VGND VPWR VPWR _26950_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21024_ _32728_/Q _32664_/Q _32600_/Q _36056_/Q _20813_/X _20950_/X VGND VGND VPWR
+ VPWR _21024_/X sky130_fd_sc_hd__mux4_1
X_25901_ _25029_/X _33370_/Q _25915_/S VGND VGND VPWR VPWR _25902_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26881_ input11/X VGND VGND VPWR VPWR _26881_/X sky130_fd_sc_hd__buf_4
XFILLER_248_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28620_ _28620_/A VGND VGND VPWR VPWR _34626_/D sky130_fd_sc_hd__clkbuf_1
X_25832_ _25832_/A VGND VGND VPWR VPWR _33337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28551_ _28641_/S VGND VGND VPWR VPWR _28570_/S sky130_fd_sc_hd__buf_4
X_25763_ _25763_/A VGND VGND VPWR VPWR _33304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22975_ _22975_/A VGND VGND VPWR VPWR _32044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27502_ _27502_/A VGND VGND VPWR VPWR _34097_/D sky130_fd_sc_hd__clkbuf_1
X_24714_ _24714_/A VGND VGND VPWR VPWR _32844_/D sky130_fd_sc_hd__clkbuf_1
X_21926_ _35057_/Q _34993_/Q _34929_/Q _34865_/Q _21756_/X _21757_/X VGND VGND VPWR
+ VPWR _21926_/X sky130_fd_sc_hd__mux4_1
X_28482_ _26981_/X _34561_/Q _28498_/S VGND VGND VPWR VPWR _28483_/A sky130_fd_sc_hd__mux2_1
X_25694_ _33273_/Q _24379_/X _25706_/S VGND VGND VPWR VPWR _25695_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27433_ _27433_/A VGND VGND VPWR VPWR _34064_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24645_ _24645_/A VGND VGND VPWR VPWR _32811_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21857_ _35311_/Q _35247_/Q _35183_/Q _32303_/Q _21606_/X _21607_/X VGND VGND VPWR
+ VPWR _21857_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20808_ _20736_/X _20806_/X _20807_/X _20741_/X VGND VGND VPWR VPWR _20808_/X sky130_fd_sc_hd__a22o_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24576_ _24576_/A VGND VGND VPWR VPWR _32780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27364_ _34032_/Q _24351_/X _27374_/S VGND VGND VPWR VPWR _27365_/A sky130_fd_sc_hd__mux2_1
X_21788_ _21749_/X _21786_/X _21787_/X _21752_/X VGND VGND VPWR VPWR _21788_/X sky130_fd_sc_hd__a22o_1
X_29103_ _29103_/A VGND VGND VPWR VPWR _34846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23527_ _23527_/A VGND VGND VPWR VPWR _32317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26315_ _26315_/A VGND VGND VPWR VPWR _33566_/D sky130_fd_sc_hd__clkbuf_1
X_20739_ _33744_/Q _33680_/Q _33616_/Q _33552_/Q _20737_/X _20738_/X VGND VGND VPWR
+ VPWR _20739_/X sky130_fd_sc_hd__mux4_1
X_27295_ _33999_/Q _24249_/X _27311_/S VGND VGND VPWR VPWR _27296_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29034_ _34823_/Q _24422_/X _29038_/S VGND VGND VPWR VPWR _29035_/A sky130_fd_sc_hd__mux2_1
X_26246_ _25140_/X _33534_/Q _26248_/S VGND VGND VPWR VPWR _26247_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23458_ _23458_/A VGND VGND VPWR VPWR _32284_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22409_ _22405_/X _22408_/X _22089_/X _22090_/X VGND VGND VPWR VPWR _22424_/B sky130_fd_sc_hd__o211a_1
XFILLER_167_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26177_ _25038_/X _33501_/Q _26185_/S VGND VGND VPWR VPWR _26178_/A sky130_fd_sc_hd__mux2_1
X_23389_ _23389_/A VGND VGND VPWR VPWR _32253_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_353_CLK clkbuf_6_44__f_CLK/X VGND VGND VPWR VPWR _33013_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25128_ input39/X VGND VGND VPWR VPWR _25128_/X sky130_fd_sc_hd__buf_2
XFILLER_164_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29936_ _35219_/Q _29067_/X _29944_/S VGND VGND VPWR VPWR _29937_/A sky130_fd_sc_hd__mux2_1
X_17950_ _33027_/Q _32963_/Q _32899_/Q _32835_/Q _17695_/X _17696_/X VGND VGND VPWR
+ VPWR _17950_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_105_CLK clkbuf_leaf_80_CLK/A VGND VGND VPWR VPWR _35666_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25059_ _25059_/A VGND VGND VPWR VPWR _32995_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16901_ _16646_/X _16899_/X _16900_/X _16649_/X VGND VGND VPWR VPWR _16901_/X sky130_fd_sc_hd__a22o_1
XFILLER_26_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17881_ _32513_/Q _32385_/Q _32065_/Q _36033_/Q _17629_/X _17770_/X VGND VGND VPWR
+ VPWR _17881_/X sky130_fd_sc_hd__mux4_1
X_29867_ _29867_/A VGND VGND VPWR VPWR _35186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19620_ _19299_/X _19618_/X _19619_/X _19302_/X VGND VGND VPWR VPWR _19620_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16832_ _16828_/X _16831_/X _16794_/X VGND VGND VPWR VPWR _16840_/C sky130_fd_sc_hd__o21ba_1
X_28818_ _28818_/A VGND VGND VPWR VPWR _34720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29798_ _29798_/A VGND VGND VPWR VPWR _35153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19551_ _20257_/A VGND VGND VPWR VPWR _19551_/X sky130_fd_sc_hd__buf_4
X_28749_ _28776_/S VGND VGND VPWR VPWR _28768_/S sky130_fd_sc_hd__clkbuf_8
X_16763_ _16448_/X _16761_/X _16762_/X _16453_/X VGND VGND VPWR VPWR _16763_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18502_ _18387_/X _18500_/X _18501_/X _18397_/X VGND VGND VPWR VPWR _18502_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19482_ _35565_/Q _35501_/Q _35437_/Q _35373_/Q _19197_/X _19198_/X VGND VGND VPWR
+ VPWR _19482_/X sky130_fd_sc_hd__mux4_1
X_31760_ _31760_/A VGND VGND VPWR VPWR _36083_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16694_ _16694_/A VGND VGND VPWR VPWR _31967_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18433_ _18429_/X _18432_/X _18400_/X VGND VGND VPWR VPWR _18434_/D sky130_fd_sc_hd__o21ba_1
X_30711_ _35586_/Q _29213_/X _30725_/S VGND VGND VPWR VPWR _30712_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31691_ _31691_/A VGND VGND VPWR VPWR _36050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33430_ _36228_/CLK _33430_/D VGND VGND VPWR VPWR _33430_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30642_ _30642_/A VGND VGND VPWR VPWR _35553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18364_ _20062_/A VGND VGND VPWR VPWR _20232_/A sky130_fd_sc_hd__buf_12
XFILLER_15_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17315_ _35825_/Q _32202_/Q _35697_/Q _35633_/Q _17313_/X _17314_/X VGND VGND VPWR
+ VPWR _17315_/X sky130_fd_sc_hd__mux4_1
X_33361_ _36232_/CLK _33361_/D VGND VGND VPWR VPWR _33361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18295_ _18295_/A VGND VGND VPWR VPWR _20069_/A sky130_fd_sc_hd__buf_2
X_30573_ _30573_/A VGND VGND VPWR VPWR _35520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35100_ _35933_/CLK _35100_/D VGND VGND VPWR VPWR _35100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32312_ _35319_/CLK _32312_/D VGND VGND VPWR VPWR _32312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17246_ _17242_/X _17245_/X _17136_/X _17137_/X VGND VGND VPWR VPWR _17263_/B sky130_fd_sc_hd__o211a_1
X_36080_ _36080_/CLK _36080_/D VGND VGND VPWR VPWR _36080_/Q sky130_fd_sc_hd__dfxtp_1
X_33292_ _36173_/CLK _33292_/D VGND VGND VPWR VPWR _33292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35031_ _35031_/CLK _35031_/D VGND VGND VPWR VPWR _35031_/Q sky130_fd_sc_hd__dfxtp_1
X_32243_ _34291_/CLK _32243_/D VGND VGND VPWR VPWR _32243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17177_ _17063_/X _17175_/X _17176_/X _17067_/X VGND VGND VPWR VPWR _17177_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_344_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _34229_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16128_ _35279_/Q _35215_/Q _35151_/Q _32271_/Q _16079_/X _16081_/X VGND VGND VPWR
+ VPWR _16128_/X sky130_fd_sc_hd__mux4_1
XFILLER_227_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32174_ _35799_/CLK _32174_/D VGND VGND VPWR VPWR _32174_/Q sky130_fd_sc_hd__dfxtp_1
X_31125_ _31125_/A VGND VGND VPWR VPWR _35782_/D sky130_fd_sc_hd__clkbuf_1
X_16059_ _16059_/A VGND VGND VPWR VPWR _17847_/A sky130_fd_sc_hd__buf_12
XFILLER_142_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31056_ _31056_/A VGND VGND VPWR VPWR _35749_/D sky130_fd_sc_hd__clkbuf_1
X_35933_ _35933_/CLK _35933_/D VGND VGND VPWR VPWR _35933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30007_ _35253_/Q _29172_/X _30007_/S VGND VGND VPWR VPWR _30008_/A sky130_fd_sc_hd__mux2_1
X_19818_ _33783_/Q _33719_/Q _33655_/Q _33591_/Q _19496_/X _19497_/X VGND VGND VPWR
+ VPWR _19818_/X sky130_fd_sc_hd__mux4_1
XFILLER_233_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35864_ _35864_/CLK _35864_/D VGND VGND VPWR VPWR _35864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34815_ _35837_/CLK _34815_/D VGND VGND VPWR VPWR _34815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19749_ _19745_/X _19748_/X _19428_/X VGND VGND VPWR VPWR _19771_/A sky130_fd_sc_hd__o21ba_1
X_35795_ _35797_/CLK _35795_/D VGND VGND VPWR VPWR _35795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22760_ _22508_/X _22758_/X _22759_/X _22511_/X VGND VGND VPWR VPWR _22760_/X sky130_fd_sc_hd__a22o_1
X_34746_ _35771_/CLK _34746_/D VGND VGND VPWR VPWR _34746_/Q sky130_fd_sc_hd__dfxtp_1
X_31958_ _35036_/CLK _31958_/D VGND VGND VPWR VPWR _31958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21711_ _34795_/Q _34731_/Q _34667_/Q _34603_/Q _21535_/X _21536_/X VGND VGND VPWR
+ VPWR _21711_/X sky130_fd_sc_hd__mux4_1
XFILLER_212_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30909_ _35680_/Q _29107_/X _30911_/S VGND VGND VPWR VPWR _30910_/A sky130_fd_sc_hd__mux2_1
X_22691_ _22460_/X _22689_/X _22690_/X _22465_/X VGND VGND VPWR VPWR _22691_/X sky130_fd_sc_hd__a22o_1
X_34677_ _35250_/CLK _34677_/D VGND VGND VPWR VPWR _34677_/Q sky130_fd_sc_hd__dfxtp_1
X_31889_ _31889_/A VGND VGND VPWR VPWR _36144_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24430_ _24430_/A VGND VGND VPWR VPWR _32713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21642_ _34537_/Q _32425_/Q _34409_/Q _34345_/Q _21472_/X _21473_/X VGND VGND VPWR
+ VPWR _21642_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33628_ _34010_/CLK _33628_/D VGND VGND VPWR VPWR _33628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24361_ _32691_/Q _24360_/X _24367_/S VGND VGND VPWR VPWR _24362_/A sky130_fd_sc_hd__mux2_1
X_33559_ _35279_/CLK _33559_/D VGND VGND VPWR VPWR _33559_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_20 _32115_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21573_ _35047_/Q _34983_/Q _34919_/Q _34855_/Q _21403_/X _21404_/X VGND VGND VPWR
+ VPWR _21573_/X sky130_fd_sc_hd__mux4_1
XANTENNA_31 _32116_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26100_ _26100_/A VGND VGND VPWR VPWR _33464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23312_ _23312_/A VGND VGND VPWR VPWR _32221_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_42 _32118_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20524_ _19449_/A _20522_/X _20523_/X _19452_/A VGND VGND VPWR VPWR _20524_/X sky130_fd_sc_hd__a22o_1
XANTENNA_53 _32126_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27080_ _27080_/A VGND VGND VPWR VPWR _33897_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_64 _32126_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24292_ input7/X VGND VGND VPWR VPWR _24292_/X sky130_fd_sc_hd__buf_4
XANTENNA_75 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_86 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26031_ _26142_/S VGND VGND VPWR VPWR _26050_/S sky130_fd_sc_hd__buf_4
XFILLER_165_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_97 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23243_ _23243_/A VGND VGND VPWR VPWR _32198_/D sky130_fd_sc_hd__clkbuf_1
X_35229_ _35293_/CLK _35229_/D VGND VGND VPWR VPWR _35229_/Q sky130_fd_sc_hd__dfxtp_1
X_20455_ _33802_/Q _33738_/Q _33674_/Q _33610_/Q _20202_/X _20203_/X VGND VGND VPWR
+ VPWR _20455_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_335_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _36088_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_181_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23174_ _23174_/A VGND VGND VPWR VPWR _32170_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20386_ _34823_/Q _34759_/Q _34695_/Q _34631_/Q _20294_/X _20295_/X VGND VGND VPWR
+ VPWR _20386_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22125_ _32759_/Q _32695_/Q _32631_/Q _36087_/Q _21872_/X _22009_/X VGND VGND VPWR
+ VPWR _22125_/X sky130_fd_sc_hd__mux4_1
XTAP_6504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27982_ _26841_/X _34324_/Q _27988_/S VGND VGND VPWR VPWR _27983_/A sky130_fd_sc_hd__mux2_1
Xoutput160 _36189_/Q VGND VGND VPWR VPWR D2[15] sky130_fd_sc_hd__buf_2
XTAP_6526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput171 _36199_/Q VGND VGND VPWR VPWR D2[25] sky130_fd_sc_hd__buf_2
XTAP_5803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput182 _36209_/Q VGND VGND VPWR VPWR D2[35] sky130_fd_sc_hd__buf_2
XFILLER_121_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29721_ _35117_/Q _29148_/X _29737_/S VGND VGND VPWR VPWR _29722_/A sky130_fd_sc_hd__mux2_1
XTAP_6548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput193 _36219_/Q VGND VGND VPWR VPWR D2[45] sky130_fd_sc_hd__buf_2
X_26933_ _26933_/A VGND VGND VPWR VPWR _33841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22056_ _22052_/X _22055_/X _21736_/X _21737_/X VGND VGND VPWR VPWR _22071_/B sky130_fd_sc_hd__o211a_1
XTAP_6559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21007_ _20674_/X _21005_/X _21006_/X _20684_/X VGND VGND VPWR VPWR _21007_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29652_ _35085_/Q _29246_/X _29652_/S VGND VGND VPWR VPWR _29653_/A sky130_fd_sc_hd__mux2_1
XTAP_5858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26864_ _26863_/X _33819_/Q _26882_/S VGND VGND VPWR VPWR _26865_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28603_ _28603_/A VGND VGND VPWR VPWR _34618_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25815_ _25815_/A VGND VGND VPWR VPWR _33329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29583_ _29652_/S VGND VGND VPWR VPWR _29602_/S sky130_fd_sc_hd__buf_4
XFILLER_60_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26795_ _33793_/Q _24404_/X _26811_/S VGND VGND VPWR VPWR _26796_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28534_ _28534_/A VGND VGND VPWR VPWR _34585_/D sky130_fd_sc_hd__clkbuf_1
X_25746_ _25746_/A VGND VGND VPWR VPWR _33296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22958_ _22957_/X _32039_/Q _22970_/S VGND VGND VPWR VPWR _22959_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21909_ _32497_/Q _32369_/Q _32049_/Q _36017_/Q _21876_/X _21664_/X VGND VGND VPWR
+ VPWR _21909_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28465_ _26956_/X _34553_/Q _28477_/S VGND VGND VPWR VPWR _28466_/A sky130_fd_sc_hd__mux2_1
X_22889_ input34/X VGND VGND VPWR VPWR _22889_/X sky130_fd_sc_hd__buf_4
X_25677_ _33265_/Q _24354_/X _25685_/S VGND VGND VPWR VPWR _25678_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27416_ _34057_/Q _24428_/X _27416_/S VGND VGND VPWR VPWR _27417_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24628_ _22945_/X _32803_/Q _24644_/S VGND VGND VPWR VPWR _24629_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28396_ _26853_/X _34520_/Q _28414_/S VGND VGND VPWR VPWR _28397_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24559_ _23047_/X _32772_/Q _24569_/S VGND VGND VPWR VPWR _24560_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27347_ _34024_/Q _24326_/X _27353_/S VGND VGND VPWR VPWR _27348_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17100_ _32491_/Q _32363_/Q _32043_/Q _36011_/Q _16923_/X _17064_/X VGND VGND VPWR
+ VPWR _17100_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18080_ _35783_/Q _35143_/Q _34503_/Q _33863_/Q _17846_/X _17847_/X VGND VGND VPWR
+ VPWR _18080_/X sky130_fd_sc_hd__mux4_1
X_27278_ _27278_/A VGND VGND VPWR VPWR _33991_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29017_ _34815_/Q _24397_/X _29017_/S VGND VGND VPWR VPWR _29018_/A sky130_fd_sc_hd__mux2_1
X_17031_ _17027_/X _17030_/X _16783_/X _16784_/X VGND VGND VPWR VPWR _17046_/B sky130_fd_sc_hd__o211a_1
XFILLER_171_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26229_ _26277_/S VGND VGND VPWR VPWR _26248_/S sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_326_CLK clkbuf_6_44__f_CLK/X VGND VGND VPWR VPWR _36021_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18982_ _35551_/Q _35487_/Q _35423_/Q _35359_/Q _18844_/X _18845_/X VGND VGND VPWR
+ VPWR _18982_/X sky130_fd_sc_hd__mux4_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _34562_/Q _32450_/Q _34434_/Q _34370_/Q _17931_/X _17932_/X VGND VGND VPWR
+ VPWR _17933_/X sky130_fd_sc_hd__mux4_1
X_29919_ _29919_/A VGND VGND VPWR VPWR _35211_/D sky130_fd_sc_hd__clkbuf_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32930_ _36067_/CLK _32930_/D VGND VGND VPWR VPWR _32930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17864_ _35072_/Q _35008_/Q _34944_/Q _34880_/Q _17862_/X _17863_/X VGND VGND VPWR
+ VPWR _17864_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19603_ _34033_/Q _33969_/Q _33905_/Q _32241_/Q _19320_/X _19321_/X VGND VGND VPWR
+ VPWR _19603_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16815_ _33507_/Q _33443_/Q _33379_/Q _33315_/Q _16770_/X _16771_/X VGND VGND VPWR
+ VPWR _16815_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32861_ _34146_/CLK _32861_/D VGND VGND VPWR VPWR _32861_/Q sky130_fd_sc_hd__dfxtp_1
X_17795_ _17795_/A VGND VGND VPWR VPWR _17795_/X sky130_fd_sc_hd__buf_6
XFILLER_226_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34600_ _34792_/CLK _34600_/D VGND VGND VPWR VPWR _34600_/Q sky130_fd_sc_hd__dfxtp_1
X_31812_ _31812_/A VGND VGND VPWR VPWR _36108_/D sky130_fd_sc_hd__clkbuf_1
X_19534_ _34287_/Q _34223_/Q _34159_/Q _34095_/Q _19389_/X _19390_/X VGND VGND VPWR
+ VPWR _19534_/X sky130_fd_sc_hd__mux4_1
X_35580_ _35580_/CLK _35580_/D VGND VGND VPWR VPWR _35580_/Q sky130_fd_sc_hd__dfxtp_1
X_16746_ _16702_/X _16744_/X _16745_/X _16708_/X VGND VGND VPWR VPWR _16746_/X sky130_fd_sc_hd__a22o_1
X_32792_ _35995_/CLK _32792_/D VGND VGND VPWR VPWR _32792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34531_ _35938_/CLK _34531_/D VGND VGND VPWR VPWR _34531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31743_ _31743_/A VGND VGND VPWR VPWR _36075_/D sky130_fd_sc_hd__clkbuf_1
X_19465_ _33773_/Q _33709_/Q _33645_/Q _33581_/Q _19143_/X _19144_/X VGND VGND VPWR
+ VPWR _19465_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16677_ _16357_/X _16675_/X _16676_/X _16361_/X VGND VGND VPWR VPWR _16677_/X sky130_fd_sc_hd__a22o_1
XFILLER_59_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18416_ _32463_/Q _32335_/Q _32015_/Q _35983_/Q _18328_/X _20163_/A VGND VGND VPWR
+ VPWR _18416_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34462_ _35743_/CLK _34462_/D VGND VGND VPWR VPWR _34462_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31674_ _36043_/Q input58/X _31678_/S VGND VGND VPWR VPWR _31675_/A sky130_fd_sc_hd__mux2_1
X_19396_ _19392_/X _19395_/X _19075_/X VGND VGND VPWR VPWR _19418_/A sky130_fd_sc_hd__o21ba_1
XFILLER_107_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36201_ _36201_/CLK _36201_/D VGND VGND VPWR VPWR _36201_/Q sky130_fd_sc_hd__dfxtp_2
X_33413_ _34053_/CLK _33413_/D VGND VGND VPWR VPWR _33413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18347_ _35790_/Q _32164_/Q _35662_/Q _35598_/Q _18345_/X _18346_/X VGND VGND VPWR
+ VPWR _18347_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30625_ _35545_/Q _29086_/X _30641_/S VGND VGND VPWR VPWR _30626_/A sky130_fd_sc_hd__mux2_1
XFILLER_226_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34393_ _35293_/CLK _34393_/D VGND VGND VPWR VPWR _34393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36132_ _36132_/CLK _36132_/D VGND VGND VPWR VPWR _36132_/Q sky130_fd_sc_hd__dfxtp_1
X_33344_ _34305_/CLK _33344_/D VGND VGND VPWR VPWR _33344_/Q sky130_fd_sc_hd__dfxtp_1
X_18278_ input77/X VGND VGND VPWR VPWR _18357_/A sky130_fd_sc_hd__buf_6
XFILLER_148_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30556_ _30556_/A VGND VGND VPWR VPWR _35512_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput40 DW[45] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_8
X_17229_ _17154_/X _17227_/X _17228_/X _17159_/X VGND VGND VPWR VPWR _17229_/X sky130_fd_sc_hd__a22o_1
X_36063_ _36063_/CLK _36063_/D VGND VGND VPWR VPWR _36063_/Q sky130_fd_sc_hd__dfxtp_1
X_33275_ _36154_/CLK _33275_/D VGND VGND VPWR VPWR _33275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_317_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _35833_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_200_1244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30487_ _30598_/S VGND VGND VPWR VPWR _30506_/S sky130_fd_sc_hd__buf_4
Xinput51 DW[55] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__buf_8
XFILLER_162_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput62 DW[7] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__buf_8
Xinput73 R2[2] VGND VGND VPWR VPWR input73/X sky130_fd_sc_hd__buf_4
X_35014_ _35079_/CLK _35014_/D VGND VGND VPWR VPWR _35014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput84 RW[1] VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__buf_6
XFILLER_239_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20240_ _34307_/Q _34243_/Q _34179_/Q _34115_/Q _20095_/X _20096_/X VGND VGND VPWR
+ VPWR _20240_/X sky130_fd_sc_hd__mux4_1
X_32226_ _36136_/CLK _32226_/D VGND VGND VPWR VPWR _32226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_928 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20171_ _33793_/Q _33729_/Q _33665_/Q _33601_/Q _19849_/X _19850_/X VGND VGND VPWR
+ VPWR _20171_/X sky130_fd_sc_hd__mux4_1
XFILLER_170_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32157_ _36200_/CLK _32157_/D VGND VGND VPWR VPWR _32157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31108_ _31108_/A VGND VGND VPWR VPWR _35774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32088_ _35040_/CLK _32088_/D VGND VGND VPWR VPWR _32088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35916_ _35981_/CLK _35916_/D VGND VGND VPWR VPWR _35916_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23930_ _23930_/A VGND VGND VPWR VPWR _32505_/D sky130_fd_sc_hd__clkbuf_1
X_31039_ _31039_/A VGND VGND VPWR VPWR _35741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_1097 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23861_ _23861_/A VGND VGND VPWR VPWR _32472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35847_ _35847_/CLK _35847_/D VGND VGND VPWR VPWR _35847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22812_ _22808_/X _22811_/X _22467_/A VGND VGND VPWR VPWR _22813_/D sky130_fd_sc_hd__o21ba_1
X_25600_ input85/X input84/X _27561_/B VGND VGND VPWR VPWR _25601_/A sky130_fd_sc_hd__or3_1
XFILLER_44_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_708 _22532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23792_ _23792_/A VGND VGND VPWR VPWR _32440_/D sky130_fd_sc_hd__clkbuf_1
X_26580_ _26580_/A VGND VGND VPWR VPWR _33691_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_1403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35778_ _35778_/CLK _35778_/D VGND VGND VPWR VPWR _35778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_719 _21749_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22743_ _33225_/Q _32585_/Q _35977_/Q _35913_/Q _20675_/X _20676_/X VGND VGND VPWR
+ VPWR _22743_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25531_ _33197_/Q _24342_/X _25547_/S VGND VGND VPWR VPWR _25532_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34729_ _34794_/CLK _34729_/D VGND VGND VPWR VPWR _34729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25462_ _25462_/A _27561_/B VGND VGND VPWR VPWR _25463_/A sky130_fd_sc_hd__or2_1
X_28250_ _34451_/Q _24261_/X _28258_/S VGND VGND VPWR VPWR _28251_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22674_ _22361_/X _22672_/X _22673_/X _22367_/X VGND VGND VPWR VPWR _22674_/X sky130_fd_sc_hd__a22o_1
XFILLER_201_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24413_ input50/X VGND VGND VPWR VPWR _24413_/X sky130_fd_sc_hd__buf_6
X_27201_ _27201_/A VGND VGND VPWR VPWR _33954_/D sky130_fd_sc_hd__clkbuf_1
X_21625_ _32745_/Q _32681_/Q _32617_/Q _36073_/Q _21519_/X _21303_/X VGND VGND VPWR
+ VPWR _21625_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25393_ _25393_/A VGND VGND VPWR VPWR _33133_/D sky130_fd_sc_hd__clkbuf_1
X_28181_ _28181_/A VGND VGND VPWR VPWR _34418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27132_ _26984_/X _33922_/Q _27146_/S VGND VGND VPWR VPWR _27133_/A sky130_fd_sc_hd__mux2_1
X_24344_ _24344_/A VGND VGND VPWR VPWR _32685_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21556_ _32487_/Q _32359_/Q _32039_/Q _36007_/Q _21523_/X _21311_/X VGND VGND VPWR
+ VPWR _21556_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20507_ _35339_/Q _35275_/Q _35211_/Q _32331_/Q _18388_/X _18390_/X VGND VGND VPWR
+ VPWR _20507_/X sky130_fd_sc_hd__mux4_1
X_27063_ _27063_/A VGND VGND VPWR VPWR _33889_/D sky130_fd_sc_hd__clkbuf_1
X_24275_ _24275_/A VGND VGND VPWR VPWR _32663_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_308_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _35578_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_166_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21487_ _32741_/Q _32677_/Q _32613_/Q _36069_/Q _21166_/X _21303_/X VGND VGND VPWR
+ VPWR _21487_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26014_ _26014_/A VGND VGND VPWR VPWR _33423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23226_ _32193_/Q _23217_/X _23350_/S VGND VGND VPWR VPWR _23227_/A sky130_fd_sc_hd__mux2_1
X_20438_ _20434_/X _20437_/X _20142_/X _20143_/X VGND VGND VPWR VPWR _20453_/B sky130_fd_sc_hd__o211a_1
XFILLER_146_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23157_ input85/X input84/X _26549_/C VGND VGND VPWR VPWR _23158_/A sky130_fd_sc_hd__or3_1
XFILLER_136_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20369_ _34055_/Q _33991_/Q _33927_/Q _32263_/Q _18358_/X _18360_/X VGND VGND VPWR
+ VPWR _20369_/X sky130_fd_sc_hd__mux4_1
XTAP_6301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1107 input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22108_ _34550_/Q _32438_/Q _34422_/Q _34358_/Q _21825_/X _21826_/X VGND VGND VPWR
+ VPWR _22108_/X sky130_fd_sc_hd__mux4_1
XTAP_7079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1118 input53/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23088_ _32142_/Q _23077_/X _23115_/S VGND VGND VPWR VPWR _23089_/A sky130_fd_sc_hd__mux2_1
XTAP_5600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27965_ _27965_/A VGND VGND VPWR VPWR _34316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1129 _31998_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29704_ _35109_/Q _29123_/X _29716_/S VGND VGND VPWR VPWR _29705_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26916_ _27018_/S VGND VGND VPWR VPWR _26944_/S sky130_fd_sc_hd__buf_4
X_22039_ _22039_/A _22039_/B _22039_/C _22039_/D VGND VGND VPWR VPWR _22040_/A sky130_fd_sc_hd__or4_1
XTAP_6389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27896_ _27896_/A VGND VGND VPWR VPWR _34283_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29635_ _29635_/A VGND VGND VPWR VPWR _35076_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26847_ input63/X VGND VGND VPWR VPWR _26847_/X sky130_fd_sc_hd__buf_4
XFILLER_57_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16600_ _32733_/Q _32669_/Q _32605_/Q _36061_/Q _16566_/X _16350_/X VGND VGND VPWR
+ VPWR _16600_/X sky130_fd_sc_hd__mux4_1
XTAP_4987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17580_ _34552_/Q _32440_/Q _34424_/Q _34360_/Q _17578_/X _17579_/X VGND VGND VPWR
+ VPWR _17580_/X sky130_fd_sc_hd__mux4_1
X_29566_ _29566_/A VGND VGND VPWR VPWR _35043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26778_ _33785_/Q _24379_/X _26790_/S VGND VGND VPWR VPWR _26779_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28517_ _28517_/A VGND VGND VPWR VPWR _34577_/D sky130_fd_sc_hd__clkbuf_1
X_16531_ _34011_/Q _33947_/Q _33883_/Q _32155_/Q _16314_/X _16315_/X VGND VGND VPWR
+ VPWR _16531_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25729_ _33290_/Q _24431_/X _25735_/S VGND VGND VPWR VPWR _25730_/A sky130_fd_sc_hd__mux2_1
X_29497_ _23313_/X _35011_/Q _29509_/S VGND VGND VPWR VPWR _29498_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19250_ _34023_/Q _33959_/Q _33895_/Q _32204_/Q _18967_/X _18968_/X VGND VGND VPWR
+ VPWR _19250_/X sky130_fd_sc_hd__mux4_1
X_16462_ _33497_/Q _33433_/Q _33369_/Q _33305_/Q _16417_/X _16418_/X VGND VGND VPWR
+ VPWR _16462_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28448_ _26931_/X _34545_/Q _28456_/S VGND VGND VPWR VPWR _28449_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18201_ _15977_/X _18199_/X _18200_/X _15987_/X VGND VGND VPWR VPWR _18201_/X sky130_fd_sc_hd__a22o_1
XFILLER_204_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19181_ _34277_/Q _34213_/Q _34149_/Q _34085_/Q _19036_/X _19037_/X VGND VGND VPWR
+ VPWR _19181_/X sky130_fd_sc_hd__mux4_1
XPHY_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28379_ _26829_/X _34512_/Q _28393_/S VGND VGND VPWR VPWR _28380_/A sky130_fd_sc_hd__mux2_1
X_16393_ _16349_/X _16391_/X _16392_/X _16355_/X VGND VGND VPWR VPWR _16393_/X sky130_fd_sc_hd__a22o_1
XPHY_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18132_ _32777_/Q _32713_/Q _32649_/Q _36105_/Q _17978_/X _16873_/A VGND VGND VPWR
+ VPWR _18132_/X sky130_fd_sc_hd__mux4_1
X_30410_ _30410_/A VGND VGND VPWR VPWR _35443_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31390_ _35908_/Q input50/X _31400_/S VGND VGND VPWR VPWR _31391_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18063_ _18063_/A _18063_/B _18063_/C _18063_/D VGND VGND VPWR VPWR _18064_/A sky130_fd_sc_hd__or4_4
X_30341_ _30341_/A VGND VGND VPWR VPWR _35410_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1048 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17014_ _17014_/A _17014_/B _17014_/C _17014_/D VGND VGND VPWR VPWR _17015_/A sky130_fd_sc_hd__or4_4
X_33060_ _36130_/CLK _33060_/D VGND VGND VPWR VPWR _33060_/Q sky130_fd_sc_hd__dfxtp_1
X_30272_ _30272_/A VGND VGND VPWR VPWR _35378_/D sky130_fd_sc_hd__clkbuf_1
X_32011_ _36185_/CLK _32011_/D VGND VGND VPWR VPWR _32011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18965_ _18789_/X _18963_/X _18964_/X _18794_/X VGND VGND VPWR VPWR _18965_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17916_ _17761_/X _17914_/X _17915_/X _17767_/X VGND VGND VPWR VPWR _17916_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33962_ _34154_/CLK _33962_/D VGND VGND VPWR VPWR _33962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18896_ _33501_/Q _33437_/Q _33373_/Q _33309_/Q _18717_/X _18718_/X VGND VGND VPWR
+ VPWR _18896_/X sky130_fd_sc_hd__mux4_1
XTAP_6890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32913_ _35985_/CLK _32913_/D VGND VGND VPWR VPWR _32913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35701_ _35828_/CLK _35701_/D VGND VGND VPWR VPWR _35701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17847_ _17847_/A VGND VGND VPWR VPWR _17847_/X sky130_fd_sc_hd__clkbuf_4
X_33893_ _36134_/CLK _33893_/D VGND VGND VPWR VPWR _33893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32844_ _35917_/CLK _32844_/D VGND VGND VPWR VPWR _32844_/Q sky130_fd_sc_hd__dfxtp_1
X_35632_ _35951_/CLK _35632_/D VGND VGND VPWR VPWR _35632_/Q sky130_fd_sc_hd__dfxtp_1
X_17778_ _17700_/X _17776_/X _17777_/X _17703_/X VGND VGND VPWR VPWR _17778_/X sky130_fd_sc_hd__a22o_1
XFILLER_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19517_ _19294_/X _19515_/X _19516_/X _19297_/X VGND VGND VPWR VPWR _19517_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16729_ _34528_/Q _32416_/Q _34400_/Q _34336_/Q _16519_/X _16520_/X VGND VGND VPWR
+ VPWR _16729_/X sky130_fd_sc_hd__mux4_1
X_35563_ _35946_/CLK _35563_/D VGND VGND VPWR VPWR _35563_/Q sky130_fd_sc_hd__dfxtp_1
X_32775_ _36103_/CLK _32775_/D VGND VGND VPWR VPWR _32775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34514_ _35028_/CLK _34514_/D VGND VGND VPWR VPWR _34514_/Q sky130_fd_sc_hd__dfxtp_1
X_19448_ _19443_/X _19446_/X _19447_/X VGND VGND VPWR VPWR _19463_/C sky130_fd_sc_hd__o21ba_1
X_31726_ _36067_/Q input14/X _31742_/S VGND VGND VPWR VPWR _31727_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_1008 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35494_ _35750_/CLK _35494_/D VGND VGND VPWR VPWR _35494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34445_ _35597_/CLK _34445_/D VGND VGND VPWR VPWR _34445_/Q sky130_fd_sc_hd__dfxtp_1
X_31657_ _31657_/A VGND VGND VPWR VPWR _36034_/D sky130_fd_sc_hd__clkbuf_1
X_19379_ _34794_/Q _34730_/Q _34666_/Q _34602_/Q _19235_/X _19236_/X VGND VGND VPWR
+ VPWR _19379_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_94_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _36189_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21410_ _21410_/A _21410_/B _21410_/C _21410_/D VGND VGND VPWR VPWR _21411_/A sky130_fd_sc_hd__or4_4
X_30608_ _35537_/Q _29061_/X _30620_/S VGND VGND VPWR VPWR _30609_/A sky130_fd_sc_hd__mux2_1
X_34376_ _35078_/CLK _34376_/D VGND VGND VPWR VPWR _34376_/Q sky130_fd_sc_hd__dfxtp_1
X_22390_ _22107_/X _22388_/X _22389_/X _22112_/X VGND VGND VPWR VPWR _22390_/X sky130_fd_sc_hd__a22o_1
X_31588_ _31678_/S VGND VGND VPWR VPWR _31607_/S sky130_fd_sc_hd__buf_4
XFILLER_241_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36115_ _36115_/CLK _36115_/D VGND VGND VPWR VPWR _36115_/Q sky130_fd_sc_hd__dfxtp_1
X_33327_ _33520_/CLK _33327_/D VGND VGND VPWR VPWR _33327_/Q sky130_fd_sc_hd__dfxtp_1
X_21341_ _34017_/Q _33953_/Q _33889_/Q _32161_/Q _21267_/X _21268_/X VGND VGND VPWR
+ VPWR _21341_/X sky130_fd_sc_hd__mux4_1
X_30539_ _30539_/A VGND VGND VPWR VPWR _35504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36046_ _36048_/CLK _36046_/D VGND VGND VPWR VPWR _36046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24060_ _24060_/A VGND VGND VPWR VPWR _32566_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21272_ _32735_/Q _32671_/Q _32607_/Q _36063_/Q _21166_/X _20950_/X VGND VGND VPWR
+ VPWR _21272_/X sky130_fd_sc_hd__mux4_1
X_33258_ _36074_/CLK _33258_/D VGND VGND VPWR VPWR _33258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23011_ _23010_/X _32056_/Q _23032_/S VGND VGND VPWR VPWR _23012_/A sky130_fd_sc_hd__mux2_1
X_20223_ _20000_/X _20221_/X _20222_/X _20003_/X VGND VGND VPWR VPWR _20223_/X sky130_fd_sc_hd__a22o_1
X_32209_ _35833_/CLK _32209_/D VGND VGND VPWR VPWR _32209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33189_ _35941_/CLK _33189_/D VGND VGND VPWR VPWR _33189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20154_ _20149_/X _20152_/X _20153_/X VGND VGND VPWR VPWR _20169_/C sky130_fd_sc_hd__o21ba_1
XFILLER_48_1290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27750_ _34214_/Q _24320_/X _27760_/S VGND VGND VPWR VPWR _27751_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24962_ _24962_/A VGND VGND VPWR VPWR _32960_/D sky130_fd_sc_hd__clkbuf_1
X_20085_ _34814_/Q _34750_/Q _34686_/Q _34622_/Q _19941_/X _19942_/X VGND VGND VPWR
+ VPWR _20085_/X sky130_fd_sc_hd__mux4_1
XTAP_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26701_ _26701_/A VGND VGND VPWR VPWR _33748_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23913_ _23913_/A VGND VGND VPWR VPWR _32497_/D sky130_fd_sc_hd__clkbuf_1
X_27681_ _27681_/A VGND VGND VPWR VPWR _34181_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24893_ _22935_/X _32928_/Q _24895_/S VGND VGND VPWR VPWR _24894_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29420_ _29420_/A VGND VGND VPWR VPWR _34974_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26632_ _26632_/A VGND VGND VPWR VPWR _33716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23844_ _23844_/A VGND VGND VPWR VPWR _32464_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_505 _17843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_516 _17970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_527 _18034_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29351_ _23297_/X _34942_/Q _29353_/S VGND VGND VPWR VPWR _29352_/A sky130_fd_sc_hd__mux2_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26563_ _26563_/A VGND VGND VPWR VPWR _33683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23775_ _23775_/A VGND VGND VPWR VPWR _32432_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_538 _20160_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20987_ _33495_/Q _33431_/Q _33367_/Q _33303_/Q _20598_/X _20599_/X VGND VGND VPWR
+ VPWR _20987_/X sky130_fd_sc_hd__mux4_1
XANTENNA_549 _20208_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1080 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28302_ _28371_/S VGND VGND VPWR VPWR _28321_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_81_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25514_ _33189_/Q _24317_/X _25526_/S VGND VGND VPWR VPWR _25515_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22726_ _34313_/Q _34249_/Q _34185_/Q _34121_/Q _20645_/X _20646_/X VGND VGND VPWR
+ VPWR _22726_/X sky130_fd_sc_hd__mux4_1
X_29282_ _23133_/X _34909_/Q _29290_/S VGND VGND VPWR VPWR _29283_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26494_ _26494_/A VGND VGND VPWR VPWR _33651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28233_ _28233_/A VGND VGND VPWR VPWR _34443_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22657_ _35334_/Q _35270_/Q _35206_/Q _32326_/Q _20688_/X _20690_/X VGND VGND VPWR
+ VPWR _22657_/X sky130_fd_sc_hd__mux4_1
X_25445_ _25445_/A VGND VGND VPWR VPWR _33158_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_85_CLK clkbuf_leaf_87_CLK/A VGND VGND VPWR VPWR _36059_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21608_ _35304_/Q _35240_/Q _35176_/Q _32296_/Q _21606_/X _21607_/X VGND VGND VPWR
+ VPWR _21608_/X sky130_fd_sc_hd__mux4_1
XFILLER_167_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28164_ _28164_/A VGND VGND VPWR VPWR _34410_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22588_ _35780_/Q _35140_/Q _34500_/Q _33860_/Q _22446_/X _22447_/X VGND VGND VPWR
+ VPWR _22588_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25376_ _25376_/A VGND VGND VPWR VPWR _33125_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27115_ _26959_/X _33914_/Q _27125_/S VGND VGND VPWR VPWR _27116_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21539_ _21396_/X _21537_/X _21538_/X _21399_/X VGND VGND VPWR VPWR _21539_/X sky130_fd_sc_hd__a22o_1
X_24327_ _32680_/Q _24326_/X _24336_/S VGND VGND VPWR VPWR _24328_/A sky130_fd_sc_hd__mux2_1
X_28095_ _27008_/X _34378_/Q _28101_/S VGND VGND VPWR VPWR _28096_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24258_ input45/X VGND VGND VPWR VPWR _24258_/X sky130_fd_sc_hd__buf_6
X_27046_ _26857_/X _33881_/Q _27062_/S VGND VGND VPWR VPWR _27047_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23209_ _32186_/Q _23148_/X _23235_/S VGND VGND VPWR VPWR _23210_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24189_ _24189_/A VGND VGND VPWR VPWR _32627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28997_ _28997_/A VGND VGND VPWR VPWR _34805_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18750_ _20162_/A VGND VGND VPWR VPWR _18750_/X sky130_fd_sc_hd__buf_4
X_27948_ _34308_/Q _24413_/X _27958_/S VGND VGND VPWR VPWR _27949_/A sky130_fd_sc_hd__mux2_1
XTAP_6175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17701_ _35836_/Q _32214_/Q _35708_/Q _35644_/Q _17666_/X _17667_/X VGND VGND VPWR
+ VPWR _17701_/X sky130_fd_sc_hd__mux4_1
XTAP_5463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18681_ _18681_/A VGND VGND VPWR VPWR _32086_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27879_ _34275_/Q _24311_/X _27895_/S VGND VGND VPWR VPWR _27880_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29618_ _29618_/A VGND VGND VPWR VPWR _35068_/D sky130_fd_sc_hd__clkbuf_1
X_17632_ _17416_/X _17630_/X _17631_/X _17420_/X VGND VGND VPWR VPWR _17632_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30890_ _35671_/Q _29079_/X _30890_/S VGND VGND VPWR VPWR _30891_/A sky130_fd_sc_hd__mux2_1
XTAP_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17563_ _17408_/X _17561_/X _17562_/X _17414_/X VGND VGND VPWR VPWR _17563_/X sky130_fd_sc_hd__a22o_1
X_29549_ _29549_/A VGND VGND VPWR VPWR _35035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19302_ _20165_/A VGND VGND VPWR VPWR _19302_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_32_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16514_ _16293_/X _16512_/X _16513_/X _16296_/X VGND VGND VPWR VPWR _16514_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32560_ _36013_/CLK _32560_/D VGND VGND VPWR VPWR _32560_/Q sky130_fd_sc_hd__dfxtp_1
X_17494_ _17847_/A VGND VGND VPWR VPWR _17494_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_220_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31511_ _31511_/A VGND VGND VPWR VPWR _35965_/D sky130_fd_sc_hd__clkbuf_1
X_19233_ _18946_/X _19231_/X _19232_/X _18949_/X VGND VGND VPWR VPWR _19233_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16445_ _35288_/Q _35224_/Q _35160_/Q _32280_/Q _16300_/X _16301_/X VGND VGND VPWR
+ VPWR _16445_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32491_ _36011_/CLK _32491_/D VGND VGND VPWR VPWR _32491_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_76_CLK clkbuf_leaf_76_CLK/A VGND VGND VPWR VPWR _36112_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_1323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34230_ _36150_/CLK _34230_/D VGND VGND VPWR VPWR _34230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19164_ _18941_/X _19162_/X _19163_/X _18944_/X VGND VGND VPWR VPWR _19164_/X sky130_fd_sc_hd__a22o_1
X_31442_ _31442_/A VGND VGND VPWR VPWR _35932_/D sky130_fd_sc_hd__clkbuf_1
X_16376_ _34518_/Q _32406_/Q _34390_/Q _34326_/Q _16166_/X _16167_/X VGND VGND VPWR
+ VPWR _16376_/X sky130_fd_sc_hd__mux4_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18115_ _18111_/X _18114_/X _17853_/X VGND VGND VPWR VPWR _18123_/C sky130_fd_sc_hd__o21ba_1
XFILLER_129_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34161_ _34227_/CLK _34161_/D VGND VGND VPWR VPWR _34161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31373_ _35900_/Q input41/X _31379_/S VGND VGND VPWR VPWR _31374_/A sky130_fd_sc_hd__mux2_1
X_19095_ _19090_/X _19093_/X _19094_/X VGND VGND VPWR VPWR _19110_/C sky130_fd_sc_hd__o21ba_1
XFILLER_8_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33112_ _34265_/CLK _33112_/D VGND VGND VPWR VPWR _33112_/Q sky130_fd_sc_hd__dfxtp_1
X_30324_ _30324_/A VGND VGND VPWR VPWR _35403_/D sky130_fd_sc_hd__clkbuf_1
X_18046_ _33030_/Q _32966_/Q _32902_/Q _32838_/Q _15980_/X _15983_/X VGND VGND VPWR
+ VPWR _18046_/X sky130_fd_sc_hd__mux4_1
X_34092_ _35315_/CLK _34092_/D VGND VGND VPWR VPWR _34092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33043_ _36115_/CLK _33043_/D VGND VGND VPWR VPWR _33043_/Q sky130_fd_sc_hd__dfxtp_1
X_30255_ _30255_/A VGND VGND VPWR VPWR _35370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30186_ _35338_/Q _29237_/X _30192_/S VGND VGND VPWR VPWR _30187_/A sky130_fd_sc_hd__mux2_1
X_19997_ _33020_/Q _32956_/Q _32892_/Q _32828_/Q _19995_/X _19996_/X VGND VGND VPWR
+ VPWR _19997_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18948_ _33182_/Q _32542_/Q _35934_/Q _35870_/Q _18668_/X _18669_/X VGND VGND VPWR
+ VPWR _18948_/X sky130_fd_sc_hd__mux4_1
X_34994_ _35826_/CLK _34994_/D VGND VGND VPWR VPWR _34994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33945_ _35284_/CLK _33945_/D VGND VGND VPWR VPWR _33945_/Q sky130_fd_sc_hd__dfxtp_1
X_18879_ _33180_/Q _32540_/Q _35932_/Q _35868_/Q _18668_/X _18669_/X VGND VGND VPWR
+ VPWR _18879_/X sky130_fd_sc_hd__mux4_1
XFILLER_227_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20910_ _33749_/Q _33685_/Q _33621_/Q _33557_/Q _20737_/X _20738_/X VGND VGND VPWR
+ VPWR _20910_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33876_ _36232_/CLK _33876_/D VGND VGND VPWR VPWR _33876_/Q sky130_fd_sc_hd__dfxtp_1
X_21890_ _34800_/Q _34736_/Q _34672_/Q _34608_/Q _21888_/X _21889_/X VGND VGND VPWR
+ VPWR _21890_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20841_ _34259_/Q _34195_/Q _34131_/Q _34067_/Q _20605_/X _20607_/X VGND VGND VPWR
+ VPWR _20841_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32827_ _32954_/CLK _32827_/D VGND VGND VPWR VPWR _32827_/Q sky130_fd_sc_hd__dfxtp_1
X_35615_ _35807_/CLK _35615_/D VGND VGND VPWR VPWR _35615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23560_ _23560_/A VGND VGND VPWR VPWR _32333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20772_ _20772_/A _20772_/B _20772_/C _20772_/D VGND VGND VPWR VPWR _20773_/A sky130_fd_sc_hd__or4_4
X_35546_ _35801_/CLK _35546_/D VGND VGND VPWR VPWR _35546_/Q sky130_fd_sc_hd__dfxtp_1
X_32758_ _36087_/CLK _32758_/D VGND VGND VPWR VPWR _32758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22511_ _22511_/A VGND VGND VPWR VPWR _22511_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_126_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31709_ _36059_/Q input5/X _31721_/S VGND VGND VPWR VPWR _31710_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35477_ _35925_/CLK _35477_/D VGND VGND VPWR VPWR _35477_/Q sky130_fd_sc_hd__dfxtp_1
X_23491_ _22972_/X _32300_/Q _23509_/S VGND VGND VPWR VPWR _23492_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_67_CLK clkbuf_leaf_73_CLK/A VGND VGND VPWR VPWR _36116_/CLK sky130_fd_sc_hd__clkbuf_16
X_32689_ _36081_/CLK _32689_/D VGND VGND VPWR VPWR _32689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22442_ _22442_/A VGND VGND VPWR VPWR _22442_/X sky130_fd_sc_hd__buf_4
X_34428_ _34620_/CLK _34428_/D VGND VGND VPWR VPWR _34428_/Q sky130_fd_sc_hd__dfxtp_1
X_25230_ _25050_/X _33057_/Q _25230_/S VGND VGND VPWR VPWR _25231_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25161_ _25161_/A VGND VGND VPWR VPWR _33028_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22373_ _22373_/A VGND VGND VPWR VPWR _22373_/X sky130_fd_sc_hd__clkbuf_4
X_34359_ _35319_/CLK _34359_/D VGND VGND VPWR VPWR _34359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24112_ _24112_/A VGND VGND VPWR VPWR _32590_/D sky130_fd_sc_hd__clkbuf_1
X_21324_ _21246_/X _21320_/X _21323_/X _21249_/X VGND VGND VPWR VPWR _21324_/X sky130_fd_sc_hd__a22o_1
X_25092_ _25091_/X _33006_/Q _25113_/S VGND VGND VPWR VPWR _25093_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28920_ _28920_/A VGND VGND VPWR VPWR _34768_/D sky130_fd_sc_hd__clkbuf_1
X_24043_ _24043_/A VGND VGND VPWR VPWR _32558_/D sky130_fd_sc_hd__clkbuf_1
X_36029_ _36029_/CLK _36029_/D VGND VGND VPWR VPWR _36029_/Q sky130_fd_sc_hd__dfxtp_1
X_21255_ _35294_/Q _35230_/Q _35166_/Q _32286_/Q _21253_/X _21254_/X VGND VGND VPWR
+ VPWR _21255_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20206_ _20206_/A VGND VGND VPWR VPWR _20206_/X sky130_fd_sc_hd__buf_4
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28851_ _26928_/X _34736_/Q _28861_/S VGND VGND VPWR VPWR _28852_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21186_ _21043_/X _21184_/X _21185_/X _21046_/X VGND VGND VPWR VPWR _21186_/X sky130_fd_sc_hd__a22o_1
X_27802_ _34239_/Q _24397_/X _27802_/S VGND VGND VPWR VPWR _27803_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20137_ _33280_/Q _36160_/Q _33152_/Q _33088_/Q _20064_/X _20065_/X VGND VGND VPWR
+ VPWR _20137_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28782_ _26826_/X _34703_/Q _28798_/S VGND VGND VPWR VPWR _28783_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25994_ _25994_/A VGND VGND VPWR VPWR _33414_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27733_ _34206_/Q _24295_/X _27739_/S VGND VGND VPWR VPWR _27734_/A sky130_fd_sc_hd__mux2_1
X_20068_ _20061_/X _20063_/X _20066_/X _20067_/X VGND VGND VPWR VPWR _20068_/X sky130_fd_sc_hd__a22o_1
XTAP_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24945_ _24945_/A VGND VGND VPWR VPWR _32952_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27664_ _27664_/A VGND VGND VPWR VPWR _34173_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24876_ _24987_/S VGND VGND VPWR VPWR _24895_/S sky130_fd_sc_hd__buf_4
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_302 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29403_ _29403_/A VGND VGND VPWR VPWR _34966_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_313 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26615_ _25084_/X _33708_/Q _26633_/S VGND VGND VPWR VPWR _26616_/A sky130_fd_sc_hd__mux2_1
XTAP_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23827_ _23827_/A VGND VGND VPWR VPWR _32457_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_324 _32141_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27595_ _27595_/A VGND VGND VPWR VPWR _34140_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_335 _32141_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_346 _36205_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29334_ _29382_/S VGND VGND VPWR VPWR _29353_/S sky130_fd_sc_hd__buf_4
XANTENNA_357 _36207_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_368 _36207_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26546_ _26546_/A VGND VGND VPWR VPWR _33676_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_379 _36208_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23758_ _23758_/A VGND VGND VPWR VPWR _32424_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22709_ _35848_/Q _32228_/Q _35720_/Q _35656_/Q _20589_/X _20591_/X VGND VGND VPWR
+ VPWR _22709_/X sky130_fd_sc_hd__mux4_1
X_29265_ _23108_/X _34901_/Q _29269_/S VGND VGND VPWR VPWR _29266_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26477_ _26477_/A VGND VGND VPWR VPWR _33643_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23689_ _23689_/A VGND VGND VPWR VPWR _32393_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_58_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _34149_/CLK sky130_fd_sc_hd__clkbuf_16
X_28216_ _26987_/X _34435_/Q _28228_/S VGND VGND VPWR VPWR _28217_/A sky130_fd_sc_hd__mux2_1
X_16230_ _17995_/A VGND VGND VPWR VPWR _16230_/X sky130_fd_sc_hd__buf_4
XFILLER_220_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25428_ _25428_/A VGND VGND VPWR VPWR _33150_/D sky130_fd_sc_hd__clkbuf_1
X_29196_ _29196_/A VGND VGND VPWR VPWR _34876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16161_ _16056_/X _16159_/X _16160_/X _16068_/X VGND VGND VPWR VPWR _16161_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28147_ _26884_/X _34402_/Q _28165_/S VGND VGND VPWR VPWR _28148_/A sky130_fd_sc_hd__mux2_1
X_25359_ _25359_/A VGND VGND VPWR VPWR _33117_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28078_ _28078_/A VGND VGND VPWR VPWR _34369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16092_ _17862_/A VGND VGND VPWR VPWR _16092_/X sky130_fd_sc_hd__buf_4
XFILLER_108_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27029_ _26832_/X _33873_/Q _27041_/S VGND VGND VPWR VPWR _27030_/A sky130_fd_sc_hd__mux2_1
X_19920_ _19848_/X _19918_/X _19919_/X _19853_/X VGND VGND VPWR VPWR _19920_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_1452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30040_ _30040_/A VGND VGND VPWR VPWR _35268_/D sky130_fd_sc_hd__clkbuf_1
X_19851_ _33784_/Q _33720_/Q _33656_/Q _33592_/Q _19849_/X _19850_/X VGND VGND VPWR
+ VPWR _19851_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_929 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18802_ _32730_/Q _32666_/Q _32602_/Q _36058_/Q _18513_/X _18650_/X VGND VGND VPWR
+ VPWR _18802_/X sky130_fd_sc_hd__mux4_1
X_19782_ _19775_/X _19780_/X _19781_/X VGND VGND VPWR VPWR _19816_/A sky130_fd_sc_hd__o21ba_1
XFILLER_228_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16994_ _17855_/A VGND VGND VPWR VPWR _16994_/X sky130_fd_sc_hd__buf_4
XFILLER_7_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18733_ _35800_/Q _32175_/Q _35672_/Q _35608_/Q _18554_/X _18555_/X VGND VGND VPWR
+ VPWR _18733_/X sky130_fd_sc_hd__mux4_1
XFILLER_231_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31991_ _36200_/CLK _31991_/D VGND VGND VPWR VPWR _31991_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33730_ _33795_/CLK _33730_/D VGND VGND VPWR VPWR _33730_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18664_ _35798_/Q _32173_/Q _35670_/Q _35606_/Q _18554_/X _18555_/X VGND VGND VPWR
+ VPWR _18664_/X sky130_fd_sc_hd__mux4_1
X_30942_ _30942_/A VGND VGND VPWR VPWR _35695_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ _17611_/X _17614_/X _17514_/X VGND VGND VPWR VPWR _17616_/D sky130_fd_sc_hd__o21ba_1
XFILLER_97_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33661_ _34044_/CLK _33661_/D VGND VGND VPWR VPWR _33661_/Q sky130_fd_sc_hd__dfxtp_1
X_30873_ _30873_/A VGND VGND VPWR VPWR _35662_/D sky130_fd_sc_hd__clkbuf_1
X_18595_ _33172_/Q _32532_/Q _35924_/Q _35860_/Q _18363_/X _18365_/X VGND VGND VPWR
+ VPWR _18595_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35400_ _35464_/CLK _35400_/D VGND VGND VPWR VPWR _35400_/Q sky130_fd_sc_hd__dfxtp_1
X_32612_ _36067_/CLK _32612_/D VGND VGND VPWR VPWR _32612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17546_ _17546_/A _17546_/B _17546_/C _17546_/D VGND VGND VPWR VPWR _17547_/A sky130_fd_sc_hd__or4_1
X_33592_ _34296_/CLK _33592_/D VGND VGND VPWR VPWR _33592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35331_ _35331_/CLK _35331_/D VGND VGND VPWR VPWR _35331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_880 _25084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_891 _25597_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32543_ _35935_/CLK _32543_/D VGND VGND VPWR VPWR _32543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17477_ _17830_/A VGND VGND VPWR VPWR _17477_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_220_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_49_CLK clkbuf_leaf_50_CLK/A VGND VGND VPWR VPWR _36128_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_177_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_895 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19216_ _34022_/Q _33958_/Q _33894_/Q _32193_/Q _18967_/X _18968_/X VGND VGND VPWR
+ VPWR _19216_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_6_53__f_CLK clkbuf_5_26_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_53__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_220_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35262_ _36105_/CLK _35262_/D VGND VGND VPWR VPWR _35262_/Q sky130_fd_sc_hd__dfxtp_1
X_16428_ _32984_/Q _32920_/Q _32856_/Q _32792_/Q _16283_/X _16284_/X VGND VGND VPWR
+ VPWR _16428_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32474_ _35994_/CLK _32474_/D VGND VGND VPWR VPWR _32474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34213_ _34277_/CLK _34213_/D VGND VGND VPWR VPWR _34213_/Q sky130_fd_sc_hd__dfxtp_1
X_31425_ _31425_/A VGND VGND VPWR VPWR _35924_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19147_ _20206_/A VGND VGND VPWR VPWR _19147_/X sky130_fd_sc_hd__clkbuf_4
X_16359_ _32470_/Q _32342_/Q _32022_/Q _35990_/Q _16217_/X _16358_/X VGND VGND VPWR
+ VPWR _16359_/X sky130_fd_sc_hd__mux4_1
X_35193_ _35320_/CLK _35193_/D VGND VGND VPWR VPWR _35193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34144_ _34777_/CLK _34144_/D VGND VGND VPWR VPWR _34144_/Q sky130_fd_sc_hd__dfxtp_1
X_31356_ _35892_/Q input32/X _31358_/S VGND VGND VPWR VPWR _31357_/A sky130_fd_sc_hd__mux2_1
X_19078_ _33250_/Q _36130_/Q _33122_/Q _33058_/Q _19005_/X _19006_/X VGND VGND VPWR
+ VPWR _19078_/X sky130_fd_sc_hd__mux4_1
XFILLER_246_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18029_ _34565_/Q _32453_/Q _34437_/Q _34373_/Q _17931_/X _17932_/X VGND VGND VPWR
+ VPWR _18029_/X sky130_fd_sc_hd__mux4_1
X_30307_ _35395_/Q _29216_/X _30319_/S VGND VGND VPWR VPWR _30308_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34075_ _34267_/CLK _34075_/D VGND VGND VPWR VPWR _34075_/Q sky130_fd_sc_hd__dfxtp_1
X_31287_ _35859_/Q input56/X _31295_/S VGND VGND VPWR VPWR _31288_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33026_ _33026_/CLK _33026_/D VGND VGND VPWR VPWR _33026_/Q sky130_fd_sc_hd__dfxtp_1
X_21040_ _20893_/X _21038_/X _21039_/X _20896_/X VGND VGND VPWR VPWR _21040_/X sky130_fd_sc_hd__a22o_1
XFILLER_82_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30238_ _35362_/Q _29113_/X _30256_/S VGND VGND VPWR VPWR _30239_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30169_ _30169_/A VGND VGND VPWR VPWR _35329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34977_ _35807_/CLK _34977_/D VGND VGND VPWR VPWR _34977_/Q sky130_fd_sc_hd__dfxtp_1
X_22991_ input30/X VGND VGND VPWR VPWR _22991_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_1290 _17847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24730_ _24730_/A VGND VGND VPWR VPWR _32850_/D sky130_fd_sc_hd__clkbuf_1
X_33928_ _34817_/CLK _33928_/D VGND VGND VPWR VPWR _33928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21942_ _22429_/A VGND VGND VPWR VPWR _21942_/X sky130_fd_sc_hd__buf_4
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21873_ _32752_/Q _32688_/Q _32624_/Q _36080_/Q _21872_/X _21656_/X VGND VGND VPWR
+ VPWR _21873_/X sky130_fd_sc_hd__mux4_1
X_24661_ _22994_/X _32819_/Q _24665_/S VGND VGND VPWR VPWR _24662_/A sky130_fd_sc_hd__mux2_1
X_33859_ _35777_/CLK _33859_/D VGND VGND VPWR VPWR _33859_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26400_ _25168_/X _33607_/Q _26404_/S VGND VGND VPWR VPWR _26401_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20824_ _20644_/X _20822_/X _20823_/X _20654_/X VGND VGND VPWR VPWR _20824_/X sky130_fd_sc_hd__a22o_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23612_ _23612_/A VGND VGND VPWR VPWR _32356_/D sky130_fd_sc_hd__clkbuf_1
X_27380_ _27380_/A VGND VGND VPWR VPWR _34039_/D sky130_fd_sc_hd__clkbuf_1
X_24592_ _22892_/X _32786_/Q _24602_/S VGND VGND VPWR VPWR _24593_/A sky130_fd_sc_hd__mux2_1
X_26331_ _25066_/X _33574_/Q _26341_/S VGND VGND VPWR VPWR _26332_/A sky130_fd_sc_hd__mux2_1
X_23543_ _23050_/X _32325_/Q _23551_/S VGND VGND VPWR VPWR _23544_/A sky130_fd_sc_hd__mux2_1
X_35529_ _35975_/CLK _35529_/D VGND VGND VPWR VPWR _35529_/Q sky130_fd_sc_hd__dfxtp_1
X_20755_ _20751_/X _20754_/X _20640_/X _20642_/X VGND VGND VPWR VPWR _20772_/B sky130_fd_sc_hd__o211a_1
XFILLER_126_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29050_ _29050_/A VGND VGND VPWR VPWR _30059_/A sky130_fd_sc_hd__buf_8
XFILLER_196_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26262_ _26262_/A VGND VGND VPWR VPWR _33541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23474_ _22948_/X _32292_/Q _23488_/S VGND VGND VPWR VPWR _23475_/A sky130_fd_sc_hd__mux2_1
X_20686_ _22369_/A VGND VGND VPWR VPWR _21754_/A sky130_fd_sc_hd__buf_12
XFILLER_17_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28001_ _26869_/X _34333_/Q _28009_/S VGND VGND VPWR VPWR _28002_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22425_ _22425_/A VGND VGND VPWR VPWR _36223_/D sky130_fd_sc_hd__clkbuf_1
X_25213_ _25213_/A VGND VGND VPWR VPWR _33048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26193_ _26193_/A VGND VGND VPWR VPWR _33508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22356_ _22148_/X _22354_/X _22355_/X _22153_/X VGND VGND VPWR VPWR _22356_/X sky130_fd_sc_hd__a22o_1
X_25144_ _25143_/X _33023_/Q _25144_/S VGND VGND VPWR VPWR _25145_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21307_ _33248_/Q _36128_/Q _33120_/Q _33056_/Q _21305_/X _21306_/X VGND VGND VPWR
+ VPWR _21307_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29952_ _29952_/A VGND VGND VPWR VPWR _35226_/D sky130_fd_sc_hd__clkbuf_1
X_25075_ input20/X VGND VGND VPWR VPWR _25075_/X sky130_fd_sc_hd__clkbuf_4
X_22287_ _33532_/Q _33468_/Q _33404_/Q _33340_/Q _22076_/X _22077_/X VGND VGND VPWR
+ VPWR _22287_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28903_ _27005_/X _34761_/Q _28903_/S VGND VGND VPWR VPWR _28904_/A sky130_fd_sc_hd__mux2_1
X_24026_ _24026_/A VGND VGND VPWR VPWR _32550_/D sky130_fd_sc_hd__clkbuf_1
X_21238_ _32990_/Q _32926_/Q _32862_/Q _32798_/Q _21236_/X _21237_/X VGND VGND VPWR
+ VPWR _21238_/X sky130_fd_sc_hd__mux4_1
X_29883_ _35194_/Q _29188_/X _29893_/S VGND VGND VPWR VPWR _29884_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28834_ _26903_/X _34728_/Q _28840_/S VGND VGND VPWR VPWR _28835_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21169_ _20949_/X _21167_/X _21168_/X _20955_/X VGND VGND VPWR VPWR _21169_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28765_ _28765_/A VGND VGND VPWR VPWR _34695_/D sky130_fd_sc_hd__clkbuf_1
X_25977_ _25977_/A VGND VGND VPWR VPWR _33406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27716_ _34198_/Q _24270_/X _27718_/S VGND VGND VPWR VPWR _27717_/A sky130_fd_sc_hd__mux2_1
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24928_ _24928_/A VGND VGND VPWR VPWR _32944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28696_ _28696_/A VGND VGND VPWR VPWR _34662_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27647_ _27647_/A VGND VGND VPWR VPWR _34165_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24859_ _24859_/A VGND VGND VPWR VPWR _32911_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_110 _32129_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_121 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17400_ _17400_/A VGND VGND VPWR VPWR _31987_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ _20062_/A VGND VGND VPWR VPWR _19307_/A sky130_fd_sc_hd__buf_12
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27578_ _27578_/A VGND VGND VPWR VPWR _34132_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_154 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_176 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_187 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29317_ _29317_/A VGND VGND VPWR VPWR _34925_/D sky130_fd_sc_hd__clkbuf_1
X_17331_ _33778_/Q _33714_/Q _33650_/Q _33586_/Q _17196_/X _17197_/X VGND VGND VPWR
+ VPWR _17331_/X sky130_fd_sc_hd__mux4_1
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26529_ _25159_/X _33668_/Q _26539_/S VGND VGND VPWR VPWR _26530_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_198 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29248_ _29248_/A VGND VGND VPWR VPWR _34893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17262_ _17258_/X _17261_/X _17161_/X VGND VGND VPWR VPWR _17263_/D sky130_fd_sc_hd__o21ba_1
XFILLER_81_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19001_ _18997_/X _19000_/X _18722_/X VGND VGND VPWR VPWR _19033_/A sky130_fd_sc_hd__o21ba_1
X_16213_ _17978_/A VGND VGND VPWR VPWR _16213_/X sky130_fd_sc_hd__buf_6
XFILLER_122_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17193_ _17193_/A _17193_/B _17193_/C _17193_/D VGND VGND VPWR VPWR _17194_/A sky130_fd_sc_hd__or4_4
X_29179_ input36/X VGND VGND VPWR VPWR _29179_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_945 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31210_ _31210_/A VGND VGND VPWR VPWR _35822_/D sky130_fd_sc_hd__clkbuf_1
X_16144_ _33488_/Q _33424_/Q _33360_/Q _33296_/Q _15998_/X _15999_/X VGND VGND VPWR
+ VPWR _16144_/X sky130_fd_sc_hd__mux4_1
X_32190_ _35814_/CLK _32190_/D VGND VGND VPWR VPWR _32190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31141_ _31273_/S VGND VGND VPWR VPWR _31160_/S sky130_fd_sc_hd__buf_4
X_16075_ _17931_/A VGND VGND VPWR VPWR _16075_/X sky130_fd_sc_hd__buf_6
XFILLER_143_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19903_ _20256_/A VGND VGND VPWR VPWR _19903_/X sky130_fd_sc_hd__clkbuf_8
X_31072_ _35757_/Q _29148_/X _31088_/S VGND VGND VPWR VPWR _31073_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34900_ _35031_/CLK _34900_/D VGND VGND VPWR VPWR _34900_/Q sky130_fd_sc_hd__dfxtp_1
X_30023_ _30023_/A VGND VGND VPWR VPWR _35260_/D sky130_fd_sc_hd__clkbuf_1
X_19834_ _19647_/X _19832_/X _19833_/X _19650_/X VGND VGND VPWR VPWR _19834_/X sky130_fd_sc_hd__a22o_1
X_35880_ _35947_/CLK _35880_/D VGND VGND VPWR VPWR _35880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34831_ _35282_/CLK _34831_/D VGND VGND VPWR VPWR _34831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16977_ _16977_/A VGND VGND VPWR VPWR _31975_/D sky130_fd_sc_hd__clkbuf_1
X_19765_ _35317_/Q _35253_/Q _35189_/Q _32309_/Q _19659_/X _19660_/X VGND VGND VPWR
+ VPWR _19765_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 DW[13] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__buf_8
XFILLER_77_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18716_ _18436_/X _18714_/X _18715_/X _18441_/X VGND VGND VPWR VPWR _18716_/X sky130_fd_sc_hd__a22o_1
XFILLER_49_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34762_ _35338_/CLK _34762_/D VGND VGND VPWR VPWR _34762_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31974_ _34970_/CLK _31974_/D VGND VGND VPWR VPWR _31974_/Q sky130_fd_sc_hd__dfxtp_1
X_19696_ _35059_/Q _34995_/Q _34931_/Q _34867_/Q _19456_/X _19457_/X VGND VGND VPWR
+ VPWR _19696_/X sky130_fd_sc_hd__mux4_1
XFILLER_188_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18647_ _18443_/X _18645_/X _18646_/X _18446_/X VGND VGND VPWR VPWR _18647_/X sky130_fd_sc_hd__a22o_1
X_30925_ _30925_/A VGND VGND VPWR VPWR _35687_/D sky130_fd_sc_hd__clkbuf_1
X_33713_ _33779_/CLK _33713_/D VGND VGND VPWR VPWR _33713_/Q sky130_fd_sc_hd__dfxtp_1
X_34693_ _35333_/CLK _34693_/D VGND VGND VPWR VPWR _34693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18578_ _18574_/X _18577_/X _18311_/X VGND VGND VPWR VPWR _18608_/A sky130_fd_sc_hd__o21ba_2
X_30856_ _23327_/X _35655_/Q _30860_/S VGND VGND VPWR VPWR _30857_/A sky130_fd_sc_hd__mux2_1
X_33644_ _34283_/CLK _33644_/D VGND VGND VPWR VPWR _33644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17529_ _33015_/Q _32951_/Q _32887_/Q _32823_/Q _17342_/X _17343_/X VGND VGND VPWR
+ VPWR _17529_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33575_ _34278_/CLK _33575_/D VGND VGND VPWR VPWR _33575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30787_ _23217_/X _35622_/Q _30797_/S VGND VGND VPWR VPWR _30788_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20540_ _35084_/Q _35020_/Q _34956_/Q _34892_/Q _18379_/X _18381_/X VGND VGND VPWR
+ VPWR _20540_/X sky130_fd_sc_hd__mux4_1
XFILLER_221_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32526_ _34317_/CLK _32526_/D VGND VGND VPWR VPWR _32526_/Q sky130_fd_sc_hd__dfxtp_1
X_35314_ _35700_/CLK _35314_/D VGND VGND VPWR VPWR _35314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32457_ _35848_/CLK _32457_/D VGND VGND VPWR VPWR _32457_/Q sky130_fd_sc_hd__dfxtp_1
X_20471_ _18277_/X _20469_/X _20470_/X _18287_/X VGND VGND VPWR VPWR _20471_/X sky130_fd_sc_hd__a22o_1
X_35245_ _35500_/CLK _35245_/D VGND VGND VPWR VPWR _35245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22210_ _35321_/Q _35257_/Q _35193_/Q _32313_/Q _21959_/X _21960_/X VGND VGND VPWR
+ VPWR _22210_/X sky130_fd_sc_hd__mux4_1
X_31408_ _35917_/Q input60/X _31408_/S VGND VGND VPWR VPWR _31409_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35176_ _35179_/CLK _35176_/D VGND VGND VPWR VPWR _35176_/Q sky130_fd_sc_hd__dfxtp_1
X_23190_ _23190_/A VGND VGND VPWR VPWR _32177_/D sky130_fd_sc_hd__clkbuf_1
X_32388_ _32901_/CLK _32388_/D VGND VGND VPWR VPWR _32388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_786 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34127_ _35021_/CLK _34127_/D VGND VGND VPWR VPWR _34127_/Q sky130_fd_sc_hd__dfxtp_1
X_22141_ _22102_/X _22139_/X _22140_/X _22105_/X VGND VGND VPWR VPWR _22141_/X sky130_fd_sc_hd__a22o_1
X_31339_ _31408_/S VGND VGND VPWR VPWR _31358_/S sky130_fd_sc_hd__buf_6
XFILLER_156_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34058_ _35273_/CLK _34058_/D VGND VGND VPWR VPWR _34058_/Q sky130_fd_sc_hd__dfxtp_1
X_22072_ _22072_/A VGND VGND VPWR VPWR _36213_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21023_ _21016_/X _21021_/X _21022_/X VGND VGND VPWR VPWR _21057_/A sky130_fd_sc_hd__o21ba_1
X_25900_ _25900_/A VGND VGND VPWR VPWR _33369_/D sky130_fd_sc_hd__clkbuf_1
X_33009_ _33009_/CLK _33009_/D VGND VGND VPWR VPWR _33009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26880_ _26880_/A VGND VGND VPWR VPWR _33824_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25831_ _25125_/X _33337_/Q _25843_/S VGND VGND VPWR VPWR _25832_/A sky130_fd_sc_hd__mux2_1
XFILLER_247_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28550_ _28550_/A VGND VGND VPWR VPWR _34593_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25762_ _25022_/X _33304_/Q _25780_/S VGND VGND VPWR VPWR _25763_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22974_ _22972_/X _32044_/Q _23001_/S VGND VGND VPWR VPWR _22975_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27501_ _26931_/X _34097_/Q _27509_/S VGND VGND VPWR VPWR _27502_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24713_ _23071_/X _32844_/Q _24715_/S VGND VGND VPWR VPWR _24714_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28481_ _28481_/A VGND VGND VPWR VPWR _34560_/D sky130_fd_sc_hd__clkbuf_1
X_21925_ _34545_/Q _32433_/Q _34417_/Q _34353_/Q _21825_/X _21826_/X VGND VGND VPWR
+ VPWR _21925_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25693_ _25693_/A VGND VGND VPWR VPWR _33272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27432_ _26829_/X _34064_/Q _27446_/S VGND VGND VPWR VPWR _27433_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24644_ _22969_/X _32811_/Q _24644_/S VGND VGND VPWR VPWR _24645_/A sky130_fd_sc_hd__mux2_1
X_21856_ _34799_/Q _34735_/Q _34671_/Q _34607_/Q _21535_/X _21536_/X VGND VGND VPWR
+ VPWR _21856_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20807_ _34258_/Q _34194_/Q _34130_/Q _34066_/Q _20605_/X _20607_/X VGND VGND VPWR
+ VPWR _20807_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27363_ _27363_/A VGND VGND VPWR VPWR _34031_/D sky130_fd_sc_hd__clkbuf_1
X_24575_ _23071_/X _32780_/Q _24577_/S VGND VGND VPWR VPWR _24576_/A sky130_fd_sc_hd__mux2_1
X_21787_ _35309_/Q _35245_/Q _35181_/Q _32301_/Q _21606_/X _21607_/X VGND VGND VPWR
+ VPWR _21787_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29102_ _34846_/Q _29101_/X _29111_/S VGND VGND VPWR VPWR _29103_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26314_ _25041_/X _33566_/Q _26320_/S VGND VGND VPWR VPWR _26315_/A sky130_fd_sc_hd__mux2_1
X_23526_ _23025_/X _32317_/Q _23530_/S VGND VGND VPWR VPWR _23527_/A sky130_fd_sc_hd__mux2_1
X_27294_ _27294_/A VGND VGND VPWR VPWR _33998_/D sky130_fd_sc_hd__clkbuf_1
X_20738_ _22503_/A VGND VGND VPWR VPWR _20738_/X sky130_fd_sc_hd__buf_6
XFILLER_243_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29033_ _29033_/A VGND VGND VPWR VPWR _34822_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26245_ _26245_/A VGND VGND VPWR VPWR _33533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20669_ _20656_/X _20661_/X _20666_/X _20668_/X VGND VGND VPWR VPWR _20669_/X sky130_fd_sc_hd__a22o_1
X_23457_ _22923_/X _32284_/Q _23467_/S VGND VGND VPWR VPWR _23458_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22408_ _22369_/X _22406_/X _22407_/X _22373_/X VGND VGND VPWR VPWR _22408_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26176_ _26176_/A VGND VGND VPWR VPWR _33500_/D sky130_fd_sc_hd__clkbuf_1
X_23388_ _32253_/Q _23294_/X _23392_/S VGND VGND VPWR VPWR _23389_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25127_ _25127_/A VGND VGND VPWR VPWR _33017_/D sky130_fd_sc_hd__clkbuf_1
X_22339_ _35773_/Q _35133_/Q _34493_/Q _33853_/Q _22093_/X _22094_/X VGND VGND VPWR
+ VPWR _22339_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29935_ _29935_/A VGND VGND VPWR VPWR _35218_/D sky130_fd_sc_hd__clkbuf_1
X_25058_ _25057_/X _32995_/Q _25082_/S VGND VGND VPWR VPWR _25059_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16900_ _33189_/Q _32549_/Q _35941_/Q _35877_/Q _16721_/X _16722_/X VGND VGND VPWR
+ VPWR _16900_/X sky130_fd_sc_hd__mux4_1
X_24009_ _24009_/A VGND VGND VPWR VPWR _32542_/D sky130_fd_sc_hd__clkbuf_1
X_17880_ _17761_/X _17878_/X _17879_/X _17767_/X VGND VGND VPWR VPWR _17880_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29866_ _35186_/Q _29163_/X _29872_/S VGND VGND VPWR VPWR _29867_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16831_ _16646_/X _16829_/X _16830_/X _16649_/X VGND VGND VPWR VPWR _16831_/X sky130_fd_sc_hd__a22o_1
X_28817_ _26878_/X _34720_/Q _28819_/S VGND VGND VPWR VPWR _28818_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29797_ _35153_/Q _29061_/X _29809_/S VGND VGND VPWR VPWR _29798_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19550_ _20256_/A VGND VGND VPWR VPWR _19550_/X sky130_fd_sc_hd__buf_6
XFILLER_232_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28748_ _28748_/A VGND VGND VPWR VPWR _34687_/D sky130_fd_sc_hd__clkbuf_1
X_16762_ _35041_/Q _34977_/Q _34913_/Q _34849_/Q _16450_/X _16451_/X VGND VGND VPWR
+ VPWR _16762_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_1171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18501_ _35025_/Q _34961_/Q _34897_/Q _34833_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _18501_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19481_ _19294_/X _19479_/X _19480_/X _19297_/X VGND VGND VPWR VPWR _19481_/X sky130_fd_sc_hd__a22o_1
X_16693_ _16693_/A _16693_/B _16693_/C _16693_/D VGND VGND VPWR VPWR _16694_/A sky130_fd_sc_hd__or4_1
X_28679_ _28679_/A VGND VGND VPWR VPWR _34654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_784 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18432_ _18387_/X _18430_/X _18431_/X _18397_/X VGND VGND VPWR VPWR _18432_/X sky130_fd_sc_hd__a22o_1
X_30710_ _30710_/A VGND VGND VPWR VPWR _35585_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31690_ _36050_/Q input45/X _31700_/S VGND VGND VPWR VPWR _31691_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _20231_/A VGND VGND VPWR VPWR _18363_/X sky130_fd_sc_hd__buf_6
X_30641_ _35553_/Q _29110_/X _30641_/S VGND VGND VPWR VPWR _30642_/A sky130_fd_sc_hd__mux2_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _17796_/A VGND VGND VPWR VPWR _17314_/X sky130_fd_sc_hd__buf_4
XFILLER_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33360_ _33940_/CLK _33360_/D VGND VGND VPWR VPWR _33360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18294_ input79/X input80/X VGND VGND VPWR VPWR _18295_/A sky130_fd_sc_hd__and2_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30572_ _23303_/X _35520_/Q _30590_/S VGND VGND VPWR VPWR _30573_/A sky130_fd_sc_hd__mux2_1
X_32311_ _35318_/CLK _32311_/D VGND VGND VPWR VPWR _32311_/Q sky130_fd_sc_hd__dfxtp_1
X_17245_ _17063_/X _17243_/X _17244_/X _17067_/X VGND VGND VPWR VPWR _17245_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33291_ _36107_/CLK _33291_/D VGND VGND VPWR VPWR _33291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35030_ _35730_/CLK _35030_/D VGND VGND VPWR VPWR _35030_/Q sky130_fd_sc_hd__dfxtp_1
X_32242_ _34222_/CLK _32242_/D VGND VGND VPWR VPWR _32242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17176_ _33005_/Q _32941_/Q _32877_/Q _32813_/Q _16989_/X _16990_/X VGND VGND VPWR
+ VPWR _17176_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16127_ _34767_/Q _34703_/Q _34639_/Q _34575_/Q _16075_/X _16076_/X VGND VGND VPWR
+ VPWR _16127_/X sky130_fd_sc_hd__mux4_1
X_32173_ _35799_/CLK _32173_/D VGND VGND VPWR VPWR _32173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31124_ _35782_/Q _29225_/X _31130_/S VGND VGND VPWR VPWR _31125_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16058_ _17846_/A VGND VGND VPWR VPWR _16058_/X sky130_fd_sc_hd__buf_8
XFILLER_115_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31055_ _35749_/Q _29123_/X _31067_/S VGND VGND VPWR VPWR _31056_/A sky130_fd_sc_hd__mux2_1
X_35932_ _35932_/CLK _35932_/D VGND VGND VPWR VPWR _35932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30006_ _30006_/A VGND VGND VPWR VPWR _35252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19817_ _19817_/A VGND VGND VPWR VPWR _32118_/D sky130_fd_sc_hd__buf_2
X_35863_ _35863_/CLK _35863_/D VGND VGND VPWR VPWR _35863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34814_ _36031_/CLK _34814_/D VGND VGND VPWR VPWR _34814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19748_ _19502_/X _19746_/X _19747_/X _19505_/X VGND VGND VPWR VPWR _19748_/X sky130_fd_sc_hd__a22o_1
X_35794_ _35922_/CLK _35794_/D VGND VGND VPWR VPWR _35794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34745_ _34745_/CLK _34745_/D VGND VGND VPWR VPWR _34745_/Q sky130_fd_sc_hd__dfxtp_1
X_31957_ _35036_/CLK _31957_/D VGND VGND VPWR VPWR _31957_/Q sky130_fd_sc_hd__dfxtp_1
X_19679_ _33267_/Q _36147_/Q _33139_/Q _33075_/Q _19358_/X _19359_/X VGND VGND VPWR
+ VPWR _19679_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_280_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _34171_/CLK sky130_fd_sc_hd__clkbuf_16
X_21710_ _21706_/X _21709_/X _21394_/X VGND VGND VPWR VPWR _21718_/C sky130_fd_sc_hd__o21ba_1
X_22690_ _35079_/Q _35015_/Q _34951_/Q _34887_/Q _22462_/X _22463_/X VGND VGND VPWR
+ VPWR _22690_/X sky130_fd_sc_hd__mux4_1
X_30908_ _30908_/A VGND VGND VPWR VPWR _35679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31888_ _23250_/X _36144_/Q _31898_/S VGND VGND VPWR VPWR _31889_/A sky130_fd_sc_hd__mux2_1
X_34676_ _34739_/CLK _34676_/D VGND VGND VPWR VPWR _34676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21641_ _21396_/X _21639_/X _21640_/X _21399_/X VGND VGND VPWR VPWR _21641_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30839_ _23300_/X _35647_/Q _30839_/S VGND VGND VPWR VPWR _30840_/A sky130_fd_sc_hd__mux2_1
X_33627_ _34266_/CLK _33627_/D VGND VGND VPWR VPWR _33627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21572_ _34535_/Q _32423_/Q _34407_/Q _34343_/Q _21472_/X _21473_/X VGND VGND VPWR
+ VPWR _21572_/X sky130_fd_sc_hd__mux4_1
X_24360_ input31/X VGND VGND VPWR VPWR _24360_/X sky130_fd_sc_hd__buf_4
X_33558_ _33685_/CLK _33558_/D VGND VGND VPWR VPWR _33558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_10 _32114_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_21 _32115_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_32 _32117_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23311_ _32221_/Q _23310_/X _23334_/S VGND VGND VPWR VPWR _23312_/A sky130_fd_sc_hd__mux2_1
X_20523_ _33292_/Q _36172_/Q _33164_/Q _33100_/Q _18328_/X _19457_/A VGND VGND VPWR
+ VPWR _20523_/X sky130_fd_sc_hd__mux4_1
XANTENNA_43 _32118_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 _32126_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32509_ _36029_/CLK _32509_/D VGND VGND VPWR VPWR _32509_/Q sky130_fd_sc_hd__dfxtp_1
X_24291_ _24291_/A VGND VGND VPWR VPWR _32668_/D sky130_fd_sc_hd__clkbuf_1
X_33489_ _36237_/CLK _33489_/D VGND VGND VPWR VPWR _33489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_65 _32126_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26030_ _26030_/A VGND VGND VPWR VPWR _33431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_87 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20454_ _20454_/A VGND VGND VPWR VPWR _32137_/D sky130_fd_sc_hd__buf_4
XANTENNA_98 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23242_ _32198_/Q _23241_/X _23268_/S VGND VGND VPWR VPWR _23243_/A sky130_fd_sc_hd__mux2_1
X_35228_ _35292_/CLK _35228_/D VGND VGND VPWR VPWR _35228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23173_ _32170_/Q _23105_/X _23182_/S VGND VGND VPWR VPWR _23174_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20385_ _20381_/X _20384_/X _20153_/X VGND VGND VPWR VPWR _20393_/C sky130_fd_sc_hd__o21ba_1
X_35159_ _36202_/CLK _35159_/D VGND VGND VPWR VPWR _35159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22124_ _22120_/X _22123_/X _22081_/X VGND VGND VPWR VPWR _22146_/A sky130_fd_sc_hd__o21ba_1
XTAP_6505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27981_ _27981_/A VGND VGND VPWR VPWR _34323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput150 _31956_/Q VGND VGND VPWR VPWR D1[6] sky130_fd_sc_hd__buf_2
XTAP_6516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput161 _36190_/Q VGND VGND VPWR VPWR D2[16] sky130_fd_sc_hd__buf_2
XFILLER_115_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput172 _36200_/Q VGND VGND VPWR VPWR D2[26] sky130_fd_sc_hd__buf_2
X_29720_ _29720_/A VGND VGND VPWR VPWR _35116_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput183 _36210_/Q VGND VGND VPWR VPWR D2[36] sky130_fd_sc_hd__buf_2
X_26932_ _26931_/X _33841_/Q _26944_/S VGND VGND VPWR VPWR _26933_/A sky130_fd_sc_hd__mux2_1
X_22055_ _22016_/X _22053_/X _22054_/X _22020_/X VGND VGND VPWR VPWR _22055_/X sky130_fd_sc_hd__a22o_1
XTAP_6549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput194 _36220_/Q VGND VGND VPWR VPWR D2[46] sky130_fd_sc_hd__buf_2
XTAP_5815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21006_ _35287_/Q _35223_/Q _35159_/Q _32279_/Q _20900_/X _20901_/X VGND VGND VPWR
+ VPWR _21006_/X sky130_fd_sc_hd__mux4_1
X_29651_ _29651_/A VGND VGND VPWR VPWR _35084_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26863_ input5/X VGND VGND VPWR VPWR _26863_/X sky130_fd_sc_hd__buf_4
XFILLER_248_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28602_ _26959_/X _34618_/Q _28612_/S VGND VGND VPWR VPWR _28603_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25814_ _25100_/X _33329_/Q _25822_/S VGND VGND VPWR VPWR _25815_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29582_ _29582_/A VGND VGND VPWR VPWR _35051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26794_ _26794_/A VGND VGND VPWR VPWR _33792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28533_ _26857_/X _34585_/Q _28549_/S VGND VGND VPWR VPWR _28534_/A sky130_fd_sc_hd__mux2_1
X_25745_ _24998_/X _33296_/Q _25759_/S VGND VGND VPWR VPWR _25746_/A sky130_fd_sc_hd__mux2_1
X_22957_ input18/X VGND VGND VPWR VPWR _22957_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_55_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_271_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _33789_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_244_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28464_ _28464_/A VGND VGND VPWR VPWR _34552_/D sky130_fd_sc_hd__clkbuf_1
X_21908_ _21655_/X _21906_/X _21907_/X _21661_/X VGND VGND VPWR VPWR _21908_/X sky130_fd_sc_hd__a22o_1
XFILLER_189_929 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25676_ _25676_/A VGND VGND VPWR VPWR _33264_/D sky130_fd_sc_hd__clkbuf_1
X_22888_ _22888_/A VGND VGND VPWR VPWR _32016_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27415_ _27415_/A VGND VGND VPWR VPWR _34056_/D sky130_fd_sc_hd__clkbuf_1
X_24627_ _24627_/A VGND VGND VPWR VPWR _32802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21839_ _21835_/X _21838_/X _21728_/X VGND VGND VPWR VPWR _21863_/A sky130_fd_sc_hd__o21ba_1
X_28395_ _28506_/S VGND VGND VPWR VPWR _28414_/S sky130_fd_sc_hd__buf_4
XFILLER_54_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27346_ _27346_/A VGND VGND VPWR VPWR _34023_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24558_ _24558_/A VGND VGND VPWR VPWR _32771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23509_ _23000_/X _32309_/Q _23509_/S VGND VGND VPWR VPWR _23510_/A sky130_fd_sc_hd__mux2_1
X_27277_ _26999_/X _33991_/Q _27281_/S VGND VGND VPWR VPWR _27278_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24489_ _24489_/A VGND VGND VPWR VPWR _32738_/D sky130_fd_sc_hd__clkbuf_1
X_29016_ _29016_/A VGND VGND VPWR VPWR _34814_/D sky130_fd_sc_hd__clkbuf_1
X_17030_ _16710_/X _17028_/X _17029_/X _16714_/X VGND VGND VPWR VPWR _17030_/X sky130_fd_sc_hd__a22o_1
X_26228_ _26228_/A VGND VGND VPWR VPWR _33525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26159_ _26159_/A VGND VGND VPWR VPWR _33492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18981_ _18941_/X _18979_/X _18980_/X _18944_/X VGND VGND VPWR VPWR _18981_/X sky130_fd_sc_hd__a22o_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29918_ _35211_/Q _29240_/X _29922_/S VGND VGND VPWR VPWR _29919_/A sky130_fd_sc_hd__mux2_1
X_17932_ _17932_/A VGND VGND VPWR VPWR _17932_/X sky130_fd_sc_hd__buf_4
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17863_ _17863_/A VGND VGND VPWR VPWR _17863_/X sky130_fd_sc_hd__buf_4
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29849_ _35178_/Q _29138_/X _29851_/S VGND VGND VPWR VPWR _29850_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19602_ _33521_/Q _33457_/Q _33393_/Q _33329_/Q _19423_/X _19424_/X VGND VGND VPWR
+ VPWR _19602_/X sky130_fd_sc_hd__mux4_1
XFILLER_213_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16814_ _16489_/X _16812_/X _16813_/X _16494_/X VGND VGND VPWR VPWR _16814_/X sky130_fd_sc_hd__a22o_1
X_17794_ _33791_/Q _33727_/Q _33663_/Q _33599_/Q _17549_/X _17550_/X VGND VGND VPWR
+ VPWR _17794_/X sky130_fd_sc_hd__mux4_1
X_32860_ _32860_/CLK _32860_/D VGND VGND VPWR VPWR _32860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31811_ _36108_/Q input59/X _31813_/S VGND VGND VPWR VPWR _31812_/A sky130_fd_sc_hd__mux2_1
X_19533_ _33775_/Q _33711_/Q _33647_/Q _33583_/Q _19496_/X _19497_/X VGND VGND VPWR
+ VPWR _19533_/X sky130_fd_sc_hd__mux4_1
X_16745_ _33249_/Q _36129_/Q _33121_/Q _33057_/Q _16705_/X _16706_/X VGND VGND VPWR
+ VPWR _16745_/X sky130_fd_sc_hd__mux4_1
X_32791_ _35991_/CLK _32791_/D VGND VGND VPWR VPWR _32791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_262_CLK clkbuf_6_57__f_CLK/X VGND VGND VPWR VPWR _36098_/CLK sky130_fd_sc_hd__clkbuf_16
X_19464_ _19464_/A VGND VGND VPWR VPWR _32108_/D sky130_fd_sc_hd__buf_2
X_34530_ _35298_/CLK _34530_/D VGND VGND VPWR VPWR _34530_/Q sky130_fd_sc_hd__dfxtp_1
X_31742_ _36075_/Q input22/X _31742_/S VGND VGND VPWR VPWR _31743_/A sky130_fd_sc_hd__mux2_1
X_16676_ _32991_/Q _32927_/Q _32863_/Q _32799_/Q _16636_/X _16637_/X VGND VGND VPWR
+ VPWR _16676_/X sky130_fd_sc_hd__mux4_1
XFILLER_234_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18415_ _18314_/X _18413_/X _18414_/X _18323_/X VGND VGND VPWR VPWR _18415_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31673_ _31673_/A VGND VGND VPWR VPWR _36042_/D sky130_fd_sc_hd__clkbuf_1
X_34461_ _35933_/CLK _34461_/D VGND VGND VPWR VPWR _34461_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19395_ _19149_/X _19393_/X _19394_/X _19152_/X VGND VGND VPWR VPWR _19395_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36200_ _36200_/CLK _36200_/D VGND VGND VPWR VPWR _36200_/Q sky130_fd_sc_hd__dfxtp_2
X_33412_ _33545_/CLK _33412_/D VGND VGND VPWR VPWR _33412_/Q sky130_fd_sc_hd__dfxtp_1
X_18346_ _20096_/A VGND VGND VPWR VPWR _18346_/X sky130_fd_sc_hd__buf_6
X_30624_ _30624_/A VGND VGND VPWR VPWR _35544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34392_ _35292_/CLK _34392_/D VGND VGND VPWR VPWR _34392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33343_ _33789_/CLK _33343_/D VGND VGND VPWR VPWR _33343_/Q sky130_fd_sc_hd__dfxtp_1
X_36131_ _36132_/CLK _36131_/D VGND VGND VPWR VPWR _36131_/Q sky130_fd_sc_hd__dfxtp_1
X_18277_ _20155_/A VGND VGND VPWR VPWR _18277_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30555_ _23277_/X _35512_/Q _30569_/S VGND VGND VPWR VPWR _30556_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17228_ _35054_/Q _34990_/Q _34926_/Q _34862_/Q _17156_/X _17157_/X VGND VGND VPWR
+ VPWR _17228_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33274_ _36154_/CLK _33274_/D VGND VGND VPWR VPWR _33274_/Q sky130_fd_sc_hd__dfxtp_1
Xinput30 DW[36] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_4
X_36062_ _36062_/CLK _36062_/D VGND VGND VPWR VPWR _36062_/Q sky130_fd_sc_hd__dfxtp_1
X_30486_ _30486_/A VGND VGND VPWR VPWR _35479_/D sky130_fd_sc_hd__clkbuf_1
Xinput41 DW[46] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__buf_6
XFILLER_238_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput52 DW[56] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__buf_8
Xinput63 DW[8] VGND VGND VPWR VPWR input63/X sky130_fd_sc_hd__buf_8
X_35013_ _35780_/CLK _35013_/D VGND VGND VPWR VPWR _35013_/Q sky130_fd_sc_hd__dfxtp_1
X_32225_ _35849_/CLK _32225_/D VGND VGND VPWR VPWR _32225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput74 R2[3] VGND VGND VPWR VPWR input74/X sky130_fd_sc_hd__buf_4
X_17159_ _17159_/A VGND VGND VPWR VPWR _17159_/X sky130_fd_sc_hd__clkbuf_4
Xinput85 RW[2] VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__buf_6
XFILLER_239_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20170_ _20170_/A VGND VGND VPWR VPWR _32128_/D sky130_fd_sc_hd__buf_4
X_32156_ _36200_/CLK _32156_/D VGND VGND VPWR VPWR _32156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31107_ _35774_/Q _29200_/X _31109_/S VGND VGND VPWR VPWR _31108_/A sky130_fd_sc_hd__mux2_1
X_32087_ _35040_/CLK _32087_/D VGND VGND VPWR VPWR _32087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35915_ _35979_/CLK _35915_/D VGND VGND VPWR VPWR _35915_/Q sky130_fd_sc_hd__dfxtp_1
X_31038_ _35741_/Q _29098_/X _31046_/S VGND VGND VPWR VPWR _31039_/A sky130_fd_sc_hd__mux2_1
XFILLER_233_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35846_ _35849_/CLK _35846_/D VGND VGND VPWR VPWR _35846_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23860_ _22910_/X _32472_/Q _23878_/S VGND VGND VPWR VPWR _23861_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_6_0__f_CLK clkbuf_5_0_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_2_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22811_ _20656_/X _22809_/X _22810_/X _20668_/X VGND VGND VPWR VPWR _22811_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35777_ _35777_/CLK _35777_/D VGND VGND VPWR VPWR _35777_/Q sky130_fd_sc_hd__dfxtp_1
X_23791_ _23010_/X _32440_/Q _23805_/S VGND VGND VPWR VPWR _23792_/A sky130_fd_sc_hd__mux2_1
XANTENNA_709 _22532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32989_ _33244_/CLK _32989_/D VGND VGND VPWR VPWR _32989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_253_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _34305_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_246_1415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25530_ _25530_/A VGND VGND VPWR VPWR _33196_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22742_ _35593_/Q _35529_/Q _35465_/Q _35401_/Q _22556_/X _22557_/X VGND VGND VPWR
+ VPWR _22742_/X sky130_fd_sc_hd__mux4_1
X_34728_ _34792_/CLK _34728_/D VGND VGND VPWR VPWR _34728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25461_ _25461_/A VGND VGND VPWR VPWR _31275_/B sky130_fd_sc_hd__buf_8
XFILLER_197_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22673_ _33287_/Q _36167_/Q _33159_/Q _33095_/Q _22364_/X _22365_/X VGND VGND VPWR
+ VPWR _22673_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34659_ _35928_/CLK _34659_/D VGND VGND VPWR VPWR _34659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27200_ _26884_/X _33954_/Q _27218_/S VGND VGND VPWR VPWR _27201_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24412_ _24412_/A VGND VGND VPWR VPWR _32707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28180_ _26934_/X _34418_/Q _28186_/S VGND VGND VPWR VPWR _28181_/A sky130_fd_sc_hd__mux2_1
X_21624_ _21618_/X _21623_/X _21375_/X VGND VGND VPWR VPWR _21646_/A sky130_fd_sc_hd__o21ba_1
X_25392_ _25088_/X _33133_/Q _25408_/S VGND VGND VPWR VPWR _25393_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27131_ _27131_/A VGND VGND VPWR VPWR _33921_/D sky130_fd_sc_hd__clkbuf_1
X_24343_ _32685_/Q _24342_/X _24367_/S VGND VGND VPWR VPWR _24344_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21555_ _21302_/X _21553_/X _21554_/X _21308_/X VGND VGND VPWR VPWR _21555_/X sky130_fd_sc_hd__a22o_1
XFILLER_138_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20506_ _34827_/Q _34763_/Q _34699_/Q _34635_/Q _20294_/X _20295_/X VGND VGND VPWR
+ VPWR _20506_/X sky130_fd_sc_hd__mux4_1
X_27062_ _26881_/X _33889_/Q _27062_/S VGND VGND VPWR VPWR _27063_/A sky130_fd_sc_hd__mux2_1
X_24274_ _32663_/Q _24273_/X _24274_/S VGND VGND VPWR VPWR _24275_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21486_ _21482_/X _21485_/X _21375_/X VGND VGND VPWR VPWR _21510_/A sky130_fd_sc_hd__o21ba_1
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1004 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26013_ _24995_/X _33423_/Q _26029_/S VGND VGND VPWR VPWR _26014_/A sky130_fd_sc_hd__mux2_1
X_20437_ _19454_/A _20435_/X _20436_/X _19459_/A VGND VGND VPWR VPWR _20437_/X sky130_fd_sc_hd__a22o_1
X_23225_ _23225_/A VGND VGND VPWR VPWR _32192_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20368_ _33543_/Q _33479_/Q _33415_/Q _33351_/Q _20129_/X _20130_/X VGND VGND VPWR
+ VPWR _20368_/X sky130_fd_sc_hd__mux4_2
X_23156_ _23156_/A VGND VGND VPWR VPWR _31140_/A sky130_fd_sc_hd__buf_8
XTAP_7036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22107_ _22460_/A VGND VGND VPWR VPWR _22107_/X sky130_fd_sc_hd__buf_2
XFILLER_136_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1108 _36201_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23087_ _23421_/S VGND VGND VPWR VPWR _23115_/S sky130_fd_sc_hd__buf_4
XANTENNA_1119 input53/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27964_ _34316_/Q _24437_/X _27966_/S VGND VGND VPWR VPWR _27965_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20299_ _34564_/Q _32452_/Q _34436_/Q _34372_/Q _20231_/X _20232_/X VGND VGND VPWR
+ VPWR _20299_/X sky130_fd_sc_hd__mux4_1
XTAP_6335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26915_ input24/X VGND VGND VPWR VPWR _26915_/X sky130_fd_sc_hd__clkbuf_4
X_29703_ _29703_/A VGND VGND VPWR VPWR _35108_/D sky130_fd_sc_hd__clkbuf_1
X_22038_ _22034_/X _22037_/X _21761_/X VGND VGND VPWR VPWR _22039_/D sky130_fd_sc_hd__o21ba_1
XTAP_6379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27895_ _34283_/Q _24335_/X _27895_/S VGND VGND VPWR VPWR _27896_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_492_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _35296_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_48_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29634_ _35076_/Q _29219_/X _29644_/S VGND VGND VPWR VPWR _29635_/A sky130_fd_sc_hd__mux2_1
XTAP_5678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26846_ _26846_/A VGND VGND VPWR VPWR _33813_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29565_ _35043_/Q _29117_/X _29581_/S VGND VGND VPWR VPWR _29566_/A sky130_fd_sc_hd__mux2_1
XTAP_4988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26777_ _26777_/A VGND VGND VPWR VPWR _33784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23989_ _22901_/X _32533_/Q _23993_/S VGND VGND VPWR VPWR _23990_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_244_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _34308_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_216_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28516_ _26832_/X _34577_/Q _28528_/S VGND VGND VPWR VPWR _28517_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16530_ _33499_/Q _33435_/Q _33371_/Q _33307_/Q _16417_/X _16418_/X VGND VGND VPWR
+ VPWR _16530_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25728_ _25728_/A VGND VGND VPWR VPWR _33289_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29496_ _29496_/A VGND VGND VPWR VPWR _35010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16461_ _16136_/X _16459_/X _16460_/X _16141_/X VGND VGND VPWR VPWR _16461_/X sky130_fd_sc_hd__a22o_1
X_28447_ _28447_/A VGND VGND VPWR VPWR _34544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25659_ _25659_/A VGND VGND VPWR VPWR _33256_/D sky130_fd_sc_hd__clkbuf_1
X_18200_ _35787_/Q _35147_/Q _34507_/Q _33867_/Q _16108_/X _16109_/X VGND VGND VPWR
+ VPWR _18200_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19180_ _33765_/Q _33701_/Q _33637_/Q _33573_/Q _19143_/X _19144_/X VGND VGND VPWR
+ VPWR _19180_/X sky130_fd_sc_hd__mux4_1
XFILLER_231_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28378_ _28378_/A VGND VGND VPWR VPWR _34511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16392_ _33239_/Q _36119_/Q _33111_/Q _33047_/Q _16352_/X _16353_/X VGND VGND VPWR
+ VPWR _16392_/X sky130_fd_sc_hd__mux4_1
XPHY_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18131_ _18127_/X _18130_/X _17834_/X VGND VGND VPWR VPWR _18153_/A sky130_fd_sc_hd__o21ba_2
XPHY_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27329_ _27329_/A VGND VGND VPWR VPWR _34015_/D sky130_fd_sc_hd__clkbuf_1
XPHY_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18062_ _18058_/X _18061_/X _17867_/X VGND VGND VPWR VPWR _18063_/D sky130_fd_sc_hd__o21ba_1
X_30340_ _23099_/X _35410_/Q _30350_/S VGND VGND VPWR VPWR _30341_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17013_ _17009_/X _17012_/X _16808_/X VGND VGND VPWR VPWR _17014_/D sky130_fd_sc_hd__o21ba_1
XFILLER_208_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30271_ _35378_/Q _29163_/X _30277_/S VGND VGND VPWR VPWR _30272_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32010_ _36194_/CLK _32010_/D VGND VGND VPWR VPWR _32010_/Q sky130_fd_sc_hd__dfxtp_1
X_18964_ _34271_/Q _34207_/Q _34143_/Q _34079_/Q _18683_/X _18684_/X VGND VGND VPWR
+ VPWR _18964_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17915_ _33282_/Q _36162_/Q _33154_/Q _33090_/Q _17764_/X _17765_/X VGND VGND VPWR
+ VPWR _17915_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_1090 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33961_ _34154_/CLK _33961_/D VGND VGND VPWR VPWR _33961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18895_ _18789_/X _18893_/X _18894_/X _18794_/X VGND VGND VPWR VPWR _18895_/X sky130_fd_sc_hd__a22o_1
XTAP_6880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_483_CLK clkbuf_6_3__f_CLK/X VGND VGND VPWR VPWR _35933_/CLK sky130_fd_sc_hd__clkbuf_16
X_35700_ _35700_/CLK _35700_/D VGND VGND VPWR VPWR _35700_/Q sky130_fd_sc_hd__dfxtp_1
X_32912_ _36049_/CLK _32912_/D VGND VGND VPWR VPWR _32912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17846_ _17846_/A VGND VGND VPWR VPWR _17846_/X sky130_fd_sc_hd__buf_4
XFILLER_26_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_868 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33892_ _34149_/CLK _33892_/D VGND VGND VPWR VPWR _33892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35631_ _35822_/CLK _35631_/D VGND VGND VPWR VPWR _35631_/Q sky130_fd_sc_hd__dfxtp_1
X_32843_ _35979_/CLK _32843_/D VGND VGND VPWR VPWR _32843_/Q sky130_fd_sc_hd__dfxtp_1
X_17777_ _35774_/Q _35134_/Q _34494_/Q _33854_/Q _17493_/X _17494_/X VGND VGND VPWR
+ VPWR _17777_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_235_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _32967_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19516_ _35758_/Q _35118_/Q _34478_/Q _33838_/Q _19440_/X _19441_/X VGND VGND VPWR
+ VPWR _19516_/X sky130_fd_sc_hd__mux4_1
X_35562_ _35562_/CLK _35562_/D VGND VGND VPWR VPWR _35562_/Q sky130_fd_sc_hd__dfxtp_1
X_16728_ _16443_/X _16726_/X _16727_/X _16446_/X VGND VGND VPWR VPWR _16728_/X sky130_fd_sc_hd__a22o_1
X_32774_ _36103_/CLK _32774_/D VGND VGND VPWR VPWR _32774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34513_ _36211_/CLK _34513_/D VGND VGND VPWR VPWR _34513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16659_ _16448_/X _16657_/X _16658_/X _16453_/X VGND VGND VPWR VPWR _16659_/X sky130_fd_sc_hd__a22o_1
X_19447_ _20153_/A VGND VGND VPWR VPWR _19447_/X sky130_fd_sc_hd__clkbuf_4
X_31725_ _31725_/A VGND VGND VPWR VPWR _36066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35493_ _35749_/CLK _35493_/D VGND VGND VPWR VPWR _35493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34444_ _35981_/CLK _34444_/D VGND VGND VPWR VPWR _34444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_1432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31656_ _36034_/Q input48/X _31670_/S VGND VGND VPWR VPWR _31657_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19378_ _19372_/X _19377_/X _19094_/X VGND VGND VPWR VPWR _19386_/C sky130_fd_sc_hd__o21ba_1
XFILLER_31_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30607_ _30607_/A VGND VGND VPWR VPWR _35536_/D sky130_fd_sc_hd__clkbuf_1
X_18329_ _18359_/A VGND VGND VPWR VPWR _20070_/A sky130_fd_sc_hd__buf_12
XFILLER_124_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34375_ _35078_/CLK _34375_/D VGND VGND VPWR VPWR _34375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31587_ _31587_/A VGND VGND VPWR VPWR _36001_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1048 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36114_ _36114_/CLK _36114_/D VGND VGND VPWR VPWR _36114_/Q sky130_fd_sc_hd__dfxtp_1
X_21340_ _33505_/Q _33441_/Q _33377_/Q _33313_/Q _21017_/X _21018_/X VGND VGND VPWR
+ VPWR _21340_/X sky130_fd_sc_hd__mux4_1
X_30538_ _23250_/X _35504_/Q _30548_/S VGND VGND VPWR VPWR _30539_/A sky130_fd_sc_hd__mux2_1
X_33326_ _36147_/CLK _33326_/D VGND VGND VPWR VPWR _33326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36045_ _36045_/CLK _36045_/D VGND VGND VPWR VPWR _36045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21271_ _21265_/X _21270_/X _21022_/X VGND VGND VPWR VPWR _21293_/A sky130_fd_sc_hd__o21ba_1
X_30469_ _23090_/X _35471_/Q _30485_/S VGND VGND VPWR VPWR _30470_/A sky130_fd_sc_hd__mux2_1
X_33257_ _36136_/CLK _33257_/D VGND VGND VPWR VPWR _33257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20222_ _35778_/Q _35138_/Q _34498_/Q _33858_/Q _20146_/X _20147_/X VGND VGND VPWR
+ VPWR _20222_/X sky130_fd_sc_hd__mux4_1
X_23010_ input37/X VGND VGND VPWR VPWR _23010_/X sky130_fd_sc_hd__buf_2
XFILLER_85_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32208_ _35638_/CLK _32208_/D VGND VGND VPWR VPWR _32208_/Q sky130_fd_sc_hd__dfxtp_1
X_33188_ _35876_/CLK _33188_/D VGND VGND VPWR VPWR _33188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20153_ _20153_/A VGND VGND VPWR VPWR _20153_/X sky130_fd_sc_hd__clkbuf_4
X_32139_ _35815_/CLK _32139_/D VGND VGND VPWR VPWR _32139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24961_ _23034_/X _32960_/Q _24979_/S VGND VGND VPWR VPWR _24962_/A sky130_fd_sc_hd__mux2_1
X_20084_ _20078_/X _20083_/X _19800_/X VGND VGND VPWR VPWR _20092_/C sky130_fd_sc_hd__o21ba_1
XFILLER_135_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26700_ _33748_/Q _24264_/X _26706_/S VGND VGND VPWR VPWR _26701_/A sky130_fd_sc_hd__mux2_1
XTAP_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_474_CLK clkbuf_6_8__f_CLK/X VGND VGND VPWR VPWR _35938_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23912_ _22988_/X _32497_/Q _23920_/S VGND VGND VPWR VPWR _23913_/A sky130_fd_sc_hd__mux2_1
X_27680_ _34181_/Q _24416_/X _27688_/S VGND VGND VPWR VPWR _27681_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24892_ _24892_/A VGND VGND VPWR VPWR _32927_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26631_ _25109_/X _33716_/Q _26633_/S VGND VGND VPWR VPWR _26632_/A sky130_fd_sc_hd__mux2_1
X_23843_ _22886_/X _32464_/Q _23857_/S VGND VGND VPWR VPWR _23844_/A sky130_fd_sc_hd__mux2_1
XTAP_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35829_ _35829_/CLK _35829_/D VGND VGND VPWR VPWR _35829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_226_CLK clkbuf_6_55__f_CLK/X VGND VGND VPWR VPWR _35843_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_506 _17900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_517 _17970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29350_ _29350_/A VGND VGND VPWR VPWR _34941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26562_ _25007_/X _33683_/Q _26570_/S VGND VGND VPWR VPWR _26563_/A sky130_fd_sc_hd__mux2_1
XANTENNA_528 _18034_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23774_ _22985_/X _32432_/Q _23784_/S VGND VGND VPWR VPWR _23775_/A sky130_fd_sc_hd__mux2_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20986_ _20736_/X _20982_/X _20985_/X _20741_/X VGND VGND VPWR VPWR _20986_/X sky130_fd_sc_hd__a22o_1
XANTENNA_539 _20160_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28301_ _28301_/A VGND VGND VPWR VPWR _34475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25513_ _25513_/A VGND VGND VPWR VPWR _33188_/D sky130_fd_sc_hd__clkbuf_1
X_22725_ _33801_/Q _33737_/Q _33673_/Q _33609_/Q _22502_/X _22503_/X VGND VGND VPWR
+ VPWR _22725_/X sky130_fd_sc_hd__mux4_1
X_29281_ _29281_/A VGND VGND VPWR VPWR _34908_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26493_ _25106_/X _33651_/Q _26497_/S VGND VGND VPWR VPWR _26494_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28232_ _27011_/X _34443_/Q _28236_/S VGND VGND VPWR VPWR _28233_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25444_ _25165_/X _33158_/Q _25450_/S VGND VGND VPWR VPWR _25445_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22656_ _34822_/Q _34758_/Q _34694_/Q _34630_/Q _22594_/X _22595_/X VGND VGND VPWR
+ VPWR _22656_/X sky130_fd_sc_hd__mux4_1
XFILLER_186_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28163_ _26909_/X _34410_/Q _28165_/S VGND VGND VPWR VPWR _28164_/A sky130_fd_sc_hd__mux2_1
X_21607_ _21607_/A VGND VGND VPWR VPWR _21607_/X sky130_fd_sc_hd__clkbuf_4
X_25375_ _25063_/X _33125_/Q _25387_/S VGND VGND VPWR VPWR _25376_/A sky130_fd_sc_hd__mux2_1
X_22587_ _35844_/Q _32223_/Q _35716_/Q _35652_/Q _22266_/X _22267_/X VGND VGND VPWR
+ VPWR _22587_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27114_ _27114_/A VGND VGND VPWR VPWR _33913_/D sky130_fd_sc_hd__clkbuf_1
X_24326_ input19/X VGND VGND VPWR VPWR _24326_/X sky130_fd_sc_hd__buf_4
XFILLER_103_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28094_ _28094_/A VGND VGND VPWR VPWR _34377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21538_ _35302_/Q _35238_/Q _35174_/Q _32294_/Q _21253_/X _21254_/X VGND VGND VPWR
+ VPWR _21538_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27045_ _27045_/A VGND VGND VPWR VPWR _33880_/D sky130_fd_sc_hd__clkbuf_1
X_24257_ _24257_/A VGND VGND VPWR VPWR _32657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21469_ _34788_/Q _34724_/Q _34660_/Q _34596_/Q _21182_/X _21183_/X VGND VGND VPWR
+ VPWR _21469_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23208_ _23346_/S VGND VGND VPWR VPWR _23235_/S sky130_fd_sc_hd__buf_4
XFILLER_134_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24188_ _22994_/X _32627_/Q _24192_/S VGND VGND VPWR VPWR _24189_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23139_ input9/X VGND VGND VPWR VPWR _23139_/X sky130_fd_sc_hd__buf_4
XTAP_6121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28996_ _34805_/Q _24366_/X _28996_/S VGND VGND VPWR VPWR _28997_/A sky130_fd_sc_hd__mux2_1
XTAP_6143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27947_ _27947_/A VGND VGND VPWR VPWR _34307_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17700_ _17855_/A VGND VGND VPWR VPWR _17700_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_465_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _35750_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_5464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18680_ _18680_/A _18680_/B _18680_/C _18680_/D VGND VGND VPWR VPWR _18681_/A sky130_fd_sc_hd__or4_4
X_27878_ _27878_/A VGND VGND VPWR VPWR _34274_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29617_ _35068_/Q _29194_/X _29623_/S VGND VGND VPWR VPWR _29618_/A sky130_fd_sc_hd__mux2_1
X_17631_ _33018_/Q _32954_/Q _32890_/Q _32826_/Q _17342_/X _17343_/X VGND VGND VPWR
+ VPWR _17631_/X sky130_fd_sc_hd__mux4_1
X_26829_ input23/X VGND VGND VPWR VPWR _26829_/X sky130_fd_sc_hd__buf_4
XTAP_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_217_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _35781_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17562_ _33272_/Q _36152_/Q _33144_/Q _33080_/Q _17411_/X _17412_/X VGND VGND VPWR
+ VPWR _17562_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29548_ _35035_/Q _29092_/X _29560_/S VGND VGND VPWR VPWR _29549_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_1031 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19301_ _33192_/Q _32552_/Q _35944_/Q _35880_/Q _19021_/X _19022_/X VGND VGND VPWR
+ VPWR _19301_/X sky130_fd_sc_hd__mux4_1
X_16513_ _33178_/Q _32538_/Q _35930_/Q _35866_/Q _16368_/X _16369_/X VGND VGND VPWR
+ VPWR _16513_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1015 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17493_ _17846_/A VGND VGND VPWR VPWR _17493_/X sky130_fd_sc_hd__buf_4
XFILLER_16_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29479_ _29479_/A VGND VGND VPWR VPWR _35002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31510_ _23294_/X _35965_/Q _31514_/S VGND VGND VPWR VPWR _31511_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19232_ _33190_/Q _32550_/Q _35942_/Q _35878_/Q _19021_/X _19022_/X VGND VGND VPWR
+ VPWR _19232_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16444_ _34776_/Q _34712_/Q _34648_/Q _34584_/Q _16229_/X _16230_/X VGND VGND VPWR
+ VPWR _16444_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32490_ _36075_/CLK _32490_/D VGND VGND VPWR VPWR _32490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19163_ _35748_/Q _35108_/Q _34468_/Q _33828_/Q _19087_/X _19088_/X VGND VGND VPWR
+ VPWR _19163_/X sky130_fd_sc_hd__mux4_1
X_31441_ _23130_/X _35932_/Q _31451_/S VGND VGND VPWR VPWR _31442_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16375_ _16074_/X _16373_/X _16374_/X _16084_/X VGND VGND VPWR VPWR _16375_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_1335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18114_ _15997_/X _18112_/X _18113_/X _16003_/X VGND VGND VPWR VPWR _18114_/X sky130_fd_sc_hd__a22o_1
XFILLER_223_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34160_ _34286_/CLK _34160_/D VGND VGND VPWR VPWR _34160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31372_ _31372_/A VGND VGND VPWR VPWR _35899_/D sky130_fd_sc_hd__clkbuf_1
X_19094_ _20153_/A VGND VGND VPWR VPWR _19094_/X sky130_fd_sc_hd__buf_2
XFILLER_144_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30323_ _35403_/Q _29240_/X _30327_/S VGND VGND VPWR VPWR _30324_/A sky130_fd_sc_hd__mux2_1
X_18045_ _32518_/Q _32390_/Q _32070_/Q _36038_/Q _17982_/X _17770_/X VGND VGND VPWR
+ VPWR _18045_/X sky130_fd_sc_hd__mux4_1
X_33111_ _36118_/CLK _33111_/D VGND VGND VPWR VPWR _33111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34091_ _34282_/CLK _34091_/D VGND VGND VPWR VPWR _34091_/Q sky130_fd_sc_hd__dfxtp_1
X_33042_ _36114_/CLK _33042_/D VGND VGND VPWR VPWR _33042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30254_ _35370_/Q _29138_/X _30256_/S VGND VGND VPWR VPWR _30255_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30185_ _30185_/A VGND VGND VPWR VPWR _35337_/D sky130_fd_sc_hd__clkbuf_1
X_19996_ _20130_/A VGND VGND VPWR VPWR _19996_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_119_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18947_ _35550_/Q _35486_/Q _35422_/Q _35358_/Q _18844_/X _18845_/X VGND VGND VPWR
+ VPWR _18947_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34993_ _35826_/CLK _34993_/D VGND VGND VPWR VPWR _34993_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_13__f_CLK clkbuf_5_6_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_57_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_95_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_456_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _34792_/CLK sky130_fd_sc_hd__clkbuf_16
X_33944_ _36185_/CLK _33944_/D VGND VGND VPWR VPWR _33944_/Q sky130_fd_sc_hd__dfxtp_1
X_18878_ _35548_/Q _35484_/Q _35420_/Q _35356_/Q _18844_/X _18845_/X VGND VGND VPWR
+ VPWR _18878_/X sky130_fd_sc_hd__mux4_1
XFILLER_227_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17829_ _17829_/A VGND VGND VPWR VPWR _17829_/X sky130_fd_sc_hd__buf_4
X_33875_ _36228_/CLK _33875_/D VGND VGND VPWR VPWR _33875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_208_CLK clkbuf_6_52__f_CLK/X VGND VGND VPWR VPWR _35849_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_48_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35614_ _35807_/CLK _35614_/D VGND VGND VPWR VPWR _35614_/Q sky130_fd_sc_hd__dfxtp_1
X_20840_ _33747_/Q _33683_/Q _33619_/Q _33555_/Q _20737_/X _20738_/X VGND VGND VPWR
+ VPWR _20840_/X sky130_fd_sc_hd__mux4_1
X_32826_ _32954_/CLK _32826_/D VGND VGND VPWR VPWR _32826_/Q sky130_fd_sc_hd__dfxtp_1
X_35545_ _35801_/CLK _35545_/D VGND VGND VPWR VPWR _35545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20771_ _20765_/X _20770_/X _20700_/X VGND VGND VPWR VPWR _20772_/D sky130_fd_sc_hd__o21ba_1
X_32757_ _36085_/CLK _32757_/D VGND VGND VPWR VPWR _32757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22510_ _34050_/Q _33986_/Q _33922_/Q _32258_/Q _22326_/X _22327_/X VGND VGND VPWR
+ VPWR _22510_/X sky130_fd_sc_hd__mux4_1
X_31708_ _31708_/A VGND VGND VPWR VPWR _36058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35476_ _35927_/CLK _35476_/D VGND VGND VPWR VPWR _35476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23490_ _23559_/S VGND VGND VPWR VPWR _23509_/S sky130_fd_sc_hd__buf_4
XFILLER_149_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32688_ _33009_/CLK _32688_/D VGND VGND VPWR VPWR _32688_/Q sky130_fd_sc_hd__dfxtp_1
X_22441_ _22369_/X _22439_/X _22440_/X _22373_/X VGND VGND VPWR VPWR _22441_/X sky130_fd_sc_hd__a22o_1
X_34427_ _35579_/CLK _34427_/D VGND VGND VPWR VPWR _34427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31639_ _36026_/Q input39/X _31649_/S VGND VGND VPWR VPWR _31640_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25160_ _25159_/X _33028_/Q _25175_/S VGND VGND VPWR VPWR _25161_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22372_ _33022_/Q _32958_/Q _32894_/Q _32830_/Q _22295_/X _22296_/X VGND VGND VPWR
+ VPWR _22372_/X sky130_fd_sc_hd__mux4_1
X_34358_ _35319_/CLK _34358_/D VGND VGND VPWR VPWR _34358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24111_ _22875_/X _32590_/Q _24129_/S VGND VGND VPWR VPWR _24112_/A sky130_fd_sc_hd__mux2_1
X_21323_ _33184_/Q _32544_/Q _35936_/Q _35872_/Q _21321_/X _21322_/X VGND VGND VPWR
+ VPWR _21323_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33309_ _33946_/CLK _33309_/D VGND VGND VPWR VPWR _33309_/Q sky130_fd_sc_hd__dfxtp_1
X_25091_ input26/X VGND VGND VPWR VPWR _25091_/X sky130_fd_sc_hd__buf_2
X_34289_ _34289_/CLK _34289_/D VGND VGND VPWR VPWR _34289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36028_ _36028_/CLK _36028_/D VGND VGND VPWR VPWR _36028_/Q sky130_fd_sc_hd__dfxtp_1
X_24042_ _22979_/X _32558_/Q _24056_/S VGND VGND VPWR VPWR _24043_/A sky130_fd_sc_hd__mux2_1
X_21254_ _21607_/A VGND VGND VPWR VPWR _21254_/X sky130_fd_sc_hd__buf_4
XFILLER_85_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20205_ _34306_/Q _34242_/Q _34178_/Q _34114_/Q _20095_/X _20096_/X VGND VGND VPWR
+ VPWR _20205_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28850_ _28850_/A VGND VGND VPWR VPWR _34735_/D sky130_fd_sc_hd__clkbuf_1
X_21185_ _35292_/Q _35228_/Q _35164_/Q _32284_/Q _20900_/X _20901_/X VGND VGND VPWR
+ VPWR _21185_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20136_ _32768_/Q _32704_/Q _32640_/Q _36096_/Q _19925_/X _20062_/X VGND VGND VPWR
+ VPWR _20136_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27801_ _27801_/A VGND VGND VPWR VPWR _34238_/D sky130_fd_sc_hd__clkbuf_1
X_28781_ _28781_/A VGND VGND VPWR VPWR _34702_/D sky130_fd_sc_hd__clkbuf_1
X_25993_ _25165_/X _33414_/Q _25999_/S VGND VGND VPWR VPWR _25994_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_447_CLK clkbuf_leaf_50_CLK/A VGND VGND VPWR VPWR _32994_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_86_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27732_ _27732_/A VGND VGND VPWR VPWR _34205_/D sky130_fd_sc_hd__clkbuf_1
X_20067_ _20067_/A VGND VGND VPWR VPWR _20067_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24944_ _23010_/X _32952_/Q _24958_/S VGND VGND VPWR VPWR _24945_/A sky130_fd_sc_hd__mux2_1
XTAP_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_969 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27663_ _34173_/Q _24391_/X _27667_/S VGND VGND VPWR VPWR _27664_/A sky130_fd_sc_hd__mux2_1
XTAP_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24875_ _24875_/A VGND VGND VPWR VPWR _32919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29402_ _23111_/X _34966_/Q _29404_/S VGND VGND VPWR VPWR _29403_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26614_ _26683_/S VGND VGND VPWR VPWR _26633_/S sky130_fd_sc_hd__buf_6
XTAP_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23826_ _23062_/X _32457_/Q _23826_/S VGND VGND VPWR VPWR _23827_/A sky130_fd_sc_hd__mux2_1
XANTENNA_303 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_314 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27594_ _34140_/Q _24289_/X _27604_/S VGND VGND VPWR VPWR _27595_/A sky130_fd_sc_hd__mux2_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_325 _32141_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_336 _32141_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_347 _36205_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26545_ _25183_/X _33676_/Q _26547_/S VGND VGND VPWR VPWR _26546_/A sky130_fd_sc_hd__mux2_1
X_29333_ _29333_/A VGND VGND VPWR VPWR _34933_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_358 _36207_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23757_ _22960_/X _32424_/Q _23763_/S VGND VGND VPWR VPWR _23758_/A sky130_fd_sc_hd__mux2_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_369 _36207_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20969_ _22532_/A VGND VGND VPWR VPWR _20969_/X sky130_fd_sc_hd__buf_4
XFILLER_13_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22708_ _22704_/X _22707_/X _22442_/X _22443_/X VGND VGND VPWR VPWR _22723_/B sky130_fd_sc_hd__o211a_1
X_29264_ _29264_/A VGND VGND VPWR VPWR _34900_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26476_ _25081_/X _33643_/Q _26476_/S VGND VGND VPWR VPWR _26477_/A sky130_fd_sc_hd__mux2_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23688_ _32393_/Q _23333_/X _23688_/S VGND VGND VPWR VPWR _23689_/A sky130_fd_sc_hd__mux2_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28215_ _28215_/A VGND VGND VPWR VPWR _34434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25427_ _25140_/X _33150_/Q _25429_/S VGND VGND VPWR VPWR _25428_/A sky130_fd_sc_hd__mux2_1
X_22639_ _34054_/Q _33990_/Q _33926_/Q _32262_/Q _22326_/X _22327_/X VGND VGND VPWR
+ VPWR _22639_/X sky130_fd_sc_hd__mux4_1
X_29195_ _34876_/Q _29194_/X _29204_/S VGND VGND VPWR VPWR _29196_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16160_ _33168_/Q _32528_/Q _35920_/Q _35856_/Q _16063_/X _16065_/X VGND VGND VPWR
+ VPWR _16160_/X sky130_fd_sc_hd__mux4_1
X_28146_ _28236_/S VGND VGND VPWR VPWR _28165_/S sky130_fd_sc_hd__buf_4
XFILLER_70_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25358_ _25038_/X _33117_/Q _25366_/S VGND VGND VPWR VPWR _25359_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24309_ _32674_/Q _24307_/X _24336_/S VGND VGND VPWR VPWR _24310_/A sky130_fd_sc_hd__mux2_1
X_28077_ _26981_/X _34369_/Q _28093_/S VGND VGND VPWR VPWR _28078_/A sky130_fd_sc_hd__mux2_1
X_16091_ _34510_/Q _32398_/Q _34382_/Q _34318_/Q _16088_/X _16090_/X VGND VGND VPWR
+ VPWR _16091_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25289_ _25137_/X _33085_/Q _25293_/S VGND VGND VPWR VPWR _25290_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27028_ _27028_/A VGND VGND VPWR VPWR _33872_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19850_ _20203_/A VGND VGND VPWR VPWR _19850_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_134_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18801_ _18795_/X _18800_/X _18722_/X VGND VGND VPWR VPWR _18825_/A sky130_fd_sc_hd__o21ba_1
X_19781_ _20134_/A VGND VGND VPWR VPWR _19781_/X sky130_fd_sc_hd__buf_2
XFILLER_150_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28979_ _28979_/A VGND VGND VPWR VPWR _34796_/D sky130_fd_sc_hd__clkbuf_1
X_16993_ _16987_/X _16992_/X _16783_/X _16784_/X VGND VGND VPWR VPWR _17014_/B sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_438_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _36134_/CLK sky130_fd_sc_hd__clkbuf_16
X_18732_ _18726_/X _18729_/X _18730_/X _18731_/X VGND VGND VPWR VPWR _18757_/B sky130_fd_sc_hd__o211a_2
XTAP_5250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31990_ _36200_/CLK _31990_/D VGND VGND VPWR VPWR _31990_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18663_ _18656_/X _18662_/X _18340_/X _18342_/X VGND VGND VPWR VPWR _18680_/B sky130_fd_sc_hd__o211a_1
X_30941_ _35695_/Q _29154_/X _30953_/S VGND VGND VPWR VPWR _30942_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17614_ _17507_/X _17612_/X _17613_/X _17512_/X VGND VGND VPWR VPWR _17614_/X sky130_fd_sc_hd__a22o_1
XFILLER_92_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33660_ _34044_/CLK _33660_/D VGND VGND VPWR VPWR _33660_/Q sky130_fd_sc_hd__dfxtp_1
X_30872_ _35662_/Q _29048_/X _30890_/S VGND VGND VPWR VPWR _30873_/A sky130_fd_sc_hd__mux2_1
X_18594_ _35540_/Q _35476_/Q _35412_/Q _35348_/Q _18491_/X _18492_/X VGND VGND VPWR
+ VPWR _18594_/X sky130_fd_sc_hd__mux4_1
XFILLER_188_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32611_ _36067_/CLK _32611_/D VGND VGND VPWR VPWR _32611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17545_ _17541_/X _17544_/X _17514_/X VGND VGND VPWR VPWR _17546_/D sky130_fd_sc_hd__o21ba_1
XFILLER_63_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33591_ _34293_/CLK _33591_/D VGND VGND VPWR VPWR _33591_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_870 _24987_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35330_ _35330_/CLK _35330_/D VGND VGND VPWR VPWR _35330_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_881 _25084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17476_ _17829_/A VGND VGND VPWR VPWR _17476_/X sky130_fd_sc_hd__buf_4
X_32542_ _35935_/CLK _32542_/D VGND VGND VPWR VPWR _32542_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_892 _25597_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19215_ _33510_/Q _33446_/Q _33382_/Q _33318_/Q _19070_/X _19071_/X VGND VGND VPWR
+ VPWR _19215_/X sky130_fd_sc_hd__mux4_1
X_35261_ _35326_/CLK _35261_/D VGND VGND VPWR VPWR _35261_/Q sky130_fd_sc_hd__dfxtp_1
X_16427_ _32472_/Q _32344_/Q _32024_/Q _35992_/Q _16217_/X _16358_/X VGND VGND VPWR
+ VPWR _16427_/X sky130_fd_sc_hd__mux4_1
X_32473_ _33635_/CLK _32473_/D VGND VGND VPWR VPWR _32473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34212_ _34276_/CLK _34212_/D VGND VGND VPWR VPWR _34212_/Q sky130_fd_sc_hd__dfxtp_1
X_31424_ _23105_/X _35924_/Q _31430_/S VGND VGND VPWR VPWR _31425_/A sky130_fd_sc_hd__mux2_1
X_16358_ _17770_/A VGND VGND VPWR VPWR _16358_/X sky130_fd_sc_hd__buf_4
X_19146_ _34276_/Q _34212_/Q _34148_/Q _34084_/Q _19036_/X _19037_/X VGND VGND VPWR
+ VPWR _19146_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_784 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35192_ _35320_/CLK _35192_/D VGND VGND VPWR VPWR _35192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31355_ _31355_/A VGND VGND VPWR VPWR _35891_/D sky130_fd_sc_hd__clkbuf_1
X_34143_ _35675_/CLK _34143_/D VGND VGND VPWR VPWR _34143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16289_ _35796_/Q _32170_/Q _35668_/Q _35604_/Q _16254_/X _16255_/X VGND VGND VPWR
+ VPWR _16289_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19077_ _32738_/Q _32674_/Q _32610_/Q _36066_/Q _18866_/X _19003_/X VGND VGND VPWR
+ VPWR _19077_/X sky130_fd_sc_hd__mux4_1
XFILLER_246_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30306_ _30306_/A VGND VGND VPWR VPWR _35394_/D sky130_fd_sc_hd__clkbuf_1
X_18028_ _17855_/X _18026_/X _18027_/X _17858_/X VGND VGND VPWR VPWR _18028_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31286_ _31286_/A VGND VGND VPWR VPWR _35858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34074_ _34074_/CLK _34074_/D VGND VGND VPWR VPWR _34074_/Q sky130_fd_sc_hd__dfxtp_1
X_33025_ _36159_/CLK _33025_/D VGND VGND VPWR VPWR _33025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30237_ _30327_/S VGND VGND VPWR VPWR _30256_/S sky130_fd_sc_hd__buf_4
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30168_ _35329_/Q _29210_/X _30184_/S VGND VGND VPWR VPWR _30169_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19979_ _35067_/Q _35003_/Q _34939_/Q _34875_/Q _19809_/X _19810_/X VGND VGND VPWR
+ VPWR _19979_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_429_CLK clkbuf_6_36__f_CLK/X VGND VGND VPWR VPWR _36139_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_132_1231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30099_ _30099_/A VGND VGND VPWR VPWR _35296_/D sky130_fd_sc_hd__clkbuf_1
X_22990_ _22990_/A VGND VGND VPWR VPWR _32049_/D sky130_fd_sc_hd__clkbuf_1
X_34976_ _35040_/CLK _34976_/D VGND VGND VPWR VPWR _34976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1280 _17834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1291 _17847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33927_ _34816_/CLK _33927_/D VGND VGND VPWR VPWR _33927_/Q sky130_fd_sc_hd__dfxtp_1
X_21941_ _32498_/Q _32370_/Q _32050_/Q _36018_/Q _21876_/X _21664_/X VGND VGND VPWR
+ VPWR _21941_/X sky130_fd_sc_hd__mux4_1
XFILLER_167_1305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24660_ _24660_/A VGND VGND VPWR VPWR _32818_/D sky130_fd_sc_hd__clkbuf_1
X_33858_ _35777_/CLK _33858_/D VGND VGND VPWR VPWR _33858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21872_ _22578_/A VGND VGND VPWR VPWR _21872_/X sky130_fd_sc_hd__buf_6
XFILLER_215_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23611_ _32356_/Q _23175_/X _23625_/S VGND VGND VPWR VPWR _23612_/A sky130_fd_sc_hd__mux2_1
X_20823_ _35730_/Q _35090_/Q _34450_/Q _33810_/Q _20649_/X _20651_/X VGND VGND VPWR
+ VPWR _20823_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32809_ _36137_/CLK _32809_/D VGND VGND VPWR VPWR _32809_/Q sky130_fd_sc_hd__dfxtp_1
X_24591_ _24591_/A VGND VGND VPWR VPWR _32785_/D sky130_fd_sc_hd__clkbuf_1
X_33789_ _33789_/CLK _33789_/D VGND VGND VPWR VPWR _33789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26330_ _26330_/A VGND VGND VPWR VPWR _33573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23542_ _23542_/A VGND VGND VPWR VPWR _32324_/D sky130_fd_sc_hd__clkbuf_1
X_35528_ _35975_/CLK _35528_/D VGND VGND VPWR VPWR _35528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20754_ _20626_/X _20752_/X _20753_/X _20637_/X VGND VGND VPWR VPWR _20754_/X sky130_fd_sc_hd__a22o_1
XFILLER_208_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26261_ _25162_/X _33541_/Q _26269_/S VGND VGND VPWR VPWR _26262_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35459_ _35909_/CLK _35459_/D VGND VGND VPWR VPWR _35459_/Q sky130_fd_sc_hd__dfxtp_1
X_23473_ _23473_/A VGND VGND VPWR VPWR _32291_/D sky130_fd_sc_hd__clkbuf_1
X_20685_ _20674_/X _20677_/X _20682_/X _20684_/X VGND VGND VPWR VPWR _20685_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28000_ _28000_/A VGND VGND VPWR VPWR _34332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25212_ _25022_/X _33048_/Q _25230_/S VGND VGND VPWR VPWR _25213_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22424_ _22424_/A _22424_/B _22424_/C _22424_/D VGND VGND VPWR VPWR _22425_/A sky130_fd_sc_hd__or4_4
X_26192_ _25060_/X _33508_/Q _26206_/S VGND VGND VPWR VPWR _26193_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25143_ input44/X VGND VGND VPWR VPWR _25143_/X sky130_fd_sc_hd__buf_2
X_22355_ _34302_/Q _34238_/Q _34174_/Q _34110_/Q _22042_/X _22043_/X VGND VGND VPWR
+ VPWR _22355_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21306_ _22503_/A VGND VGND VPWR VPWR _21306_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_156_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29951_ _35226_/Q _29089_/X _29965_/S VGND VGND VPWR VPWR _29952_/A sky130_fd_sc_hd__mux2_1
X_25074_ _25074_/A VGND VGND VPWR VPWR _33000_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22286_ _22148_/X _22284_/X _22285_/X _22153_/X VGND VGND VPWR VPWR _22286_/X sky130_fd_sc_hd__a22o_1
XFILLER_156_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28902_ _28902_/A VGND VGND VPWR VPWR _34760_/D sky130_fd_sc_hd__clkbuf_1
X_24025_ _22954_/X _32550_/Q _24035_/S VGND VGND VPWR VPWR _24026_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21237_ _22430_/A VGND VGND VPWR VPWR _21237_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_85_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29882_ _29882_/A VGND VGND VPWR VPWR _35193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28833_ _28833_/A VGND VGND VPWR VPWR _34727_/D sky130_fd_sc_hd__clkbuf_1
X_21168_ _33244_/Q _36124_/Q _33116_/Q _33052_/Q _20952_/X _20953_/X VGND VGND VPWR
+ VPWR _21168_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20119_ _19802_/X _20117_/X _20118_/X _19805_/X VGND VGND VPWR VPWR _20119_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28764_ _26999_/X _34695_/Q _28768_/S VGND VGND VPWR VPWR _28765_/A sky130_fd_sc_hd__mux2_1
X_25976_ _25140_/X _33406_/Q _25978_/S VGND VGND VPWR VPWR _25977_/A sky130_fd_sc_hd__mux2_1
X_21099_ _22465_/A VGND VGND VPWR VPWR _21099_/X sky130_fd_sc_hd__buf_4
XFILLER_213_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27715_ _27715_/A VGND VGND VPWR VPWR _34197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24927_ _22985_/X _32944_/Q _24937_/S VGND VGND VPWR VPWR _24928_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28695_ _26897_/X _34662_/Q _28705_/S VGND VGND VPWR VPWR _28696_/A sky130_fd_sc_hd__mux2_1
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24858_ _22883_/X _32911_/Q _24874_/S VGND VGND VPWR VPWR _24859_/A sky130_fd_sc_hd__mux2_1
XANTENNA_100 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27646_ _34165_/Q _24366_/X _27646_/S VGND VGND VPWR VPWR _27647_/A sky130_fd_sc_hd__mux2_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1080 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_111 _32129_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23809_ _23809_/A VGND VGND VPWR VPWR _32448_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_133 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27577_ _34132_/Q _24264_/X _27583_/S VGND VGND VPWR VPWR _27578_/A sky130_fd_sc_hd__mux2_1
XANTENNA_144 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24789_ _24789_/A VGND VGND VPWR VPWR _32878_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_166 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17330_ _17330_/A VGND VGND VPWR VPWR _31985_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26528_ _26528_/A VGND VGND VPWR VPWR _33667_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_177 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29316_ _23241_/X _34925_/Q _29332_/S VGND VGND VPWR VPWR _29317_/A sky130_fd_sc_hd__mux2_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_188 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_199 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17261_ _17154_/X _17259_/X _17260_/X _17159_/X VGND VGND VPWR VPWR _17261_/X sky130_fd_sc_hd__a22o_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29247_ _34893_/Q _29246_/X _29247_/S VGND VGND VPWR VPWR _29248_/A sky130_fd_sc_hd__mux2_1
X_26459_ _26459_/A VGND VGND VPWR VPWR _33634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16212_ _16208_/X _16211_/X _16011_/X VGND VGND VPWR VPWR _16238_/A sky130_fd_sc_hd__o21ba_1
X_19000_ _18796_/X _18998_/X _18999_/X _18799_/X VGND VGND VPWR VPWR _19000_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29178_ _29178_/A VGND VGND VPWR VPWR _34870_/D sky130_fd_sc_hd__clkbuf_1
X_17192_ _17188_/X _17191_/X _17161_/X VGND VGND VPWR VPWR _17193_/D sky130_fd_sc_hd__o21ba_1
XFILLER_220_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_957 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16143_ _17860_/A VGND VGND VPWR VPWR _16143_/X sky130_fd_sc_hd__buf_4
X_28129_ _28129_/A VGND VGND VPWR VPWR _34393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31140_ _31140_/A _31140_/B VGND VGND VPWR VPWR _31273_/S sky130_fd_sc_hd__nor2_8
XFILLER_5_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16074_ _17149_/A VGND VGND VPWR VPWR _16074_/X sky130_fd_sc_hd__buf_4
XFILLER_115_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19902_ _19647_/X _19900_/X _19901_/X _19650_/X VGND VGND VPWR VPWR _19902_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31071_ _31071_/A VGND VGND VPWR VPWR _35756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30022_ _35260_/Q _29194_/X _30028_/S VGND VGND VPWR VPWR _30023_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19833_ _35767_/Q _35127_/Q _34487_/Q _33847_/Q _19793_/X _19794_/X VGND VGND VPWR
+ VPWR _19833_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34830_ _35026_/CLK _34830_/D VGND VGND VPWR VPWR _34830_/Q sky130_fd_sc_hd__dfxtp_1
X_19764_ _34805_/Q _34741_/Q _34677_/Q _34613_/Q _19588_/X _19589_/X VGND VGND VPWR
+ VPWR _19764_/X sky130_fd_sc_hd__mux4_1
X_16976_ _16976_/A _16976_/B _16976_/C _16976_/D VGND VGND VPWR VPWR _16977_/A sky130_fd_sc_hd__or4_4
XFILLER_232_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18715_ _34264_/Q _34200_/Q _34136_/Q _34072_/Q _18683_/X _18684_/X VGND VGND VPWR
+ VPWR _18715_/X sky130_fd_sc_hd__mux4_1
X_34761_ _35337_/CLK _34761_/D VGND VGND VPWR VPWR _34761_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 DW[14] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__buf_6
XTAP_5091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31973_ _34970_/CLK _31973_/D VGND VGND VPWR VPWR _31973_/Q sky130_fd_sc_hd__dfxtp_1
X_19695_ _34547_/Q _32435_/Q _34419_/Q _34355_/Q _19525_/X _19526_/X VGND VGND VPWR
+ VPWR _19695_/X sky130_fd_sc_hd__mux4_1
XFILLER_209_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33712_ _33775_/CLK _33712_/D VGND VGND VPWR VPWR _33712_/Q sky130_fd_sc_hd__dfxtp_1
X_18646_ _34006_/Q _33942_/Q _33878_/Q _32150_/Q _18614_/X _18615_/X VGND VGND VPWR
+ VPWR _18646_/X sky130_fd_sc_hd__mux4_1
X_30924_ _35687_/Q _29129_/X _30932_/S VGND VGND VPWR VPWR _30925_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34692_ _35332_/CLK _34692_/D VGND VGND VPWR VPWR _34692_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33643_ _34281_/CLK _33643_/D VGND VGND VPWR VPWR _33643_/Q sky130_fd_sc_hd__dfxtp_1
X_18577_ _18443_/X _18575_/X _18576_/X _18446_/X VGND VGND VPWR VPWR _18577_/X sky130_fd_sc_hd__a22o_1
X_30855_ _30855_/A VGND VGND VPWR VPWR _35654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17528_ _32503_/Q _32375_/Q _32055_/Q _36023_/Q _17276_/X _17417_/X VGND VGND VPWR
+ VPWR _17528_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33574_ _33702_/CLK _33574_/D VGND VGND VPWR VPWR _33574_/Q sky130_fd_sc_hd__dfxtp_1
X_30786_ _30786_/A VGND VGND VPWR VPWR _35621_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35313_ _35313_/CLK _35313_/D VGND VGND VPWR VPWR _35313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32525_ _36045_/CLK _32525_/D VGND VGND VPWR VPWR _32525_/Q sky130_fd_sc_hd__dfxtp_1
X_17459_ _17347_/X _17457_/X _17458_/X _17350_/X VGND VGND VPWR VPWR _17459_/X sky130_fd_sc_hd__a22o_1
XFILLER_220_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35244_ _35304_/CLK _35244_/D VGND VGND VPWR VPWR _35244_/Q sky130_fd_sc_hd__dfxtp_1
X_32456_ _35337_/CLK _32456_/D VGND VGND VPWR VPWR _32456_/Q sky130_fd_sc_hd__dfxtp_1
X_20470_ _35786_/Q _35146_/Q _34506_/Q _33866_/Q _18408_/X _18409_/X VGND VGND VPWR
+ VPWR _20470_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31407_ _31407_/A VGND VGND VPWR VPWR _35916_/D sky130_fd_sc_hd__clkbuf_1
X_19129_ _35555_/Q _35491_/Q _35427_/Q _35363_/Q _18844_/X _18845_/X VGND VGND VPWR
+ VPWR _19129_/X sky130_fd_sc_hd__mux4_1
X_35175_ _36005_/CLK _35175_/D VGND VGND VPWR VPWR _35175_/Q sky130_fd_sc_hd__dfxtp_1
X_32387_ _36037_/CLK _32387_/D VGND VGND VPWR VPWR _32387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34126_ _35021_/CLK _34126_/D VGND VGND VPWR VPWR _34126_/Q sky130_fd_sc_hd__dfxtp_1
X_22140_ _35319_/Q _35255_/Q _35191_/Q _32311_/Q _21959_/X _21960_/X VGND VGND VPWR
+ VPWR _22140_/X sky130_fd_sc_hd__mux4_1
XFILLER_146_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31338_ _31338_/A VGND VGND VPWR VPWR _35883_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34057_ _34057_/CLK _34057_/D VGND VGND VPWR VPWR _34057_/Q sky130_fd_sc_hd__dfxtp_1
X_22071_ _22071_/A _22071_/B _22071_/C _22071_/D VGND VGND VPWR VPWR _22072_/A sky130_fd_sc_hd__or4_4
XTAP_6709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31269_ _35851_/Q input58/X _31273_/S VGND VGND VPWR VPWR _31270_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21022_ _22434_/A VGND VGND VPWR VPWR _21022_/X sky130_fd_sc_hd__clkbuf_4
X_33008_ _33009_/CLK _33008_/D VGND VGND VPWR VPWR _33008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25830_ _25830_/A VGND VGND VPWR VPWR _33336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25761_ _25872_/S VGND VGND VPWR VPWR _25780_/S sky130_fd_sc_hd__buf_4
X_34959_ _35026_/CLK _34959_/D VGND VGND VPWR VPWR _34959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22973_ _23075_/S VGND VGND VPWR VPWR _23001_/S sky130_fd_sc_hd__buf_4
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24712_ _24712_/A VGND VGND VPWR VPWR _32843_/D sky130_fd_sc_hd__clkbuf_1
X_27500_ _27500_/A VGND VGND VPWR VPWR _34096_/D sky130_fd_sc_hd__clkbuf_1
X_28480_ _26977_/X _34560_/Q _28498_/S VGND VGND VPWR VPWR _28481_/A sky130_fd_sc_hd__mux2_1
X_21924_ _21749_/X _21922_/X _21923_/X _21752_/X VGND VGND VPWR VPWR _21924_/X sky130_fd_sc_hd__a22o_1
XFILLER_216_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25692_ _33272_/Q _24376_/X _25706_/S VGND VGND VPWR VPWR _25693_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27431_ _27431_/A VGND VGND VPWR VPWR _34063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24643_ _24643_/A VGND VGND VPWR VPWR _32810_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21855_ _21849_/X _21854_/X _21747_/X VGND VGND VPWR VPWR _21863_/C sky130_fd_sc_hd__o21ba_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20806_ _33746_/Q _33682_/Q _33618_/Q _33554_/Q _20737_/X _20738_/X VGND VGND VPWR
+ VPWR _20806_/X sky130_fd_sc_hd__mux4_1
X_27362_ _34031_/Q _24348_/X _27374_/S VGND VGND VPWR VPWR _27363_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24574_ _24574_/A VGND VGND VPWR VPWR _32779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21786_ _34797_/Q _34733_/Q _34669_/Q _34605_/Q _21535_/X _21536_/X VGND VGND VPWR
+ VPWR _21786_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29101_ input8/X VGND VGND VPWR VPWR _29101_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26313_ _26313_/A VGND VGND VPWR VPWR _33565_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23525_ _23525_/A VGND VGND VPWR VPWR _32316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27293_ _33998_/Q _24244_/X _27311_/S VGND VGND VPWR VPWR _27294_/A sky130_fd_sc_hd__mux2_1
X_20737_ _22502_/A VGND VGND VPWR VPWR _20737_/X sky130_fd_sc_hd__buf_6
XFILLER_196_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29032_ _34822_/Q _24419_/X _29038_/S VGND VGND VPWR VPWR _29033_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26244_ _25137_/X _33533_/Q _26248_/S VGND VGND VPWR VPWR _26245_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23456_ _23456_/A VGND VGND VPWR VPWR _32283_/D sky130_fd_sc_hd__clkbuf_1
X_20668_ _22465_/A VGND VGND VPWR VPWR _20668_/X sky130_fd_sc_hd__buf_4
XFILLER_184_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22407_ _33023_/Q _32959_/Q _32895_/Q _32831_/Q _22295_/X _22296_/X VGND VGND VPWR
+ VPWR _22407_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26175_ _25035_/X _33500_/Q _26185_/S VGND VGND VPWR VPWR _26176_/A sky130_fd_sc_hd__mux2_1
X_23387_ _23387_/A VGND VGND VPWR VPWR _32252_/D sky130_fd_sc_hd__clkbuf_1
X_20599_ _22396_/A VGND VGND VPWR VPWR _20599_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_136_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25126_ _25125_/X _33017_/Q _25144_/S VGND VGND VPWR VPWR _25127_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22338_ _35837_/Q _32216_/Q _35709_/Q _35645_/Q _22266_/X _22267_/X VGND VGND VPWR
+ VPWR _22338_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29934_ _35218_/Q _29064_/X _29944_/S VGND VGND VPWR VPWR _29935_/A sky130_fd_sc_hd__mux2_1
X_25057_ input14/X VGND VGND VPWR VPWR _25057_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_151_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22269_ _35771_/Q _35131_/Q _34491_/Q _33851_/Q _22093_/X _22094_/X VGND VGND VPWR
+ VPWR _22269_/X sky130_fd_sc_hd__mux4_1
X_24008_ _22929_/X _32542_/Q _24014_/S VGND VGND VPWR VPWR _24009_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29865_ _29865_/A VGND VGND VPWR VPWR _35185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16830_ _33187_/Q _32547_/Q _35939_/Q _35875_/Q _16721_/X _16722_/X VGND VGND VPWR
+ VPWR _16830_/X sky130_fd_sc_hd__mux4_1
X_28816_ _28816_/A VGND VGND VPWR VPWR _34719_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29796_ _29796_/A VGND VGND VPWR VPWR _35152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28747_ _26974_/X _34687_/Q _28747_/S VGND VGND VPWR VPWR _28748_/A sky130_fd_sc_hd__mux2_1
X_16761_ _34529_/Q _32417_/Q _34401_/Q _34337_/Q _16519_/X _16520_/X VGND VGND VPWR
+ VPWR _16761_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25959_ _26007_/S VGND VGND VPWR VPWR _25978_/S sky130_fd_sc_hd__buf_4
XFILLER_4_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18500_ _34513_/Q _32401_/Q _34385_/Q _34321_/Q _18466_/X _18467_/X VGND VGND VPWR
+ VPWR _18500_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_1183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19480_ _35757_/Q _35117_/Q _34477_/Q _33837_/Q _19440_/X _19441_/X VGND VGND VPWR
+ VPWR _19480_/X sky130_fd_sc_hd__mux4_1
X_16692_ _16688_/X _16691_/X _16455_/X VGND VGND VPWR VPWR _16693_/D sky130_fd_sc_hd__o21ba_1
XFILLER_234_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28678_ _26872_/X _34654_/Q _28684_/S VGND VGND VPWR VPWR _28679_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18431_ _35023_/Q _34959_/Q _34895_/Q _34831_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _18431_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27629_ _27629_/A VGND VGND VPWR VPWR _34156_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30640_ _30640_/A VGND VGND VPWR VPWR _35552_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18362_ _20278_/A VGND VGND VPWR VPWR _20231_/A sky130_fd_sc_hd__buf_12
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17313_ _17795_/A VGND VGND VPWR VPWR _17313_/X sky130_fd_sc_hd__buf_6
X_30571_ _30598_/S VGND VGND VPWR VPWR _30590_/S sky130_fd_sc_hd__buf_4
XFILLER_25_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18293_ _18277_/X _18284_/X _18287_/X _18292_/X VGND VGND VPWR VPWR _18293_/X sky130_fd_sc_hd__a22o_1
XFILLER_109_1074 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32310_ _35318_/CLK _32310_/D VGND VGND VPWR VPWR _32310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17244_ _33007_/Q _32943_/Q _32879_/Q _32815_/Q _16989_/X _16990_/X VGND VGND VPWR
+ VPWR _17244_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33290_ _36172_/CLK _33290_/D VGND VGND VPWR VPWR _33290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17175_ _32493_/Q _32365_/Q _32045_/Q _36013_/Q _16923_/X _17064_/X VGND VGND VPWR
+ VPWR _17175_/X sky130_fd_sc_hd__mux4_1
X_32241_ _34032_/CLK _32241_/D VGND VGND VPWR VPWR _32241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16126_ _16122_/X _16125_/X _16071_/X VGND VGND VPWR VPWR _16134_/C sky130_fd_sc_hd__o21ba_1
X_32172_ _35669_/CLK _32172_/D VGND VGND VPWR VPWR _32172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31123_ _31123_/A VGND VGND VPWR VPWR _35781_/D sky130_fd_sc_hd__clkbuf_1
X_16057_ _16057_/A VGND VGND VPWR VPWR _17846_/A sky130_fd_sc_hd__buf_12
XFILLER_170_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31054_ _31054_/A VGND VGND VPWR VPWR _35748_/D sky130_fd_sc_hd__clkbuf_1
X_35931_ _35931_/CLK _35931_/D VGND VGND VPWR VPWR _35931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30005_ _35252_/Q _29169_/X _30007_/S VGND VGND VPWR VPWR _30006_/A sky130_fd_sc_hd__mux2_1
X_19816_ _19816_/A _19816_/B _19816_/C _19816_/D VGND VGND VPWR VPWR _19817_/A sky130_fd_sc_hd__or4_4
X_35862_ _36118_/CLK _35862_/D VGND VGND VPWR VPWR _35862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34813_ _36028_/CLK _34813_/D VGND VGND VPWR VPWR _34813_/Q sky130_fd_sc_hd__dfxtp_1
X_19747_ _34037_/Q _33973_/Q _33909_/Q _32245_/Q _19673_/X _19674_/X VGND VGND VPWR
+ VPWR _19747_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35793_ _35793_/CLK _35793_/D VGND VGND VPWR VPWR _35793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16959_ _16955_/X _16958_/X _16783_/X _16784_/X VGND VGND VPWR VPWR _16976_/B sky130_fd_sc_hd__o211a_1
XFILLER_244_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34744_ _35318_/CLK _34744_/D VGND VGND VPWR VPWR _34744_/Q sky130_fd_sc_hd__dfxtp_1
X_31956_ _35036_/CLK _31956_/D VGND VGND VPWR VPWR _31956_/Q sky130_fd_sc_hd__dfxtp_1
X_19678_ _32755_/Q _32691_/Q _32627_/Q _36083_/Q _19572_/X _19356_/X VGND VGND VPWR
+ VPWR _19678_/X sky130_fd_sc_hd__mux4_1
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18629_ _35541_/Q _35477_/Q _35413_/Q _35349_/Q _18491_/X _18492_/X VGND VGND VPWR
+ VPWR _18629_/X sky130_fd_sc_hd__mux4_1
X_30907_ _35679_/Q _29104_/X _30911_/S VGND VGND VPWR VPWR _30908_/A sky130_fd_sc_hd__mux2_1
X_34675_ _35242_/CLK _34675_/D VGND VGND VPWR VPWR _34675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31887_ _31887_/A VGND VGND VPWR VPWR _36143_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21640_ _35305_/Q _35241_/Q _35177_/Q _32297_/Q _21606_/X _21607_/X VGND VGND VPWR
+ VPWR _21640_/X sky130_fd_sc_hd__mux4_1
X_33626_ _33692_/CLK _33626_/D VGND VGND VPWR VPWR _33626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30838_ _30838_/A VGND VGND VPWR VPWR _35646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1084 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33557_ _33685_/CLK _33557_/D VGND VGND VPWR VPWR _33557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21571_ _21396_/X _21569_/X _21570_/X _21399_/X VGND VGND VPWR VPWR _21571_/X sky130_fd_sc_hd__a22o_1
X_30769_ _30769_/A VGND VGND VPWR VPWR _35613_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_11 _32114_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _32115_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23310_ input48/X VGND VGND VPWR VPWR _23310_/X sky130_fd_sc_hd__buf_4
X_20522_ _32780_/Q _32716_/Q _32652_/Q _36108_/Q _20278_/X _19173_/A VGND VGND VPWR
+ VPWR _20522_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32508_ _36028_/CLK _32508_/D VGND VGND VPWR VPWR _32508_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_33 _32117_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_44 _32118_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24290_ _32668_/Q _24289_/X _24305_/S VGND VGND VPWR VPWR _24291_/A sky130_fd_sc_hd__mux2_1
X_33488_ _33940_/CLK _33488_/D VGND VGND VPWR VPWR _33488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_55 _32126_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_66 _32126_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_77 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23241_ input25/X VGND VGND VPWR VPWR _23241_/X sky130_fd_sc_hd__buf_4
X_35227_ _36201_/CLK _35227_/D VGND VGND VPWR VPWR _35227_/Q sky130_fd_sc_hd__dfxtp_1
X_20453_ _20453_/A _20453_/B _20453_/C _20453_/D VGND VGND VPWR VPWR _20454_/A sky130_fd_sc_hd__or4_1
XANTENNA_88 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32439_ _35319_/CLK _32439_/D VGND VGND VPWR VPWR _32439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_99 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23172_ _23172_/A VGND VGND VPWR VPWR _32169_/D sky130_fd_sc_hd__clkbuf_1
X_35158_ _35286_/CLK _35158_/D VGND VGND VPWR VPWR _35158_/Q sky130_fd_sc_hd__dfxtp_1
X_20384_ _18297_/X _20382_/X _20383_/X _18303_/X VGND VGND VPWR VPWR _20384_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34109_ _36157_/CLK _34109_/D VGND VGND VPWR VPWR _34109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22123_ _21802_/X _22121_/X _22122_/X _21805_/X VGND VGND VPWR VPWR _22123_/X sky130_fd_sc_hd__a22o_1
XFILLER_216_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35089_ _35729_/CLK _35089_/D VGND VGND VPWR VPWR _35089_/Q sky130_fd_sc_hd__dfxtp_1
X_27980_ _26838_/X _34323_/Q _27988_/S VGND VGND VPWR VPWR _27981_/A sky130_fd_sc_hd__mux2_1
Xoutput140 _32005_/Q VGND VGND VPWR VPWR D1[55] sky130_fd_sc_hd__buf_2
XTAP_6506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput151 _31957_/Q VGND VGND VPWR VPWR D1[7] sky130_fd_sc_hd__buf_2
XTAP_6517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput162 _36191_/Q VGND VGND VPWR VPWR D2[17] sky130_fd_sc_hd__buf_2
XFILLER_217_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput173 _36201_/Q VGND VGND VPWR VPWR D2[27] sky130_fd_sc_hd__buf_2
XFILLER_134_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26931_ input29/X VGND VGND VPWR VPWR _26931_/X sky130_fd_sc_hd__buf_4
X_22054_ _33013_/Q _32949_/Q _32885_/Q _32821_/Q _21942_/X _21943_/X VGND VGND VPWR
+ VPWR _22054_/X sky130_fd_sc_hd__mux4_1
XFILLER_248_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput184 _36211_/Q VGND VGND VPWR VPWR D2[37] sky130_fd_sc_hd__buf_2
Xoutput195 _36221_/Q VGND VGND VPWR VPWR D2[47] sky130_fd_sc_hd__buf_2
XTAP_5805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21005_ _34775_/Q _34711_/Q _34647_/Q _34583_/Q _20829_/X _20830_/X VGND VGND VPWR
+ VPWR _21005_/X sky130_fd_sc_hd__mux4_1
XFILLER_247_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29650_ _35084_/Q _29243_/X _29652_/S VGND VGND VPWR VPWR _29651_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1028 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26862_ _26862_/A VGND VGND VPWR VPWR _33818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28601_ _28601_/A VGND VGND VPWR VPWR _34617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25813_ _25813_/A VGND VGND VPWR VPWR _33328_/D sky130_fd_sc_hd__clkbuf_1
X_26793_ _33792_/Q _24400_/X _26811_/S VGND VGND VPWR VPWR _26794_/A sky130_fd_sc_hd__mux2_1
X_29581_ _35051_/Q _29141_/X _29581_/S VGND VGND VPWR VPWR _29582_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25744_ _25744_/A VGND VGND VPWR VPWR _33295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28532_ _28532_/A VGND VGND VPWR VPWR _34584_/D sky130_fd_sc_hd__clkbuf_1
X_22956_ _22956_/A VGND VGND VPWR VPWR _32038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21907_ _33265_/Q _36145_/Q _33137_/Q _33073_/Q _21658_/X _21659_/X VGND VGND VPWR
+ VPWR _21907_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28463_ _26953_/X _34552_/Q _28477_/S VGND VGND VPWR VPWR _28464_/A sky130_fd_sc_hd__mux2_1
X_25675_ _33264_/Q _24351_/X _25685_/S VGND VGND VPWR VPWR _25676_/A sky130_fd_sc_hd__mux2_1
X_22887_ _22886_/X _32016_/Q _22908_/S VGND VGND VPWR VPWR _22888_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27414_ _34056_/Q _24425_/X _27416_/S VGND VGND VPWR VPWR _27415_/A sky130_fd_sc_hd__mux2_1
X_24626_ _22941_/X _32802_/Q _24644_/S VGND VGND VPWR VPWR _24627_/A sky130_fd_sc_hd__mux2_1
X_28394_ _28394_/A VGND VGND VPWR VPWR _34519_/D sky130_fd_sc_hd__clkbuf_1
X_21838_ _21802_/X _21836_/X _21837_/X _21805_/X VGND VGND VPWR VPWR _21838_/X sky130_fd_sc_hd__a22o_1
XFILLER_231_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27345_ _34023_/Q _24323_/X _27353_/S VGND VGND VPWR VPWR _27346_/A sky130_fd_sc_hd__mux2_1
X_24557_ _23044_/X _32771_/Q _24569_/S VGND VGND VPWR VPWR _24558_/A sky130_fd_sc_hd__mux2_1
X_21769_ _34029_/Q _33965_/Q _33901_/Q _32237_/Q _21620_/X _21621_/X VGND VGND VPWR
+ VPWR _21769_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23508_ _23508_/A VGND VGND VPWR VPWR _32308_/D sky130_fd_sc_hd__clkbuf_1
X_27276_ _27276_/A VGND VGND VPWR VPWR _33990_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24488_ _22941_/X _32738_/Q _24506_/S VGND VGND VPWR VPWR _24489_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29015_ _34814_/Q _24394_/X _29017_/S VGND VGND VPWR VPWR _29016_/A sky130_fd_sc_hd__mux2_1
X_26227_ _25112_/X _33525_/Q _26227_/S VGND VGND VPWR VPWR _26228_/A sky130_fd_sc_hd__mux2_1
X_23439_ _23439_/A VGND VGND VPWR VPWR _32275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26158_ _25010_/X _33492_/Q _26164_/S VGND VGND VPWR VPWR _26159_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25109_ input32/X VGND VGND VPWR VPWR _25109_/X sky130_fd_sc_hd__buf_2
XFILLER_152_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18980_ _35743_/Q _35103_/Q _34463_/Q _33823_/Q _18734_/X _18735_/X VGND VGND VPWR
+ VPWR _18980_/X sky130_fd_sc_hd__mux4_1
X_26089_ _26089_/A VGND VGND VPWR VPWR _33459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29917_ _29917_/A VGND VGND VPWR VPWR _35210_/D sky130_fd_sc_hd__clkbuf_1
X_17931_ _17931_/A VGND VGND VPWR VPWR _17931_/X sky130_fd_sc_hd__buf_6
XFILLER_112_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17862_ _17862_/A VGND VGND VPWR VPWR _17862_/X sky130_fd_sc_hd__buf_4
X_29848_ _29848_/A VGND VGND VPWR VPWR _35177_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19601_ _19495_/X _19599_/X _19600_/X _19500_/X VGND VGND VPWR VPWR _19601_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16813_ _34275_/Q _34211_/Q _34147_/Q _34083_/Q _16736_/X _16737_/X VGND VGND VPWR
+ VPWR _16813_/X sky130_fd_sc_hd__mux4_1
X_29779_ _35145_/Q _29234_/X _29779_/S VGND VGND VPWR VPWR _29780_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17793_ _17793_/A VGND VGND VPWR VPWR _31998_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_213_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31810_ _31810_/A VGND VGND VPWR VPWR _36107_/D sky130_fd_sc_hd__clkbuf_1
X_19532_ _19532_/A VGND VGND VPWR VPWR _32110_/D sky130_fd_sc_hd__buf_2
X_16744_ _32737_/Q _32673_/Q _32609_/Q _36065_/Q _16566_/X _16703_/X VGND VGND VPWR
+ VPWR _16744_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32790_ _36116_/CLK _32790_/D VGND VGND VPWR VPWR _32790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19463_ _19463_/A _19463_/B _19463_/C _19463_/D VGND VGND VPWR VPWR _19464_/A sky130_fd_sc_hd__or4_1
XFILLER_62_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31741_ _31741_/A VGND VGND VPWR VPWR _36074_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16675_ _32479_/Q _32351_/Q _32031_/Q _35999_/Q _16570_/X _16358_/X VGND VGND VPWR
+ VPWR _16675_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18414_ _33231_/Q _36111_/Q _33103_/Q _33039_/Q _18320_/X _18321_/X VGND VGND VPWR
+ VPWR _18414_/X sky130_fd_sc_hd__mux4_1
X_34460_ _35738_/CLK _34460_/D VGND VGND VPWR VPWR _34460_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31672_ _36042_/Q input57/X _31678_/S VGND VGND VPWR VPWR _31673_/A sky130_fd_sc_hd__mux2_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19394_ _34027_/Q _33963_/Q _33899_/Q _32235_/Q _19320_/X _19321_/X VGND VGND VPWR
+ VPWR _19394_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33411_ _33545_/CLK _33411_/D VGND VGND VPWR VPWR _33411_/Q sky130_fd_sc_hd__dfxtp_1
X_18345_ _20095_/A VGND VGND VPWR VPWR _18345_/X sky130_fd_sc_hd__buf_8
X_30623_ _35544_/Q _29082_/X _30641_/S VGND VGND VPWR VPWR _30624_/A sky130_fd_sc_hd__mux2_1
X_34391_ _36196_/CLK _34391_/D VGND VGND VPWR VPWR _34391_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36130_ _36130_/CLK _36130_/D VGND VGND VPWR VPWR _36130_/Q sky130_fd_sc_hd__dfxtp_1
X_33342_ _34302_/CLK _33342_/D VGND VGND VPWR VPWR _33342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18276_ _20061_/A VGND VGND VPWR VPWR _20155_/A sky130_fd_sc_hd__buf_12
X_30554_ _30554_/A VGND VGND VPWR VPWR _35511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput20 DW[27] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__buf_4
X_17227_ _34542_/Q _32430_/Q _34414_/Q _34350_/Q _17225_/X _17226_/X VGND VGND VPWR
+ VPWR _17227_/X sky130_fd_sc_hd__mux4_1
X_36061_ _36127_/CLK _36061_/D VGND VGND VPWR VPWR _36061_/Q sky130_fd_sc_hd__dfxtp_1
X_33273_ _36088_/CLK _33273_/D VGND VGND VPWR VPWR _33273_/Q sky130_fd_sc_hd__dfxtp_1
Xinput31 DW[37] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_4
XFILLER_239_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30485_ _23114_/X _35479_/Q _30485_/S VGND VGND VPWR VPWR _30486_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput42 DW[47] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__buf_6
X_35012_ _35779_/CLK _35012_/D VGND VGND VPWR VPWR _35012_/Q sky130_fd_sc_hd__dfxtp_1
Xinput53 DW[57] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_16
X_32224_ _35845_/CLK _32224_/D VGND VGND VPWR VPWR _32224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput64 DW[9] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__buf_8
Xinput75 R2[4] VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__buf_2
XFILLER_122_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17158_ _35052_/Q _34988_/Q _34924_/Q _34860_/Q _17156_/X _17157_/X VGND VGND VPWR
+ VPWR _17158_/X sky130_fd_sc_hd__mux4_1
Xinput86 RW[3] VGND VGND VPWR VPWR input86/X sky130_fd_sc_hd__buf_2
XFILLER_196_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16109_ _17847_/A VGND VGND VPWR VPWR _16109_/X sky130_fd_sc_hd__buf_4
XFILLER_196_1183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32155_ _34202_/CLK _32155_/D VGND VGND VPWR VPWR _32155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17089_ _17956_/A VGND VGND VPWR VPWR _17089_/X sky130_fd_sc_hd__buf_6
XFILLER_115_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31106_ _31106_/A VGND VGND VPWR VPWR _35773_/D sky130_fd_sc_hd__clkbuf_1
X_32086_ _35040_/CLK _32086_/D VGND VGND VPWR VPWR _32086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35914_ _35978_/CLK _35914_/D VGND VGND VPWR VPWR _35914_/Q sky130_fd_sc_hd__dfxtp_1
X_31037_ _31037_/A VGND VGND VPWR VPWR _35740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35845_ _35845_/CLK _35845_/D VGND VGND VPWR VPWR _35845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22810_ _35083_/Q _35019_/Q _34955_/Q _34891_/Q _20679_/X _20681_/X VGND VGND VPWR
+ VPWR _22810_/X sky130_fd_sc_hd__mux4_1
X_35776_ _35777_/CLK _35776_/D VGND VGND VPWR VPWR _35776_/Q sky130_fd_sc_hd__dfxtp_1
X_23790_ _23790_/A VGND VGND VPWR VPWR _32439_/D sky130_fd_sc_hd__clkbuf_1
X_32988_ _33244_/CLK _32988_/D VGND VGND VPWR VPWR _32988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22741_ _20577_/X _22739_/X _22740_/X _20587_/X VGND VGND VPWR VPWR _22741_/X sky130_fd_sc_hd__a22o_1
X_34727_ _34792_/CLK _34727_/D VGND VGND VPWR VPWR _34727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_812 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31939_ _31939_/A VGND VGND VPWR VPWR _36168_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25460_ _30329_/A _30329_/B _29049_/B VGND VGND VPWR VPWR _25461_/A sky130_fd_sc_hd__or3_1
X_22672_ _32775_/Q _32711_/Q _32647_/Q _36103_/Q _22578_/X _22362_/X VGND VGND VPWR
+ VPWR _22672_/X sky130_fd_sc_hd__mux4_1
X_34658_ _35928_/CLK _34658_/D VGND VGND VPWR VPWR _34658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24411_ _32707_/Q _24410_/X _24429_/S VGND VGND VPWR VPWR _24412_/A sky130_fd_sc_hd__mux2_1
X_33609_ _34817_/CLK _33609_/D VGND VGND VPWR VPWR _33609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21623_ _21449_/X _21619_/X _21622_/X _21452_/X VGND VGND VPWR VPWR _21623_/X sky130_fd_sc_hd__a22o_1
XFILLER_240_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25391_ _25391_/A VGND VGND VPWR VPWR _33132_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34589_ _35034_/CLK _34589_/D VGND VGND VPWR VPWR _34589_/Q sky130_fd_sc_hd__dfxtp_1
X_27130_ _26981_/X _33921_/Q _27146_/S VGND VGND VPWR VPWR _27131_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24342_ input25/X VGND VGND VPWR VPWR _24342_/X sky130_fd_sc_hd__buf_6
XFILLER_21_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21554_ _33255_/Q _36135_/Q _33127_/Q _33063_/Q _21305_/X _21306_/X VGND VGND VPWR
+ VPWR _21554_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20505_ _20501_/X _20504_/X _20153_/A VGND VGND VPWR VPWR _20513_/C sky130_fd_sc_hd__o21ba_1
XFILLER_154_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27061_ _27061_/A VGND VGND VPWR VPWR _33888_/D sky130_fd_sc_hd__clkbuf_1
X_24273_ input64/X VGND VGND VPWR VPWR _24273_/X sky130_fd_sc_hd__clkbuf_8
X_21485_ _21449_/X _21483_/X _21484_/X _21452_/X VGND VGND VPWR VPWR _21485_/X sky130_fd_sc_hd__a22o_1
XFILLER_222_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26012_ _26012_/A VGND VGND VPWR VPWR _33422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23224_ _32192_/Q _23223_/X _23235_/S VGND VGND VPWR VPWR _23225_/A sky130_fd_sc_hd__mux2_1
X_20436_ _33033_/Q _32969_/Q _32905_/Q _32841_/Q _18280_/X _18283_/X VGND VGND VPWR
+ VPWR _20436_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23155_ _30329_/A _30329_/B _29049_/B VGND VGND VPWR VPWR _23156_/A sky130_fd_sc_hd__or3b_1
XFILLER_134_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20367_ _20201_/X _20365_/X _20366_/X _20206_/X VGND VGND VPWR VPWR _20367_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22106_ _22102_/X _22103_/X _22104_/X _22105_/X VGND VGND VPWR VPWR _22106_/X sky130_fd_sc_hd__a22o_1
XTAP_7059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27963_ _27963_/A VGND VGND VPWR VPWR _34315_/D sky130_fd_sc_hd__clkbuf_1
X_23086_ _27833_/A _31275_/A VGND VGND VPWR VPWR _23421_/S sky130_fd_sc_hd__nor2_8
XANTENNA_1109 _36201_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20298_ _20155_/X _20296_/X _20297_/X _20158_/X VGND VGND VPWR VPWR _20298_/X sky130_fd_sc_hd__a22o_1
XTAP_6336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29702_ _35108_/Q _29120_/X _29716_/S VGND VGND VPWR VPWR _29703_/A sky130_fd_sc_hd__mux2_1
XTAP_6358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26914_ _26914_/A VGND VGND VPWR VPWR _33835_/D sky130_fd_sc_hd__clkbuf_1
X_22037_ _21754_/X _22035_/X _22036_/X _21759_/X VGND VGND VPWR VPWR _22037_/X sky130_fd_sc_hd__a22o_1
XTAP_6369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27894_ _27894_/A VGND VGND VPWR VPWR _34282_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29633_ _29633_/A VGND VGND VPWR VPWR _35075_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26845_ _26844_/X _33813_/Q _26851_/S VGND VGND VPWR VPWR _26846_/A sky130_fd_sc_hd__mux2_1
XTAP_5679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29564_ _29564_/A VGND VGND VPWR VPWR _35042_/D sky130_fd_sc_hd__clkbuf_1
X_23988_ _23988_/A VGND VGND VPWR VPWR _32532_/D sky130_fd_sc_hd__clkbuf_1
X_26776_ _33784_/Q _24376_/X _26790_/S VGND VGND VPWR VPWR _26777_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28515_ _28515_/A VGND VGND VPWR VPWR _34576_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25727_ _33289_/Q _24428_/X _25727_/S VGND VGND VPWR VPWR _25728_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22939_ _22938_/X _32033_/Q _22939_/S VGND VGND VPWR VPWR _22940_/A sky130_fd_sc_hd__mux2_1
X_29495_ _23310_/X _35010_/Q _29509_/S VGND VGND VPWR VPWR _29496_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16460_ _34265_/Q _34201_/Q _34137_/Q _34073_/Q _16383_/X _16384_/X VGND VGND VPWR
+ VPWR _16460_/X sky130_fd_sc_hd__mux4_1
X_28446_ _26928_/X _34544_/Q _28456_/S VGND VGND VPWR VPWR _28447_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25658_ _33256_/Q _24326_/X _25664_/S VGND VGND VPWR VPWR _25659_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16391_ _32727_/Q _32663_/Q _32599_/Q _36055_/Q _16213_/X _16350_/X VGND VGND VPWR
+ VPWR _16391_/X sky130_fd_sc_hd__mux4_1
X_24609_ _22917_/X _32794_/Q _24623_/S VGND VGND VPWR VPWR _24610_/A sky130_fd_sc_hd__mux2_1
XPHY_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25589_ _33225_/Q _24428_/X _25589_/S VGND VGND VPWR VPWR _25590_/A sky130_fd_sc_hd__mux2_1
X_28377_ _26826_/X _34511_/Q _28393_/S VGND VGND VPWR VPWR _28378_/A sky130_fd_sc_hd__mux2_1
XPHY_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18130_ _17908_/X _18128_/X _18129_/X _17911_/X VGND VGND VPWR VPWR _18130_/X sky130_fd_sc_hd__a22o_1
XPHY_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27328_ _34015_/Q _24298_/X _27332_/S VGND VGND VPWR VPWR _27329_/A sky130_fd_sc_hd__mux2_1
XPHY_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18061_ _17860_/X _18059_/X _18060_/X _17865_/X VGND VGND VPWR VPWR _18061_/X sky130_fd_sc_hd__a22o_1
X_27259_ _27259_/A VGND VGND VPWR VPWR _33982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17012_ _16801_/X _17010_/X _17011_/X _16806_/X VGND VGND VPWR VPWR _17012_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30270_ _30270_/A VGND VGND VPWR VPWR _35377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_180_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _35982_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_113_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18963_ _33759_/Q _33695_/Q _33631_/Q _33567_/Q _18790_/X _18791_/X VGND VGND VPWR
+ VPWR _18963_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17914_ _32770_/Q _32706_/Q _32642_/Q _36098_/Q _17625_/X _17762_/X VGND VGND VPWR
+ VPWR _17914_/X sky130_fd_sc_hd__mux4_1
X_33960_ _34153_/CLK _33960_/D VGND VGND VPWR VPWR _33960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18894_ _34269_/Q _34205_/Q _34141_/Q _34077_/Q _18683_/X _18684_/X VGND VGND VPWR
+ VPWR _18894_/X sky130_fd_sc_hd__mux4_1
XTAP_6870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32911_ _35985_/CLK _32911_/D VGND VGND VPWR VPWR _32911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17845_ _35840_/Q _32219_/Q _35712_/Q _35648_/Q _17666_/X _17667_/X VGND VGND VPWR
+ VPWR _17845_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33891_ _36130_/CLK _33891_/D VGND VGND VPWR VPWR _33891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35630_ _35822_/CLK _35630_/D VGND VGND VPWR VPWR _35630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32842_ _35979_/CLK _32842_/D VGND VGND VPWR VPWR _32842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17776_ _35838_/Q _32217_/Q _35710_/Q _35646_/Q _17666_/X _17667_/X VGND VGND VPWR
+ VPWR _17776_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_1411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19515_ _35822_/Q _32199_/Q _35694_/Q _35630_/Q _19260_/X _19261_/X VGND VGND VPWR
+ VPWR _19515_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35561_ _35562_/CLK _35561_/D VGND VGND VPWR VPWR _35561_/Q sky130_fd_sc_hd__dfxtp_1
X_16727_ _35296_/Q _35232_/Q _35168_/Q _32288_/Q _16653_/X _16654_/X VGND VGND VPWR
+ VPWR _16727_/X sky130_fd_sc_hd__mux4_1
X_32773_ _36103_/CLK _32773_/D VGND VGND VPWR VPWR _32773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34512_ _35281_/CLK _34512_/D VGND VGND VPWR VPWR _34512_/Q sky130_fd_sc_hd__dfxtp_1
X_19446_ _19299_/X _19444_/X _19445_/X _19302_/X VGND VGND VPWR VPWR _19446_/X sky130_fd_sc_hd__a22o_1
X_31724_ _36066_/Q input13/X _31742_/S VGND VGND VPWR VPWR _31725_/A sky130_fd_sc_hd__mux2_1
X_16658_ _35038_/Q _34974_/Q _34910_/Q _34846_/Q _16450_/X _16451_/X VGND VGND VPWR
+ VPWR _16658_/X sky130_fd_sc_hd__mux4_1
X_35492_ _35555_/CLK _35492_/D VGND VGND VPWR VPWR _35492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34443_ _35147_/CLK _34443_/D VGND VGND VPWR VPWR _34443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31655_ _31655_/A VGND VGND VPWR VPWR _36033_/D sky130_fd_sc_hd__clkbuf_1
X_19377_ _19299_/X _19373_/X _19376_/X _19302_/X VGND VGND VPWR VPWR _19377_/X sky130_fd_sc_hd__a22o_1
X_16589_ _16448_/X _16587_/X _16588_/X _16453_/X VGND VGND VPWR VPWR _16589_/X sky130_fd_sc_hd__a22o_1
XFILLER_245_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_1122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30606_ _35536_/Q _29058_/X _30620_/S VGND VGND VPWR VPWR _30607_/A sky130_fd_sc_hd__mux2_1
X_18328_ _20282_/A VGND VGND VPWR VPWR _18328_/X sky130_fd_sc_hd__buf_6
X_34374_ _35078_/CLK _34374_/D VGND VGND VPWR VPWR _34374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31586_ _36001_/Q input11/X _31586_/S VGND VGND VPWR VPWR _31587_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_6_36__f_CLK clkbuf_5_18_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_36__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_176_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36113_ _36114_/CLK _36113_/D VGND VGND VPWR VPWR _36113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33325_ _34293_/CLK _33325_/D VGND VGND VPWR VPWR _33325_/Q sky130_fd_sc_hd__dfxtp_1
X_18259_ _35853_/Q _32233_/Q _35725_/Q _35661_/Q _15989_/X _15991_/X VGND VGND VPWR
+ VPWR _18259_/X sky130_fd_sc_hd__mux4_1
X_30537_ _30537_/A VGND VGND VPWR VPWR _35503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36044_ _36045_/CLK _36044_/D VGND VGND VPWR VPWR _36044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33256_ _36136_/CLK _33256_/D VGND VGND VPWR VPWR _33256_/Q sky130_fd_sc_hd__dfxtp_1
X_21270_ _21096_/X _21266_/X _21269_/X _21099_/X VGND VGND VPWR VPWR _21270_/X sky130_fd_sc_hd__a22o_1
XFILLER_198_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30468_ _30468_/A VGND VGND VPWR VPWR _35470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20221_ _35842_/Q _32221_/Q _35714_/Q _35650_/Q _19966_/X _19967_/X VGND VGND VPWR
+ VPWR _20221_/X sky130_fd_sc_hd__mux4_1
X_32207_ _35828_/CLK _32207_/D VGND VGND VPWR VPWR _32207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_171_CLK clkbuf_leaf_76_CLK/A VGND VGND VPWR VPWR _34124_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_171_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33187_ _35938_/CLK _33187_/D VGND VGND VPWR VPWR _33187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30399_ _23244_/X _35438_/Q _30413_/S VGND VGND VPWR VPWR _30400_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20152_ _20005_/X _20150_/X _20151_/X _20008_/X VGND VGND VPWR VPWR _20152_/X sky130_fd_sc_hd__a22o_1
X_32138_ _35815_/CLK _32138_/D VGND VGND VPWR VPWR _32138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24960_ _24987_/S VGND VGND VPWR VPWR _24979_/S sky130_fd_sc_hd__buf_6
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32069_ _36037_/CLK _32069_/D VGND VGND VPWR VPWR _32069_/Q sky130_fd_sc_hd__dfxtp_1
X_20083_ _20005_/X _20079_/X _20082_/X _20008_/X VGND VGND VPWR VPWR _20083_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23911_ _23911_/A VGND VGND VPWR VPWR _32496_/D sky130_fd_sc_hd__clkbuf_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24891_ _22932_/X _32927_/Q _24895_/S VGND VGND VPWR VPWR _24892_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23842_ _23842_/A VGND VGND VPWR VPWR _32463_/D sky130_fd_sc_hd__clkbuf_1
X_26630_ _26630_/A VGND VGND VPWR VPWR _33715_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35828_ _35828_/CLK _35828_/D VGND VGND VPWR VPWR _35828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_507 _17900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26561_ _26561_/A VGND VGND VPWR VPWR _33682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_518 _17970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23773_ _23773_/A VGND VGND VPWR VPWR _32431_/D sky130_fd_sc_hd__clkbuf_1
X_35759_ _35760_/CLK _35759_/D VGND VGND VPWR VPWR _35759_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_529 _18154_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20985_ _34263_/Q _34199_/Q _34135_/Q _34071_/Q _20983_/X _20984_/X VGND VGND VPWR
+ VPWR _20985_/X sky130_fd_sc_hd__mux4_2
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28300_ _34475_/Q _24335_/X _28300_/S VGND VGND VPWR VPWR _28301_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22724_ _22724_/A VGND VGND VPWR VPWR _36232_/D sky130_fd_sc_hd__clkbuf_1
X_25512_ _33188_/Q _24314_/X _25526_/S VGND VGND VPWR VPWR _25513_/A sky130_fd_sc_hd__mux2_1
X_29280_ _23130_/X _34908_/Q _29290_/S VGND VGND VPWR VPWR _29281_/A sky130_fd_sc_hd__mux2_1
X_26492_ _26492_/A VGND VGND VPWR VPWR _33650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_1279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28231_ _28231_/A VGND VGND VPWR VPWR _34442_/D sky130_fd_sc_hd__clkbuf_1
X_25443_ _25443_/A VGND VGND VPWR VPWR _33157_/D sky130_fd_sc_hd__clkbuf_1
X_22655_ _22651_/X _22654_/X _22453_/X VGND VGND VPWR VPWR _22663_/C sky130_fd_sc_hd__o21ba_1
XFILLER_129_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21606_ _22312_/A VGND VGND VPWR VPWR _21606_/X sky130_fd_sc_hd__buf_4
XFILLER_199_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28162_ _28162_/A VGND VGND VPWR VPWR _34409_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25374_ _25374_/A VGND VGND VPWR VPWR _33124_/D sky130_fd_sc_hd__clkbuf_1
X_22586_ _22581_/X _22585_/X _22442_/X _22443_/X VGND VGND VPWR VPWR _22603_/B sky130_fd_sc_hd__o211a_1
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27113_ _26956_/X _33913_/Q _27125_/S VGND VGND VPWR VPWR _27114_/A sky130_fd_sc_hd__mux2_1
X_24325_ _24325_/A VGND VGND VPWR VPWR _32679_/D sky130_fd_sc_hd__clkbuf_1
X_28093_ _27005_/X _34377_/Q _28093_/S VGND VGND VPWR VPWR _28094_/A sky130_fd_sc_hd__mux2_1
X_21537_ _34790_/Q _34726_/Q _34662_/Q _34598_/Q _21535_/X _21536_/X VGND VGND VPWR
+ VPWR _21537_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27044_ _26853_/X _33880_/Q _27062_/S VGND VGND VPWR VPWR _27045_/A sky130_fd_sc_hd__mux2_1
X_24256_ _32657_/Q _24255_/X _24274_/S VGND VGND VPWR VPWR _24257_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_958 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21468_ _21464_/X _21467_/X _21394_/X VGND VGND VPWR VPWR _21478_/C sky130_fd_sc_hd__o21ba_1
X_23207_ _23207_/A VGND VGND VPWR VPWR _32185_/D sky130_fd_sc_hd__clkbuf_1
X_20419_ _34568_/Q _32456_/Q _34440_/Q _34376_/Q _20231_/X _20232_/X VGND VGND VPWR
+ VPWR _20419_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_162_CLK clkbuf_6_30__f_CLK/X VGND VGND VPWR VPWR _36171_/CLK sky130_fd_sc_hd__clkbuf_16
X_24187_ _24187_/A VGND VGND VPWR VPWR _32626_/D sky130_fd_sc_hd__clkbuf_1
X_21399_ _21752_/A VGND VGND VPWR VPWR _21399_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23138_ _23138_/A VGND VGND VPWR VPWR _32158_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28995_ _28995_/A VGND VGND VPWR VPWR _34804_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27946_ _34307_/Q _24410_/X _27958_/S VGND VGND VPWR VPWR _27947_/A sky130_fd_sc_hd__mux2_1
XTAP_6155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23069_ _23068_/X _32075_/Q _23075_/S VGND VGND VPWR VPWR _23070_/A sky130_fd_sc_hd__mux2_1
XTAP_5410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27877_ _34274_/Q _24307_/X _27895_/S VGND VGND VPWR VPWR _27878_/A sky130_fd_sc_hd__mux2_1
XTAP_5476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17630_ _32506_/Q _32378_/Q _32058_/Q _36026_/Q _17629_/X _17417_/X VGND VGND VPWR
+ VPWR _17630_/X sky130_fd_sc_hd__mux4_1
X_29616_ _29616_/A VGND VGND VPWR VPWR _35067_/D sky130_fd_sc_hd__clkbuf_1
X_26828_ _26828_/A VGND VGND VPWR VPWR _33807_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17561_ _32760_/Q _32696_/Q _32632_/Q _36088_/Q _17272_/X _17409_/X VGND VGND VPWR
+ VPWR _17561_/X sky130_fd_sc_hd__mux4_1
X_29547_ _29547_/A VGND VGND VPWR VPWR _35034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26759_ _33776_/Q _24351_/X _26769_/S VGND VGND VPWR VPWR _26760_/A sky130_fd_sc_hd__mux2_1
X_19300_ _35560_/Q _35496_/Q _35432_/Q _35368_/Q _19197_/X _19198_/X VGND VGND VPWR
+ VPWR _19300_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_1043 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16512_ _35546_/Q _35482_/Q _35418_/Q _35354_/Q _16191_/X _16192_/X VGND VGND VPWR
+ VPWR _16512_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29478_ _23283_/X _35002_/Q _29488_/S VGND VGND VPWR VPWR _29479_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17492_ _35830_/Q _32208_/Q _35702_/Q _35638_/Q _17313_/X _17314_/X VGND VGND VPWR
+ VPWR _17492_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19231_ _35558_/Q _35494_/Q _35430_/Q _35366_/Q _19197_/X _19198_/X VGND VGND VPWR
+ VPWR _19231_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28429_ _26903_/X _34536_/Q _28435_/S VGND VGND VPWR VPWR _28430_/A sky130_fd_sc_hd__mux2_1
X_16443_ _17149_/A VGND VGND VPWR VPWR _16443_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19162_ _35812_/Q _32188_/Q _35684_/Q _35620_/Q _18907_/X _18908_/X VGND VGND VPWR
+ VPWR _19162_/X sky130_fd_sc_hd__mux4_1
X_31440_ _31440_/A VGND VGND VPWR VPWR _35931_/D sky130_fd_sc_hd__clkbuf_1
X_16374_ _35286_/Q _35222_/Q _35158_/Q _32278_/Q _16300_/X _16301_/X VGND VGND VPWR
+ VPWR _16374_/X sky130_fd_sc_hd__mux4_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18113_ _33224_/Q _32584_/Q _35976_/Q _35912_/Q _16075_/X _16076_/X VGND VGND VPWR
+ VPWR _18113_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31371_ _35899_/Q input40/X _31379_/S VGND VGND VPWR VPWR _31372_/A sky130_fd_sc_hd__mux2_1
X_19093_ _18946_/X _19091_/X _19092_/X _18949_/X VGND VGND VPWR VPWR _19093_/X sky130_fd_sc_hd__a22o_1
XFILLER_12_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33110_ _36117_/CLK _33110_/D VGND VGND VPWR VPWR _33110_/Q sky130_fd_sc_hd__dfxtp_1
X_30322_ _30322_/A VGND VGND VPWR VPWR _35402_/D sky130_fd_sc_hd__clkbuf_1
X_18044_ _17761_/X _18042_/X _18043_/X _17767_/X VGND VGND VPWR VPWR _18044_/X sky130_fd_sc_hd__a22o_1
XFILLER_172_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34090_ _34154_/CLK _34090_/D VGND VGND VPWR VPWR _34090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33041_ _36114_/CLK _33041_/D VGND VGND VPWR VPWR _33041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_153_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _35334_/CLK sky130_fd_sc_hd__clkbuf_16
X_30253_ _30253_/A VGND VGND VPWR VPWR _35369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30184_ _35337_/Q _29234_/X _30184_/S VGND VGND VPWR VPWR _30185_/A sky130_fd_sc_hd__mux2_1
X_19995_ _20129_/A VGND VGND VPWR VPWR _19995_/X sky130_fd_sc_hd__buf_4
XFILLER_99_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18946_ _20160_/A VGND VGND VPWR VPWR _18946_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34992_ _35953_/CLK _34992_/D VGND VGND VPWR VPWR _34992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33943_ _36220_/CLK _33943_/D VGND VGND VPWR VPWR _33943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18877_ _18588_/X _18875_/X _18876_/X _18591_/X VGND VGND VPWR VPWR _18877_/X sky130_fd_sc_hd__a22o_1
XFILLER_227_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17828_ _17548_/X _17826_/X _17827_/X _17553_/X VGND VGND VPWR VPWR _17828_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33874_ _34004_/CLK _33874_/D VGND VGND VPWR VPWR _33874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35613_ _35745_/CLK _35613_/D VGND VGND VPWR VPWR _35613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32825_ _32954_/CLK _32825_/D VGND VGND VPWR VPWR _32825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17759_ _17555_/X _17757_/X _17758_/X _17558_/X VGND VGND VPWR VPWR _17759_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35544_ _36001_/CLK _35544_/D VGND VGND VPWR VPWR _35544_/Q sky130_fd_sc_hd__dfxtp_1
X_20770_ _20687_/X _20768_/X _20769_/X _20697_/X VGND VGND VPWR VPWR _20770_/X sky130_fd_sc_hd__a22o_1
XFILLER_165_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32756_ _36149_/CLK _32756_/D VGND VGND VPWR VPWR _32756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19429_ _19422_/X _19427_/X _19428_/X VGND VGND VPWR VPWR _19463_/A sky130_fd_sc_hd__o21ba_1
X_31707_ _36058_/Q input4/X _31721_/S VGND VGND VPWR VPWR _31708_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35475_ _35922_/CLK _35475_/D VGND VGND VPWR VPWR _35475_/Q sky130_fd_sc_hd__dfxtp_1
X_32687_ _36078_/CLK _32687_/D VGND VGND VPWR VPWR _32687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22440_ _33024_/Q _32960_/Q _32896_/Q _32832_/Q _22295_/X _22296_/X VGND VGND VPWR
+ VPWR _22440_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34426_ _35579_/CLK _34426_/D VGND VGND VPWR VPWR _34426_/Q sky130_fd_sc_hd__dfxtp_1
X_31638_ _31638_/A VGND VGND VPWR VPWR _36025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22371_ _32510_/Q _32382_/Q _32062_/Q _36030_/Q _22229_/X _22370_/X VGND VGND VPWR
+ VPWR _22371_/X sky130_fd_sc_hd__mux4_1
X_34357_ _34805_/CLK _34357_/D VGND VGND VPWR VPWR _34357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31569_ _31569_/A VGND VGND VPWR VPWR _35992_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_392_CLK clkbuf_6_34__f_CLK/X VGND VGND VPWR VPWR _35054_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24110_ _24242_/S VGND VGND VPWR VPWR _24129_/S sky130_fd_sc_hd__clkbuf_4
X_21322_ _22532_/A VGND VGND VPWR VPWR _21322_/X sky130_fd_sc_hd__buf_4
X_33308_ _34074_/CLK _33308_/D VGND VGND VPWR VPWR _33308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25090_ _25090_/A VGND VGND VPWR VPWR _33005_/D sky130_fd_sc_hd__clkbuf_1
X_34288_ _34288_/CLK _34288_/D VGND VGND VPWR VPWR _34288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36027_ _36027_/CLK _36027_/D VGND VGND VPWR VPWR _36027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24041_ _24041_/A VGND VGND VPWR VPWR _32557_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_144_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _35789_/CLK sky130_fd_sc_hd__clkbuf_16
X_33239_ _36118_/CLK _33239_/D VGND VGND VPWR VPWR _33239_/Q sky130_fd_sc_hd__dfxtp_1
X_21253_ _22312_/A VGND VGND VPWR VPWR _21253_/X sky130_fd_sc_hd__buf_6
XFILLER_190_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20204_ _33794_/Q _33730_/Q _33666_/Q _33602_/Q _20202_/X _20203_/X VGND VGND VPWR
+ VPWR _20204_/X sky130_fd_sc_hd__mux4_1
X_21184_ _34780_/Q _34716_/Q _34652_/Q _34588_/Q _21182_/X _21183_/X VGND VGND VPWR
+ VPWR _21184_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27800_ _34238_/Q _24394_/X _27802_/S VGND VGND VPWR VPWR _27801_/A sky130_fd_sc_hd__mux2_1
X_20135_ _20128_/X _20133_/X _20134_/X VGND VGND VPWR VPWR _20169_/A sky130_fd_sc_hd__o21ba_1
X_28780_ _26821_/X _34702_/Q _28798_/S VGND VGND VPWR VPWR _28781_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25992_ _25992_/A VGND VGND VPWR VPWR _33413_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27731_ _34205_/Q _24292_/X _27739_/S VGND VGND VPWR VPWR _27732_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20066_ _33278_/Q _36158_/Q _33150_/Q _33086_/Q _20064_/X _20065_/X VGND VGND VPWR
+ VPWR _20066_/X sky130_fd_sc_hd__mux4_1
XFILLER_161_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24943_ _24943_/A VGND VGND VPWR VPWR _32951_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27662_ _27662_/A VGND VGND VPWR VPWR _34172_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24874_ _22907_/X _32919_/Q _24874_/S VGND VGND VPWR VPWR _24875_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29401_ _29401_/A VGND VGND VPWR VPWR _34965_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26613_ _26613_/A VGND VGND VPWR VPWR _33707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23825_ _23825_/A VGND VGND VPWR VPWR _32456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_304 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27593_ _27593_/A VGND VGND VPWR VPWR _34139_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_315 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_326 _32141_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_337 _32141_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29332_ _23267_/X _34933_/Q _29332_/S VGND VGND VPWR VPWR _29333_/A sky130_fd_sc_hd__mux2_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26544_ _26544_/A VGND VGND VPWR VPWR _33675_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_348 _36205_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23756_ _23756_/A VGND VGND VPWR VPWR _32423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20968_ _22531_/A VGND VGND VPWR VPWR _20968_/X sky130_fd_sc_hd__buf_6
XANTENNA_359 _36207_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22707_ _21754_/A _22705_/X _22706_/X _21759_/A VGND VGND VPWR VPWR _22707_/X sky130_fd_sc_hd__a22o_1
XFILLER_14_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29263_ _23105_/X _34900_/Q _29269_/S VGND VGND VPWR VPWR _29264_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23687_ _23687_/A VGND VGND VPWR VPWR _32392_/D sky130_fd_sc_hd__clkbuf_1
X_26475_ _26475_/A VGND VGND VPWR VPWR _33642_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20899_ _34772_/Q _34708_/Q _34644_/Q _34580_/Q _20829_/X _20830_/X VGND VGND VPWR
+ VPWR _20899_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28214_ _26984_/X _34434_/Q _28228_/S VGND VGND VPWR VPWR _28215_/A sky130_fd_sc_hd__mux2_1
X_22638_ _33542_/Q _33478_/Q _33414_/Q _33350_/Q _22429_/X _22430_/X VGND VGND VPWR
+ VPWR _22638_/X sky130_fd_sc_hd__mux4_1
X_25426_ _25426_/A VGND VGND VPWR VPWR _33149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29194_ input41/X VGND VGND VPWR VPWR _29194_/X sky130_fd_sc_hd__clkbuf_4
X_28145_ _28145_/A VGND VGND VPWR VPWR _34401_/D sky130_fd_sc_hd__clkbuf_1
X_25357_ _25357_/A VGND VGND VPWR VPWR _33116_/D sky130_fd_sc_hd__clkbuf_1
X_22569_ _22569_/A _22569_/B _22569_/C _22569_/D VGND VGND VPWR VPWR _22570_/A sky130_fd_sc_hd__or4_4
Xclkbuf_leaf_383_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _36141_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_167_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16090_ _16873_/A VGND VGND VPWR VPWR _16090_/X sky130_fd_sc_hd__buf_4
X_24308_ _24401_/A VGND VGND VPWR VPWR _24336_/S sky130_fd_sc_hd__clkbuf_4
X_28076_ _28076_/A VGND VGND VPWR VPWR _34368_/D sky130_fd_sc_hd__clkbuf_1
X_25288_ _25288_/A VGND VGND VPWR VPWR _33084_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27027_ _26829_/X _33872_/Q _27041_/S VGND VGND VPWR VPWR _27028_/A sky130_fd_sc_hd__mux2_1
X_24239_ _24239_/A VGND VGND VPWR VPWR _32651_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_135_CLK clkbuf_6_22__f_CLK/X VGND VGND VPWR VPWR _35792_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_177_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18800_ _18796_/X _18797_/X _18798_/X _18799_/X VGND VGND VPWR VPWR _18800_/X sky130_fd_sc_hd__a22o_1
XFILLER_218_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19780_ _19502_/X _19778_/X _19779_/X _19505_/X VGND VGND VPWR VPWR _19780_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28978_ _34796_/Q _24338_/X _28996_/S VGND VGND VPWR VPWR _28979_/A sky130_fd_sc_hd__mux2_1
X_16992_ _16710_/X _16988_/X _16991_/X _16714_/X VGND VGND VPWR VPWR _16992_/X sky130_fd_sc_hd__a22o_1
XFILLER_235_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18731_ _20143_/A VGND VGND VPWR VPWR _18731_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27929_ _34299_/Q _24385_/X _27937_/S VGND VGND VPWR VPWR _27930_/A sky130_fd_sc_hd__mux2_1
XTAP_5251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18662_ _18657_/X _18659_/X _18660_/X _18661_/X VGND VGND VPWR VPWR _18662_/X sky130_fd_sc_hd__a22o_1
X_30940_ _30940_/A VGND VGND VPWR VPWR _35694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17613_ _35065_/Q _35001_/Q _34937_/Q _34873_/Q _17509_/X _17510_/X VGND VGND VPWR
+ VPWR _17613_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18593_ _20160_/A VGND VGND VPWR VPWR _18593_/X sky130_fd_sc_hd__buf_4
X_30871_ _31003_/S VGND VGND VPWR VPWR _30890_/S sky130_fd_sc_hd__buf_4
XFILLER_40_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32610_ _36067_/CLK _32610_/D VGND VGND VPWR VPWR _32610_/Q sky130_fd_sc_hd__dfxtp_1
X_17544_ _17507_/X _17542_/X _17543_/X _17512_/X VGND VGND VPWR VPWR _17544_/X sky130_fd_sc_hd__a22o_1
XTAP_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33590_ _34293_/CLK _33590_/D VGND VGND VPWR VPWR _33590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_860 _24363_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32541_ _35869_/CLK _32541_/D VGND VGND VPWR VPWR _32541_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_871 _24987_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_882 _25084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17475_ _17195_/X _17473_/X _17474_/X _17200_/X VGND VGND VPWR VPWR _17475_/X sky130_fd_sc_hd__a22o_1
XANTENNA_893 _25735_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19214_ _19142_/X _19212_/X _19213_/X _19147_/X VGND VGND VPWR VPWR _19214_/X sky130_fd_sc_hd__a22o_1
XFILLER_242_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35260_ _35326_/CLK _35260_/D VGND VGND VPWR VPWR _35260_/Q sky130_fd_sc_hd__dfxtp_1
X_16426_ _16349_/X _16424_/X _16425_/X _16355_/X VGND VGND VPWR VPWR _16426_/X sky130_fd_sc_hd__a22o_1
X_32472_ _35994_/CLK _32472_/D VGND VGND VPWR VPWR _32472_/Q sky130_fd_sc_hd__dfxtp_1
X_34211_ _34276_/CLK _34211_/D VGND VGND VPWR VPWR _34211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31423_ _31423_/A VGND VGND VPWR VPWR _35923_/D sky130_fd_sc_hd__clkbuf_1
X_19145_ _33764_/Q _33700_/Q _33636_/Q _33572_/Q _19143_/X _19144_/X VGND VGND VPWR
+ VPWR _19145_/X sky130_fd_sc_hd__mux4_1
X_16357_ _17908_/A VGND VGND VPWR VPWR _16357_/X sky130_fd_sc_hd__buf_4
X_35191_ _35320_/CLK _35191_/D VGND VGND VPWR VPWR _35191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_374_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _36078_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34142_ _34142_/CLK _34142_/D VGND VGND VPWR VPWR _34142_/Q sky130_fd_sc_hd__dfxtp_1
X_31354_ _35891_/Q input31/X _31358_/S VGND VGND VPWR VPWR _31355_/A sky130_fd_sc_hd__mux2_1
X_19076_ _19069_/X _19074_/X _19075_/X VGND VGND VPWR VPWR _19110_/A sky130_fd_sc_hd__o21ba_1
XFILLER_121_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16288_ _17855_/A VGND VGND VPWR VPWR _16288_/X sky130_fd_sc_hd__buf_4
Xclkbuf_5_31_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_31_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_117_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18027_ _35333_/Q _35269_/Q _35205_/Q _32325_/Q _17712_/X _17713_/X VGND VGND VPWR
+ VPWR _18027_/X sky130_fd_sc_hd__mux4_1
X_30305_ _35394_/Q _29213_/X _30319_/S VGND VGND VPWR VPWR _30306_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_126_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _34197_/CLK sky130_fd_sc_hd__clkbuf_16
X_34073_ _34265_/CLK _34073_/D VGND VGND VPWR VPWR _34073_/Q sky130_fd_sc_hd__dfxtp_1
X_31285_ _35858_/Q input45/X _31295_/S VGND VGND VPWR VPWR _31286_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33024_ _36159_/CLK _33024_/D VGND VGND VPWR VPWR _33024_/Q sky130_fd_sc_hd__dfxtp_1
X_30236_ _30236_/A VGND VGND VPWR VPWR _35361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30167_ _30167_/A VGND VGND VPWR VPWR _35328_/D sky130_fd_sc_hd__clkbuf_1
X_19978_ _34555_/Q _32443_/Q _34427_/Q _34363_/Q _19878_/X _19879_/X VGND VGND VPWR
+ VPWR _19978_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18929_ _34014_/Q _33950_/Q _33886_/Q _32158_/Q _18614_/X _18615_/X VGND VGND VPWR
+ VPWR _18929_/X sky130_fd_sc_hd__mux4_1
X_30098_ _35296_/Q _29107_/X _30100_/S VGND VGND VPWR VPWR _30099_/A sky130_fd_sc_hd__mux2_1
XANTENNA_1270 _31003_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_34975_ _35040_/CLK _34975_/D VGND VGND VPWR VPWR _34975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1281 _17834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1292 _17932_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21940_ _21655_/X _21938_/X _21939_/X _21661_/X VGND VGND VPWR VPWR _21940_/X sky130_fd_sc_hd__a22o_1
X_33926_ _34243_/CLK _33926_/D VGND VGND VPWR VPWR _33926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33857_ _35777_/CLK _33857_/D VGND VGND VPWR VPWR _33857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21871_ _21867_/X _21870_/X _21728_/X VGND VGND VPWR VPWR _21897_/A sky130_fd_sc_hd__o21ba_1
XFILLER_131_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23610_ _23610_/A VGND VGND VPWR VPWR _32355_/D sky130_fd_sc_hd__clkbuf_1
X_20822_ _35794_/Q _32168_/Q _35666_/Q _35602_/Q _20645_/X _20646_/X VGND VGND VPWR
+ VPWR _20822_/X sky130_fd_sc_hd__mux4_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32808_ _36009_/CLK _32808_/D VGND VGND VPWR VPWR _32808_/Q sky130_fd_sc_hd__dfxtp_1
X_24590_ _22889_/X _32785_/Q _24602_/S VGND VGND VPWR VPWR _24591_/A sky130_fd_sc_hd__mux2_1
X_33788_ _34044_/CLK _33788_/D VGND VGND VPWR VPWR _33788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23541_ _23047_/X _32324_/Q _23551_/S VGND VGND VPWR VPWR _23542_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35527_ _35590_/CLK _35527_/D VGND VGND VPWR VPWR _35527_/Q sky130_fd_sc_hd__dfxtp_1
X_20753_ _32976_/Q _32912_/Q _32848_/Q _32784_/Q _20633_/X _20635_/X VGND VGND VPWR
+ VPWR _20753_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32739_ _36067_/CLK _32739_/D VGND VGND VPWR VPWR _32739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26260_ _26260_/A VGND VGND VPWR VPWR _33540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1099 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35458_ _35970_/CLK _35458_/D VGND VGND VPWR VPWR _35458_/Q sky130_fd_sc_hd__dfxtp_1
X_23472_ _22945_/X _32291_/Q _23488_/S VGND VGND VPWR VPWR _23473_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20684_ _21752_/A VGND VGND VPWR VPWR _20684_/X sky130_fd_sc_hd__buf_4
XFILLER_51_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25211_ _25322_/S VGND VGND VPWR VPWR _25230_/S sky130_fd_sc_hd__buf_4
X_22423_ _22419_/X _22422_/X _22114_/X VGND VGND VPWR VPWR _22424_/D sky130_fd_sc_hd__o21ba_1
XFILLER_137_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34409_ _34987_/CLK _34409_/D VGND VGND VPWR VPWR _34409_/Q sky130_fd_sc_hd__dfxtp_1
X_26191_ _26191_/A VGND VGND VPWR VPWR _33507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35389_ _35517_/CLK _35389_/D VGND VGND VPWR VPWR _35389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_365_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _33520_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25142_ _25142_/A VGND VGND VPWR VPWR _33022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22354_ _33790_/Q _33726_/Q _33662_/Q _33598_/Q _22149_/X _22150_/X VGND VGND VPWR
+ VPWR _22354_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21305_ _22502_/A VGND VGND VPWR VPWR _21305_/X sky130_fd_sc_hd__buf_4
XFILLER_237_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_117_CLK clkbuf_6_20__f_CLK/X VGND VGND VPWR VPWR _35280_/CLK sky130_fd_sc_hd__clkbuf_16
X_29950_ _29950_/A VGND VGND VPWR VPWR _35225_/D sky130_fd_sc_hd__clkbuf_1
X_25073_ _25072_/X _33000_/Q _25082_/S VGND VGND VPWR VPWR _25074_/A sky130_fd_sc_hd__mux2_1
X_22285_ _34300_/Q _34236_/Q _34172_/Q _34108_/Q _22042_/X _22043_/X VGND VGND VPWR
+ VPWR _22285_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28901_ _27002_/X _34760_/Q _28903_/S VGND VGND VPWR VPWR _28902_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24024_ _24024_/A VGND VGND VPWR VPWR _32549_/D sky130_fd_sc_hd__clkbuf_1
X_21236_ _22429_/A VGND VGND VPWR VPWR _21236_/X sky130_fd_sc_hd__buf_4
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29881_ _35193_/Q _29185_/X _29893_/S VGND VGND VPWR VPWR _29882_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28832_ _26900_/X _34727_/Q _28840_/S VGND VGND VPWR VPWR _28833_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21167_ _32732_/Q _32668_/Q _32604_/Q _36060_/Q _21166_/X _20950_/X VGND VGND VPWR
+ VPWR _21167_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_1471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20118_ _35327_/Q _35263_/Q _35199_/Q _32319_/Q _20012_/X _20013_/X VGND VGND VPWR
+ VPWR _20118_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28763_ _28763_/A VGND VGND VPWR VPWR _34694_/D sky130_fd_sc_hd__clkbuf_1
X_25975_ _25975_/A VGND VGND VPWR VPWR _33405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21098_ _34010_/Q _33946_/Q _33882_/Q _32154_/Q _20914_/X _20915_/X VGND VGND VPWR
+ VPWR _21098_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27714_ _34197_/Q _24267_/X _27718_/S VGND VGND VPWR VPWR _27715_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20049_ _35069_/Q _35005_/Q _34941_/Q _34877_/Q _19809_/X _19810_/X VGND VGND VPWR
+ VPWR _20049_/X sky130_fd_sc_hd__mux4_1
X_24926_ _24926_/A VGND VGND VPWR VPWR _32943_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28694_ _28694_/A VGND VGND VPWR VPWR _34661_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27645_ _27645_/A VGND VGND VPWR VPWR _34164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24857_ _24857_/A VGND VGND VPWR VPWR _32910_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_101 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_112 _32129_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23808_ _23034_/X _32448_/Q _23826_/S VGND VGND VPWR VPWR _23809_/A sky130_fd_sc_hd__mux2_1
XANTENNA_134 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27576_ _27576_/A VGND VGND VPWR VPWR _34131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_226_1403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24788_ _22979_/X _32878_/Q _24802_/S VGND VGND VPWR VPWR _24789_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_156 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29315_ _29315_/A VGND VGND VPWR VPWR _34924_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26527_ _25156_/X _33667_/Q _26539_/S VGND VGND VPWR VPWR _26528_/A sky130_fd_sc_hd__mux2_1
XANTENNA_178 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23739_ _23739_/A VGND VGND VPWR VPWR _32415_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_189 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29246_ input60/X VGND VGND VPWR VPWR _29246_/X sky130_fd_sc_hd__buf_2
X_17260_ _35055_/Q _34991_/Q _34927_/Q _34863_/Q _17156_/X _17157_/X VGND VGND VPWR
+ VPWR _17260_/X sky130_fd_sc_hd__mux4_1
XFILLER_187_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26458_ _25053_/X _33634_/Q _26476_/S VGND VGND VPWR VPWR _26459_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16211_ _16143_/X _16209_/X _16210_/X _16146_/X VGND VGND VPWR VPWR _16211_/X sky130_fd_sc_hd__a22o_1
XFILLER_220_1002 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25409_ _25409_/A VGND VGND VPWR VPWR _33141_/D sky130_fd_sc_hd__clkbuf_1
X_29177_ _34870_/Q _29175_/X _29204_/S VGND VGND VPWR VPWR _29178_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17191_ _17154_/X _17189_/X _17190_/X _17159_/X VGND VGND VPWR VPWR _17191_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_356_CLK clkbuf_6_41__f_CLK/X VGND VGND VPWR VPWR _35827_/CLK sky130_fd_sc_hd__clkbuf_16
X_26389_ _26389_/A VGND VGND VPWR VPWR _33601_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16142_ _16136_/X _16139_/X _16140_/X _16141_/X VGND VGND VPWR VPWR _16142_/X sky130_fd_sc_hd__a22o_1
X_28128_ _26857_/X _34393_/Q _28144_/S VGND VGND VPWR VPWR _28129_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_108_CLK clkbuf_6_22__f_CLK/X VGND VGND VPWR VPWR _35728_/CLK sky130_fd_sc_hd__clkbuf_16
X_16073_ _17761_/A VGND VGND VPWR VPWR _17149_/A sky130_fd_sc_hd__buf_12
XFILLER_142_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28059_ _28059_/A VGND VGND VPWR VPWR _34360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19901_ _35769_/Q _35129_/Q _34489_/Q _33849_/Q _19793_/X _19794_/X VGND VGND VPWR
+ VPWR _19901_/X sky130_fd_sc_hd__mux4_1
X_31070_ _35756_/Q _29144_/X _31088_/S VGND VGND VPWR VPWR _31071_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30021_ _30021_/A VGND VGND VPWR VPWR _35259_/D sky130_fd_sc_hd__clkbuf_1
X_19832_ _35831_/Q _32209_/Q _35703_/Q _35639_/Q _19613_/X _19614_/X VGND VGND VPWR
+ VPWR _19832_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19763_ _19759_/X _19762_/X _19447_/X VGND VGND VPWR VPWR _19771_/C sky130_fd_sc_hd__o21ba_1
XFILLER_111_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16975_ _16971_/X _16974_/X _16808_/X VGND VGND VPWR VPWR _16976_/D sky130_fd_sc_hd__o21ba_1
XFILLER_7_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18714_ _33752_/Q _33688_/Q _33624_/Q _33560_/Q _18437_/X _18438_/X VGND VGND VPWR
+ VPWR _18714_/X sky130_fd_sc_hd__mux4_1
X_34760_ _35337_/CLK _34760_/D VGND VGND VPWR VPWR _34760_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31972_ _34970_/CLK _31972_/D VGND VGND VPWR VPWR _31972_/Q sky130_fd_sc_hd__dfxtp_1
X_19694_ _19449_/X _19692_/X _19693_/X _19452_/X VGND VGND VPWR VPWR _19694_/X sky130_fd_sc_hd__a22o_1
XTAP_5081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 DW[15] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__buf_8
XFILLER_77_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33711_ _33775_/CLK _33711_/D VGND VGND VPWR VPWR _33711_/Q sky130_fd_sc_hd__dfxtp_1
X_18645_ _33494_/Q _33430_/Q _33366_/Q _33302_/Q _18298_/X _18299_/X VGND VGND VPWR
+ VPWR _18645_/X sky130_fd_sc_hd__mux4_1
XFILLER_209_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30923_ _30923_/A VGND VGND VPWR VPWR _35686_/D sky130_fd_sc_hd__clkbuf_1
X_34691_ _35331_/CLK _34691_/D VGND VGND VPWR VPWR _34691_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33642_ _34281_/CLK _33642_/D VGND VGND VPWR VPWR _33642_/Q sky130_fd_sc_hd__dfxtp_1
X_18576_ _34004_/Q _33940_/Q _33876_/Q _32148_/Q _18408_/X _18409_/X VGND VGND VPWR
+ VPWR _18576_/X sky130_fd_sc_hd__mux4_1
X_30854_ _23322_/X _35654_/Q _30860_/S VGND VGND VPWR VPWR _30855_/A sky130_fd_sc_hd__mux2_1
XTAP_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17527_ _17408_/X _17525_/X _17526_/X _17414_/X VGND VGND VPWR VPWR _17527_/X sky130_fd_sc_hd__a22o_1
XFILLER_205_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33573_ _33702_/CLK _33573_/D VGND VGND VPWR VPWR _33573_/Q sky130_fd_sc_hd__dfxtp_1
X_30785_ _23199_/X _35621_/Q _30797_/S VGND VGND VPWR VPWR _30786_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_1394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35312_ _35757_/CLK _35312_/D VGND VGND VPWR VPWR _35312_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_690 _22443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32524_ _36109_/CLK _32524_/D VGND VGND VPWR VPWR _32524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17458_ _35765_/Q _35125_/Q _34485_/Q _33845_/Q _17140_/X _17141_/X VGND VGND VPWR
+ VPWR _17458_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_1378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16409_ _35031_/Q _34967_/Q _34903_/Q _34839_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _16409_/X sky130_fd_sc_hd__mux4_1
X_35243_ _35307_/CLK _35243_/D VGND VGND VPWR VPWR _35243_/Q sky130_fd_sc_hd__dfxtp_1
X_32455_ _35078_/CLK _32455_/D VGND VGND VPWR VPWR _32455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_347_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _33779_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17389_ _33203_/Q _32563_/Q _35955_/Q _35891_/Q _17074_/X _17075_/X VGND VGND VPWR
+ VPWR _17389_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31406_ _35916_/Q input59/X _31408_/S VGND VGND VPWR VPWR _31407_/A sky130_fd_sc_hd__mux2_1
X_19128_ _18941_/X _19126_/X _19127_/X _18944_/X VGND VGND VPWR VPWR _19128_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35174_ _35239_/CLK _35174_/D VGND VGND VPWR VPWR _35174_/Q sky130_fd_sc_hd__dfxtp_1
X_32386_ _32962_/CLK _32386_/D VGND VGND VPWR VPWR _32386_/Q sky130_fd_sc_hd__dfxtp_1
X_34125_ _34317_/CLK _34125_/D VGND VGND VPWR VPWR _34125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31337_ _35883_/Q input22/X _31337_/S VGND VGND VPWR VPWR _31338_/A sky130_fd_sc_hd__mux2_1
X_19059_ _35297_/Q _35233_/Q _35169_/Q _32289_/Q _18953_/X _18954_/X VGND VGND VPWR
+ VPWR _19059_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34056_ _34243_/CLK _34056_/D VGND VGND VPWR VPWR _34056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22070_ _22066_/X _22069_/X _21761_/X VGND VGND VPWR VPWR _22071_/D sky130_fd_sc_hd__o21ba_1
X_31268_ _31268_/A VGND VGND VPWR VPWR _35850_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21021_ _20743_/X _21019_/X _21020_/X _20746_/X VGND VGND VPWR VPWR _21021_/X sky130_fd_sc_hd__a22o_1
X_33007_ _33007_/CLK _33007_/D VGND VGND VPWR VPWR _33007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30219_ _35353_/Q _29086_/X _30235_/S VGND VGND VPWR VPWR _30220_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31199_ _31199_/A VGND VGND VPWR VPWR _35817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25760_ _25760_/A VGND VGND VPWR VPWR _33303_/D sky130_fd_sc_hd__clkbuf_1
X_22972_ input24/X VGND VGND VPWR VPWR _22972_/X sky130_fd_sc_hd__buf_4
XFILLER_101_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34958_ _35026_/CLK _34958_/D VGND VGND VPWR VPWR _34958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24711_ _23068_/X _32843_/Q _24715_/S VGND VGND VPWR VPWR _24712_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21923_ _35313_/Q _35249_/Q _35185_/Q _32305_/Q _21606_/X _21607_/X VGND VGND VPWR
+ VPWR _21923_/X sky130_fd_sc_hd__mux4_1
X_33909_ _36149_/CLK _33909_/D VGND VGND VPWR VPWR _33909_/Q sky130_fd_sc_hd__dfxtp_1
X_25691_ _25691_/A VGND VGND VPWR VPWR _33271_/D sky130_fd_sc_hd__clkbuf_1
X_34889_ _35781_/CLK _34889_/D VGND VGND VPWR VPWR _34889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27430_ _26826_/X _34063_/Q _27446_/S VGND VGND VPWR VPWR _27431_/A sky130_fd_sc_hd__mux2_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21854_ _21599_/X _21852_/X _21853_/X _21602_/X VGND VGND VPWR VPWR _21854_/X sky130_fd_sc_hd__a22o_1
X_24642_ _22966_/X _32810_/Q _24644_/S VGND VGND VPWR VPWR _24643_/A sky130_fd_sc_hd__mux2_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20805_ _20805_/A VGND VGND VPWR VPWR _36177_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27361_ _27361_/A VGND VGND VPWR VPWR _34030_/D sky130_fd_sc_hd__clkbuf_1
X_24573_ _23068_/X _32779_/Q _24577_/S VGND VGND VPWR VPWR _24574_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21785_ _21781_/X _21784_/X _21747_/X VGND VGND VPWR VPWR _21793_/C sky130_fd_sc_hd__o21ba_1
X_29100_ _29100_/A VGND VGND VPWR VPWR _34845_/D sky130_fd_sc_hd__clkbuf_1
X_26312_ _25038_/X _33565_/Q _26320_/S VGND VGND VPWR VPWR _26313_/A sky130_fd_sc_hd__mux2_1
X_20736_ _22455_/A VGND VGND VPWR VPWR _20736_/X sky130_fd_sc_hd__buf_4
XFILLER_211_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23524_ _23022_/X _32316_/Q _23530_/S VGND VGND VPWR VPWR _23525_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27292_ _27424_/S VGND VGND VPWR VPWR _27311_/S sky130_fd_sc_hd__buf_4
XFILLER_180_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29031_ _29031_/A VGND VGND VPWR VPWR _34821_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26243_ _26243_/A VGND VGND VPWR VPWR _33532_/D sky130_fd_sc_hd__clkbuf_1
X_23455_ _22920_/X _32283_/Q _23467_/S VGND VGND VPWR VPWR _23456_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20667_ _22373_/A VGND VGND VPWR VPWR _22465_/A sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_338_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _36152_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_196_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22406_ _32511_/Q _32383_/Q _32063_/Q _36031_/Q _22229_/X _22370_/X VGND VGND VPWR
+ VPWR _22406_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23386_ _32252_/Q _23289_/X _23392_/S VGND VGND VPWR VPWR _23387_/A sky130_fd_sc_hd__mux2_1
X_26174_ _26174_/A VGND VGND VPWR VPWR _33499_/D sky130_fd_sc_hd__clkbuf_1
X_20598_ _22395_/A VGND VGND VPWR VPWR _20598_/X sky130_fd_sc_hd__buf_4
X_22337_ _22333_/X _22336_/X _22089_/X _22090_/X VGND VGND VPWR VPWR _22352_/B sky130_fd_sc_hd__o211a_1
X_25125_ input38/X VGND VGND VPWR VPWR _25125_/X sky130_fd_sc_hd__buf_2
XFILLER_139_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29933_ _29933_/A VGND VGND VPWR VPWR _35217_/D sky130_fd_sc_hd__clkbuf_1
X_25056_ _25056_/A VGND VGND VPWR VPWR _32994_/D sky130_fd_sc_hd__clkbuf_1
X_22268_ _35835_/Q _32213_/Q _35707_/Q _35643_/Q _22266_/X _22267_/X VGND VGND VPWR
+ VPWR _22268_/X sky130_fd_sc_hd__mux4_1
X_24007_ _24007_/A VGND VGND VPWR VPWR _32541_/D sky130_fd_sc_hd__clkbuf_1
X_21219_ _34525_/Q _32413_/Q _34397_/Q _34333_/Q _21119_/X _21120_/X VGND VGND VPWR
+ VPWR _21219_/X sky130_fd_sc_hd__mux4_1
X_29864_ _35185_/Q _29160_/X _29872_/S VGND VGND VPWR VPWR _29865_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22199_ _22195_/X _22198_/X _22089_/X _22090_/X VGND VGND VPWR VPWR _22216_/B sky130_fd_sc_hd__o211a_1
XFILLER_116_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28815_ _26875_/X _34719_/Q _28819_/S VGND VGND VPWR VPWR _28816_/A sky130_fd_sc_hd__mux2_1
X_29795_ _35152_/Q _29058_/X _29809_/S VGND VGND VPWR VPWR _29796_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28746_ _28746_/A VGND VGND VPWR VPWR _34686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16760_ _16443_/X _16758_/X _16759_/X _16446_/X VGND VGND VPWR VPWR _16760_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25958_ _25958_/A VGND VGND VPWR VPWR _33397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24909_ _24909_/A VGND VGND VPWR VPWR _32935_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16691_ _16448_/X _16689_/X _16690_/X _16453_/X VGND VGND VPWR VPWR _16691_/X sky130_fd_sc_hd__a22o_1
X_28677_ _28677_/A VGND VGND VPWR VPWR _34653_/D sky130_fd_sc_hd__clkbuf_1
X_25889_ _25889_/A VGND VGND VPWR VPWR _33364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18430_ _34511_/Q _32399_/Q _34383_/Q _34319_/Q _18388_/X _18390_/X VGND VGND VPWR
+ VPWR _18430_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27628_ _34156_/Q _24338_/X _27646_/S VGND VGND VPWR VPWR _27629_/A sky130_fd_sc_hd__mux2_1
XFILLER_234_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _35534_/Q _35470_/Q _35406_/Q _35342_/Q _18358_/X _18360_/X VGND VGND VPWR
+ VPWR _18361_/X sky130_fd_sc_hd__mux4_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27559_ _27017_/X _34125_/Q _27559_/S VGND VGND VPWR VPWR _27560_/A sky130_fd_sc_hd__mux2_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17312_ _17308_/X _17311_/X _17136_/X _17137_/X VGND VGND VPWR VPWR _17329_/B sky130_fd_sc_hd__o211a_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18292_ _34254_/Q _34190_/Q _34126_/Q _34062_/Q _18289_/X _18291_/X VGND VGND VPWR
+ VPWR _18292_/X sky130_fd_sc_hd__mux4_1
X_30570_ _30570_/A VGND VGND VPWR VPWR _35519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29229_ _34887_/Q _29228_/X _29235_/S VGND VGND VPWR VPWR _29230_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17243_ _32495_/Q _32367_/Q _32047_/Q _36015_/Q _16923_/X _17064_/X VGND VGND VPWR
+ VPWR _17243_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_329_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _36086_/CLK sky130_fd_sc_hd__clkbuf_16
X_32240_ _36146_/CLK _32240_/D VGND VGND VPWR VPWR _32240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17174_ _17055_/X _17172_/X _17173_/X _17061_/X VGND VGND VPWR VPWR _17174_/X sky130_fd_sc_hd__a22o_1
X_16125_ _16056_/X _16123_/X _16124_/X _16068_/X VGND VGND VPWR VPWR _16125_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32171_ _34149_/CLK _32171_/D VGND VGND VPWR VPWR _32171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31122_ _35781_/Q _29222_/X _31130_/S VGND VGND VPWR VPWR _31123_/A sky130_fd_sc_hd__mux2_1
X_16056_ _17860_/A VGND VGND VPWR VPWR _16056_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_115_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31053_ _35748_/Q _29120_/X _31067_/S VGND VGND VPWR VPWR _31054_/A sky130_fd_sc_hd__mux2_1
X_35930_ _35931_/CLK _35930_/D VGND VGND VPWR VPWR _35930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30004_ _30004_/A VGND VGND VPWR VPWR _35251_/D sky130_fd_sc_hd__clkbuf_1
X_19815_ _19806_/X _19813_/X _19814_/X VGND VGND VPWR VPWR _19816_/D sky130_fd_sc_hd__o21ba_1
XFILLER_150_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35861_ _35927_/CLK _35861_/D VGND VGND VPWR VPWR _35861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34812_ _35772_/CLK _34812_/D VGND VGND VPWR VPWR _34812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16958_ _16710_/X _16956_/X _16957_/X _16714_/X VGND VGND VPWR VPWR _16958_/X sky130_fd_sc_hd__a22o_1
X_19746_ _33525_/Q _33461_/Q _33397_/Q _33333_/Q _19423_/X _19424_/X VGND VGND VPWR
+ VPWR _19746_/X sky130_fd_sc_hd__mux4_1
XFILLER_244_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35792_ _35792_/CLK _35792_/D VGND VGND VPWR VPWR _35792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31955_ _35036_/CLK _31955_/D VGND VGND VPWR VPWR _31955_/Q sky130_fd_sc_hd__dfxtp_1
X_19677_ _19671_/X _19676_/X _19428_/X VGND VGND VPWR VPWR _19699_/A sky130_fd_sc_hd__o21ba_1
X_34743_ _35575_/CLK _34743_/D VGND VGND VPWR VPWR _34743_/Q sky130_fd_sc_hd__dfxtp_1
X_16889_ _16702_/X _16887_/X _16888_/X _16708_/X VGND VGND VPWR VPWR _16889_/X sky130_fd_sc_hd__a22o_1
XFILLER_168_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18628_ _18588_/X _18626_/X _18627_/X _18591_/X VGND VGND VPWR VPWR _18628_/X sky130_fd_sc_hd__a22o_1
XFILLER_25_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30906_ _30906_/A VGND VGND VPWR VPWR _35678_/D sky130_fd_sc_hd__clkbuf_1
X_34674_ _34932_/CLK _34674_/D VGND VGND VPWR VPWR _34674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31886_ _23247_/X _36143_/Q _31898_/S VGND VGND VPWR VPWR _31887_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33625_ _35671_/CLK _33625_/D VGND VGND VPWR VPWR _33625_/Q sky130_fd_sc_hd__dfxtp_1
X_30837_ _23297_/X _35646_/Q _30839_/S VGND VGND VPWR VPWR _30838_/A sky130_fd_sc_hd__mux2_1
X_18559_ _35539_/Q _35475_/Q _35411_/Q _35347_/Q _18491_/X _18492_/X VGND VGND VPWR
+ VPWR _18559_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33556_ _33685_/CLK _33556_/D VGND VGND VPWR VPWR _33556_/Q sky130_fd_sc_hd__dfxtp_1
X_21570_ _35303_/Q _35239_/Q _35175_/Q _32295_/Q _21253_/X _21254_/X VGND VGND VPWR
+ VPWR _21570_/X sky130_fd_sc_hd__mux4_1
X_30768_ _23133_/X _35613_/Q _30776_/S VGND VGND VPWR VPWR _30769_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_1096 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_12 _32115_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20521_ _20517_/X _20520_/X _20134_/A VGND VGND VPWR VPWR _20543_/A sky130_fd_sc_hd__o21ba_1
X_32507_ _36092_/CLK _32507_/D VGND VGND VPWR VPWR _32507_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_23 _32115_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 _32117_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33487_ _33490_/CLK _33487_/D VGND VGND VPWR VPWR _33487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30699_ _30699_/A VGND VGND VPWR VPWR _35580_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_45 _32118_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_56 _32126_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_67 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23240_ _23240_/A VGND VGND VPWR VPWR _32197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20452_ _20448_/X _20451_/X _20167_/X VGND VGND VPWR VPWR _20453_/D sky130_fd_sc_hd__o21ba_1
X_32438_ _35768_/CLK _32438_/D VGND VGND VPWR VPWR _32438_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_78 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35226_ _35226_/CLK _35226_/D VGND VGND VPWR VPWR _35226_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_89 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23171_ _32169_/Q _23102_/X _23182_/S VGND VGND VPWR VPWR _23172_/A sky130_fd_sc_hd__mux2_1
X_35157_ _36202_/CLK _35157_/D VGND VGND VPWR VPWR _35157_/Q sky130_fd_sc_hd__dfxtp_1
X_20383_ _33223_/Q _32583_/Q _35975_/Q _35911_/Q _20080_/X _20081_/X VGND VGND VPWR
+ VPWR _20383_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32369_ _36078_/CLK _32369_/D VGND VGND VPWR VPWR _32369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34108_ _36157_/CLK _34108_/D VGND VGND VPWR VPWR _34108_/Q sky130_fd_sc_hd__dfxtp_1
X_22122_ _34039_/Q _33975_/Q _33911_/Q _32247_/Q _21973_/X _21974_/X VGND VGND VPWR
+ VPWR _22122_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35088_ _35279_/CLK _35088_/D VGND VGND VPWR VPWR _35088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput130 _31996_/Q VGND VGND VPWR VPWR D1[46] sky130_fd_sc_hd__buf_2
Xoutput141 _32006_/Q VGND VGND VPWR VPWR D1[56] sky130_fd_sc_hd__buf_2
XTAP_6507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput152 _31958_/Q VGND VGND VPWR VPWR D1[8] sky130_fd_sc_hd__buf_2
XFILLER_88_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput163 _36192_/Q VGND VGND VPWR VPWR D2[18] sky130_fd_sc_hd__buf_2
X_34039_ _34039_/CLK _34039_/D VGND VGND VPWR VPWR _34039_/Q sky130_fd_sc_hd__dfxtp_1
X_26930_ _26930_/A VGND VGND VPWR VPWR _33840_/D sky130_fd_sc_hd__clkbuf_1
X_22053_ _32501_/Q _32373_/Q _32053_/Q _36021_/Q _21876_/X _22017_/X VGND VGND VPWR
+ VPWR _22053_/X sky130_fd_sc_hd__mux4_1
XTAP_6529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput174 _36202_/Q VGND VGND VPWR VPWR D2[28] sky130_fd_sc_hd__buf_2
XFILLER_86_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput185 _36212_/Q VGND VGND VPWR VPWR D2[38] sky130_fd_sc_hd__buf_2
XTAP_5806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput196 _36222_/Q VGND VGND VPWR VPWR D2[48] sky130_fd_sc_hd__buf_2
X_21004_ _21000_/X _21003_/X _20671_/X VGND VGND VPWR VPWR _21012_/C sky130_fd_sc_hd__o21ba_1
XTAP_5817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26861_ _26860_/X _33818_/Q _26882_/S VGND VGND VPWR VPWR _26862_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28600_ _26956_/X _34617_/Q _28612_/S VGND VGND VPWR VPWR _28601_/A sky130_fd_sc_hd__mux2_1
X_25812_ _25097_/X _33328_/Q _25822_/S VGND VGND VPWR VPWR _25813_/A sky130_fd_sc_hd__mux2_1
X_29580_ _29580_/A VGND VGND VPWR VPWR _35050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26792_ _26819_/S VGND VGND VPWR VPWR _26811_/S sky130_fd_sc_hd__buf_6
XFILLER_247_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28531_ _26853_/X _34584_/Q _28549_/S VGND VGND VPWR VPWR _28532_/A sky130_fd_sc_hd__mux2_1
X_25743_ _24995_/X _33295_/Q _25759_/S VGND VGND VPWR VPWR _25744_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22955_ _22954_/X _32038_/Q _22970_/S VGND VGND VPWR VPWR _22956_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28462_ _28462_/A VGND VGND VPWR VPWR _34551_/D sky130_fd_sc_hd__clkbuf_1
X_21906_ _32753_/Q _32689_/Q _32625_/Q _36081_/Q _21872_/X _21656_/X VGND VGND VPWR
+ VPWR _21906_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25674_ _25674_/A VGND VGND VPWR VPWR _33263_/D sky130_fd_sc_hd__clkbuf_1
X_22886_ input23/X VGND VGND VPWR VPWR _22886_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_216_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27413_ _27413_/A VGND VGND VPWR VPWR _34055_/D sky130_fd_sc_hd__clkbuf_1
X_24625_ _24715_/S VGND VGND VPWR VPWR _24644_/S sky130_fd_sc_hd__buf_4
X_28393_ _26850_/X _34519_/Q _28393_/S VGND VGND VPWR VPWR _28394_/A sky130_fd_sc_hd__mux2_1
X_21837_ _34031_/Q _33967_/Q _33903_/Q _32239_/Q _21620_/X _21621_/X VGND VGND VPWR
+ VPWR _21837_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27344_ _27344_/A VGND VGND VPWR VPWR _34022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24556_ _24556_/A VGND VGND VPWR VPWR _32770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21768_ _33517_/Q _33453_/Q _33389_/Q _33325_/Q _21723_/X _21724_/X VGND VGND VPWR
+ VPWR _21768_/X sky130_fd_sc_hd__mux4_2
XFILLER_178_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20719_ _20715_/X _20718_/X _20640_/X _20642_/X VGND VGND VPWR VPWR _20734_/B sky130_fd_sc_hd__o211a_1
X_23507_ _22997_/X _32308_/Q _23509_/S VGND VGND VPWR VPWR _23508_/A sky130_fd_sc_hd__mux2_1
X_27275_ _26996_/X _33990_/Q _27281_/S VGND VGND VPWR VPWR _27276_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21699_ _21655_/X _21697_/X _21698_/X _21661_/X VGND VGND VPWR VPWR _21699_/X sky130_fd_sc_hd__a22o_1
X_24487_ _24577_/S VGND VGND VPWR VPWR _24506_/S sky130_fd_sc_hd__buf_4
XFILLER_106_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29014_ _29014_/A VGND VGND VPWR VPWR _34813_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26226_ _26226_/A VGND VGND VPWR VPWR _33524_/D sky130_fd_sc_hd__clkbuf_1
X_23438_ _22895_/X _32275_/Q _23446_/S VGND VGND VPWR VPWR _23439_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26157_ _26157_/A VGND VGND VPWR VPWR _33491_/D sky130_fd_sc_hd__clkbuf_1
X_23369_ _32244_/Q _23264_/X _23371_/S VGND VGND VPWR VPWR _23370_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25108_ _25108_/A VGND VGND VPWR VPWR _33011_/D sky130_fd_sc_hd__clkbuf_1
X_26088_ _25106_/X _33459_/Q _26092_/S VGND VGND VPWR VPWR _26089_/A sky130_fd_sc_hd__mux2_1
X_17930_ _17855_/X _17928_/X _17929_/X _17858_/X VGND VGND VPWR VPWR _17930_/X sky130_fd_sc_hd__a22o_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29916_ _35210_/Q _29237_/X _29922_/S VGND VGND VPWR VPWR _29917_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25039_ _25038_/X _32989_/Q _25051_/S VGND VGND VPWR VPWR _25040_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17861_ _34560_/Q _32448_/Q _34432_/Q _34368_/Q _17578_/X _17579_/X VGND VGND VPWR
+ VPWR _17861_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29847_ _35177_/Q _29135_/X _29851_/S VGND VGND VPWR VPWR _29848_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_975 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16812_ _33763_/Q _33699_/Q _33635_/Q _33571_/Q _16490_/X _16491_/X VGND VGND VPWR
+ VPWR _16812_/X sky130_fd_sc_hd__mux4_1
X_19600_ _34289_/Q _34225_/Q _34161_/Q _34097_/Q _19389_/X _19390_/X VGND VGND VPWR
+ VPWR _19600_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29778_ _29778_/A VGND VGND VPWR VPWR _35144_/D sky130_fd_sc_hd__clkbuf_1
X_17792_ _17792_/A _17792_/B _17792_/C _17792_/D VGND VGND VPWR VPWR _17793_/A sky130_fd_sc_hd__or4_2
XFILLER_226_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19531_ _19531_/A _19531_/B _19531_/C _19531_/D VGND VGND VPWR VPWR _19532_/A sky130_fd_sc_hd__or4_1
XFILLER_93_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28729_ _26946_/X _34678_/Q _28747_/S VGND VGND VPWR VPWR _28730_/A sky130_fd_sc_hd__mux2_1
X_16743_ _16739_/X _16742_/X _16422_/X VGND VGND VPWR VPWR _16765_/A sky130_fd_sc_hd__o21ba_1
XFILLER_47_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19462_ _19453_/X _19460_/X _19461_/X VGND VGND VPWR VPWR _19463_/D sky130_fd_sc_hd__o21ba_1
X_31740_ _36074_/Q input21/X _31742_/S VGND VGND VPWR VPWR _31741_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16674_ _16349_/X _16672_/X _16673_/X _16355_/X VGND VGND VPWR VPWR _16674_/X sky130_fd_sc_hd__a22o_1
X_18413_ _32719_/Q _32655_/Q _32591_/Q _36047_/Q _20162_/A _20013_/A VGND VGND VPWR
+ VPWR _18413_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31671_ _31671_/A VGND VGND VPWR VPWR _36041_/D sky130_fd_sc_hd__clkbuf_1
X_19393_ _33515_/Q _33451_/Q _33387_/Q _33323_/Q _19070_/X _19071_/X VGND VGND VPWR
+ VPWR _19393_/X sky130_fd_sc_hd__mux4_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33410_ _34050_/CLK _33410_/D VGND VGND VPWR VPWR _33410_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _20155_/A VGND VGND VPWR VPWR _18344_/X sky130_fd_sc_hd__buf_4
X_30622_ _30733_/S VGND VGND VPWR VPWR _30641_/S sky130_fd_sc_hd__buf_4
X_34390_ _34706_/CLK _34390_/D VGND VGND VPWR VPWR _34390_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1063 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33341_ _33789_/CLK _33341_/D VGND VGND VPWR VPWR _33341_/Q sky130_fd_sc_hd__dfxtp_1
X_18275_ input79/X input80/X VGND VGND VPWR VPWR _20061_/A sky130_fd_sc_hd__nor2b_4
X_30553_ _23274_/X _35511_/Q _30569_/S VGND VGND VPWR VPWR _30554_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17226_ _17932_/A VGND VGND VPWR VPWR _17226_/X sky130_fd_sc_hd__buf_4
X_36060_ _36127_/CLK _36060_/D VGND VGND VPWR VPWR _36060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33272_ _36152_/CLK _33272_/D VGND VGND VPWR VPWR _33272_/Q sky130_fd_sc_hd__dfxtp_1
Xinput10 DW[18] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__buf_8
X_30484_ _30484_/A VGND VGND VPWR VPWR _35478_/D sky130_fd_sc_hd__clkbuf_1
Xinput21 DW[28] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__buf_4
XFILLER_128_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput32 DW[38] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__buf_4
X_35011_ _35075_/CLK _35011_/D VGND VGND VPWR VPWR _35011_/Q sky130_fd_sc_hd__dfxtp_1
Xinput43 DW[48] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__buf_6
X_32223_ _35780_/CLK _32223_/D VGND VGND VPWR VPWR _32223_/Q sky130_fd_sc_hd__dfxtp_1
Xinput54 DW[58] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__buf_12
XFILLER_174_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17157_ _17157_/A VGND VGND VPWR VPWR _17157_/X sky130_fd_sc_hd__clkbuf_4
Xinput65 R1[0] VGND VGND VPWR VPWR input65/X sky130_fd_sc_hd__clkbuf_1
Xinput76 R2[5] VGND VGND VPWR VPWR input76/X sky130_fd_sc_hd__buf_2
XFILLER_115_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput87 RW[4] VGND VGND VPWR VPWR input87/X sky130_fd_sc_hd__buf_2
XFILLER_157_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16108_ _17846_/A VGND VGND VPWR VPWR _16108_/X sky130_fd_sc_hd__buf_6
XFILLER_196_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32154_ _33946_/CLK _32154_/D VGND VGND VPWR VPWR _32154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17088_ _33771_/Q _33707_/Q _33643_/Q _33579_/Q _16843_/X _16844_/X VGND VGND VPWR
+ VPWR _17088_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31105_ _35773_/Q _29197_/X _31109_/S VGND VGND VPWR VPWR _31106_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16039_ input69/X VGND VGND VPWR VPWR _17842_/A sky130_fd_sc_hd__buf_12
XFILLER_233_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32085_ _35040_/CLK _32085_/D VGND VGND VPWR VPWR _32085_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_30_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _36194_/CLK sky130_fd_sc_hd__clkbuf_16
X_35913_ _35977_/CLK _35913_/D VGND VGND VPWR VPWR _35913_/Q sky130_fd_sc_hd__dfxtp_1
X_31036_ _35740_/Q _29095_/X _31046_/S VGND VGND VPWR VPWR _31037_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35844_ _35845_/CLK _35844_/D VGND VGND VPWR VPWR _35844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_59__f_CLK clkbuf_5_29_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_59__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_19729_ _33204_/Q _32564_/Q _35956_/Q _35892_/Q _19727_/X _19728_/X VGND VGND VPWR
+ VPWR _19729_/X sky130_fd_sc_hd__mux4_1
XFILLER_211_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35775_ _35837_/CLK _35775_/D VGND VGND VPWR VPWR _35775_/Q sky130_fd_sc_hd__dfxtp_1
X_32987_ _36121_/CLK _32987_/D VGND VGND VPWR VPWR _32987_/Q sky130_fd_sc_hd__dfxtp_1
X_22740_ _35785_/Q _35145_/Q _34505_/Q _33865_/Q _22446_/X _22447_/X VGND VGND VPWR
+ VPWR _22740_/X sky130_fd_sc_hd__mux4_1
X_34726_ _35302_/CLK _34726_/D VGND VGND VPWR VPWR _34726_/Q sky130_fd_sc_hd__dfxtp_1
X_31938_ _23330_/X _36168_/Q _31940_/S VGND VGND VPWR VPWR _31939_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22671_ _22667_/X _22670_/X _22434_/X VGND VGND VPWR VPWR _22693_/A sky130_fd_sc_hd__o21ba_1
XFILLER_198_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34657_ _35098_/CLK _34657_/D VGND VGND VPWR VPWR _34657_/Q sky130_fd_sc_hd__dfxtp_1
X_31869_ _23220_/X _36135_/Q _31877_/S VGND VGND VPWR VPWR _31870_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_97_CLK clkbuf_leaf_99_CLK/A VGND VGND VPWR VPWR _35031_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24410_ input49/X VGND VGND VPWR VPWR _24410_/X sky130_fd_sc_hd__clkbuf_8
X_21622_ _34025_/Q _33961_/Q _33897_/Q _32226_/Q _21620_/X _21621_/X VGND VGND VPWR
+ VPWR _21622_/X sky130_fd_sc_hd__mux4_1
X_33608_ _34817_/CLK _33608_/D VGND VGND VPWR VPWR _33608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_1272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25390_ _25084_/X _33132_/Q _25408_/S VGND VGND VPWR VPWR _25391_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34588_ _34781_/CLK _34588_/D VGND VGND VPWR VPWR _34588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24341_ _24341_/A VGND VGND VPWR VPWR _32684_/D sky130_fd_sc_hd__clkbuf_1
X_21553_ _32743_/Q _32679_/Q _32615_/Q _36071_/Q _21519_/X _21303_/X VGND VGND VPWR
+ VPWR _21553_/X sky130_fd_sc_hd__mux4_1
X_33539_ _34050_/CLK _33539_/D VGND VGND VPWR VPWR _33539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20504_ _18297_/X _20502_/X _20503_/X _18303_/X VGND VGND VPWR VPWR _20504_/X sky130_fd_sc_hd__a22o_1
X_24272_ _24272_/A VGND VGND VPWR VPWR _32662_/D sky130_fd_sc_hd__clkbuf_1
X_27060_ _26878_/X _33888_/Q _27062_/S VGND VGND VPWR VPWR _27061_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21484_ _34021_/Q _33957_/Q _33893_/Q _32182_/Q _21267_/X _21268_/X VGND VGND VPWR
+ VPWR _21484_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26011_ _24989_/X _33422_/Q _26029_/S VGND VGND VPWR VPWR _26012_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23223_ input19/X VGND VGND VPWR VPWR _23223_/X sky130_fd_sc_hd__buf_4
X_35209_ _35273_/CLK _35209_/D VGND VGND VPWR VPWR _35209_/Q sky130_fd_sc_hd__dfxtp_1
X_20435_ _32521_/Q _32393_/Q _32073_/Q _36041_/Q _20282_/X _19307_/A VGND VGND VPWR
+ VPWR _20435_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36189_ _36189_/CLK _36189_/D VGND VGND VPWR VPWR _36189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23154_ _23154_/A VGND VGND VPWR VPWR _32163_/D sky130_fd_sc_hd__clkbuf_1
XTAP_7005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20366_ _34311_/Q _34247_/Q _34183_/Q _34119_/Q _20095_/X _20096_/X VGND VGND VPWR
+ VPWR _20366_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22105_ _22458_/A VGND VGND VPWR VPWR _22105_/X sky130_fd_sc_hd__clkbuf_4
XTAP_7049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27962_ _34315_/Q _24434_/X _27966_/S VGND VGND VPWR VPWR _27963_/A sky130_fd_sc_hd__mux2_1
X_23085_ _23085_/A VGND VGND VPWR VPWR _31275_/A sky130_fd_sc_hd__buf_6
X_20297_ _35332_/Q _35268_/Q _35204_/Q _32324_/Q _20012_/X _20013_/X VGND VGND VPWR
+ VPWR _20297_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_21_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _34779_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29701_ _29701_/A VGND VGND VPWR VPWR _35107_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26913_ _26912_/X _33835_/Q _26913_/S VGND VGND VPWR VPWR _26914_/A sky130_fd_sc_hd__mux2_1
X_22036_ _35060_/Q _34996_/Q _34932_/Q _34868_/Q _21756_/X _21757_/X VGND VGND VPWR
+ VPWR _22036_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27893_ _34282_/Q _24332_/X _27895_/S VGND VGND VPWR VPWR _27894_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29632_ _35075_/Q _29216_/X _29644_/S VGND VGND VPWR VPWR _29633_/A sky130_fd_sc_hd__mux2_1
XTAP_5647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26844_ input62/X VGND VGND VPWR VPWR _26844_/X sky130_fd_sc_hd__buf_4
XFILLER_57_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29563_ _35042_/Q _29113_/X _29581_/S VGND VGND VPWR VPWR _29564_/A sky130_fd_sc_hd__mux2_1
XTAP_4968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26775_ _26775_/A VGND VGND VPWR VPWR _33783_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23987_ _22898_/X _32532_/Q _23993_/S VGND VGND VPWR VPWR _23988_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28514_ _26829_/X _34576_/Q _28528_/S VGND VGND VPWR VPWR _28515_/A sky130_fd_sc_hd__mux2_1
X_25726_ _25726_/A VGND VGND VPWR VPWR _33288_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29494_ _29494_/A VGND VGND VPWR VPWR _35009_/D sky130_fd_sc_hd__clkbuf_1
X_22938_ input11/X VGND VGND VPWR VPWR _22938_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_232_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28445_ _28445_/A VGND VGND VPWR VPWR _34543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25657_ _25657_/A VGND VGND VPWR VPWR _33255_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22869_ _34573_/Q _32461_/Q _34445_/Q _34381_/Q _20663_/X _20665_/X VGND VGND VPWR
+ VPWR _22869_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_88_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _35669_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_73_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24608_ _24608_/A VGND VGND VPWR VPWR _32793_/D sky130_fd_sc_hd__clkbuf_1
XPHY_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16390_ _16386_/X _16389_/X _16011_/X VGND VGND VPWR VPWR _16412_/A sky130_fd_sc_hd__o21ba_2
X_28376_ _28376_/A VGND VGND VPWR VPWR _34510_/D sky130_fd_sc_hd__clkbuf_1
XPHY_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25588_ _25588_/A VGND VGND VPWR VPWR _33224_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27327_ _27327_/A VGND VGND VPWR VPWR _34014_/D sky130_fd_sc_hd__clkbuf_1
XPHY_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24539_ _24539_/A VGND VGND VPWR VPWR _32762_/D sky130_fd_sc_hd__clkbuf_1
XPHY_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18060_ _35078_/Q _35014_/Q _34950_/Q _34886_/Q _17862_/X _17863_/X VGND VGND VPWR
+ VPWR _18060_/X sky130_fd_sc_hd__mux4_1
X_27258_ _26971_/X _33982_/Q _27260_/S VGND VGND VPWR VPWR _27259_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17011_ _35048_/Q _34984_/Q _34920_/Q _34856_/Q _16803_/X _16804_/X VGND VGND VPWR
+ VPWR _17011_/X sky130_fd_sc_hd__mux4_1
X_26209_ _25084_/X _33516_/Q _26227_/S VGND VGND VPWR VPWR _26210_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27189_ _26869_/X _33949_/Q _27197_/S VGND VGND VPWR VPWR _27190_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18962_ _18962_/A VGND VGND VPWR VPWR _32094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_12_CLK clkbuf_6_3__f_CLK/X VGND VGND VPWR VPWR _35803_/CLK sky130_fd_sc_hd__clkbuf_16
X_17913_ _17907_/X _17912_/X _17834_/X VGND VGND VPWR VPWR _17937_/A sky130_fd_sc_hd__o21ba_1
XFILLER_117_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18893_ _33757_/Q _33693_/Q _33629_/Q _33565_/Q _18790_/X _18791_/X VGND VGND VPWR
+ VPWR _18893_/X sky130_fd_sc_hd__mux4_1
XTAP_6860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1095 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17844_ _17838_/X _17841_/X _17842_/X _17843_/X VGND VGND VPWR VPWR _17869_/B sky130_fd_sc_hd__o211a_1
X_32910_ _35982_/CLK _32910_/D VGND VGND VPWR VPWR _32910_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33890_ _34146_/CLK _33890_/D VGND VGND VPWR VPWR _33890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32841_ _36107_/CLK _32841_/D VGND VGND VPWR VPWR _32841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17775_ _17768_/X _17774_/X _17489_/X _17490_/X VGND VGND VPWR VPWR _17792_/B sky130_fd_sc_hd__o211a_1
XFILLER_54_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19514_ _19510_/X _19513_/X _19436_/X _19437_/X VGND VGND VPWR VPWR _19531_/B sky130_fd_sc_hd__o211a_1
X_16726_ _34784_/Q _34720_/Q _34656_/Q _34592_/Q _16582_/X _16583_/X VGND VGND VPWR
+ VPWR _16726_/X sky130_fd_sc_hd__mux4_1
X_32772_ _33026_/CLK _32772_/D VGND VGND VPWR VPWR _32772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35560_ _35819_/CLK _35560_/D VGND VGND VPWR VPWR _35560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34511_ _35728_/CLK _34511_/D VGND VGND VPWR VPWR _34511_/Q sky130_fd_sc_hd__dfxtp_1
X_19445_ _33196_/Q _32556_/Q _35948_/Q _35884_/Q _19374_/X _19375_/X VGND VGND VPWR
+ VPWR _19445_/X sky130_fd_sc_hd__mux4_1
X_31723_ _31813_/S VGND VGND VPWR VPWR _31742_/S sky130_fd_sc_hd__buf_4
X_16657_ _34526_/Q _32414_/Q _34398_/Q _34334_/Q _16519_/X _16520_/X VGND VGND VPWR
+ VPWR _16657_/X sky130_fd_sc_hd__mux4_1
X_35491_ _35552_/CLK _35491_/D VGND VGND VPWR VPWR _35491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_79_CLK clkbuf_leaf_80_CLK/A VGND VGND VPWR VPWR _35925_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34442_ _35787_/CLK _34442_/D VGND VGND VPWR VPWR _34442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31654_ _36033_/Q input47/X _31670_/S VGND VGND VPWR VPWR _31655_/A sky130_fd_sc_hd__mux2_1
X_19376_ _33194_/Q _32554_/Q _35946_/Q _35882_/Q _19374_/X _19375_/X VGND VGND VPWR
+ VPWR _19376_/X sky130_fd_sc_hd__mux4_1
X_16588_ _35036_/Q _34972_/Q _34908_/Q _34844_/Q _16450_/X _16451_/X VGND VGND VPWR
+ VPWR _16588_/X sky130_fd_sc_hd__mux4_1
X_30605_ _30605_/A VGND VGND VPWR VPWR _35535_/D sky130_fd_sc_hd__clkbuf_1
X_18327_ _18357_/A VGND VGND VPWR VPWR _20282_/A sky130_fd_sc_hd__buf_12
X_34373_ _35781_/CLK _34373_/D VGND VGND VPWR VPWR _34373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31585_ _31585_/A VGND VGND VPWR VPWR _36000_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36112_ _36112_/CLK _36112_/D VGND VGND VPWR VPWR _36112_/Q sky130_fd_sc_hd__dfxtp_1
X_33324_ _34292_/CLK _33324_/D VGND VGND VPWR VPWR _33324_/Q sky130_fd_sc_hd__dfxtp_1
X_18258_ _18254_/X _18257_/X _17842_/A _17843_/A VGND VGND VPWR VPWR _18273_/B sky130_fd_sc_hd__o211a_1
XFILLER_148_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_1167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30536_ _23247_/X _35503_/Q _30548_/S VGND VGND VPWR VPWR _30537_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17209_ _33262_/Q _36142_/Q _33134_/Q _33070_/Q _17058_/X _17059_/X VGND VGND VPWR
+ VPWR _17209_/X sky130_fd_sc_hd__mux4_1
X_36043_ _36172_/CLK _36043_/D VGND VGND VPWR VPWR _36043_/Q sky130_fd_sc_hd__dfxtp_1
X_33255_ _33255_/CLK _33255_/D VGND VGND VPWR VPWR _33255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18189_ _34059_/Q _33995_/Q _33931_/Q _32267_/Q _16058_/X _16060_/X VGND VGND VPWR
+ VPWR _18189_/X sky130_fd_sc_hd__mux4_1
X_30467_ _23077_/X _35470_/Q _30485_/S VGND VGND VPWR VPWR _30468_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20220_ _20216_/X _20219_/X _20142_/X _20143_/X VGND VGND VPWR VPWR _20237_/B sky130_fd_sc_hd__o211a_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32206_ _35700_/CLK _32206_/D VGND VGND VPWR VPWR _32206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33186_ _35938_/CLK _33186_/D VGND VGND VPWR VPWR _33186_/Q sky130_fd_sc_hd__dfxtp_1
X_30398_ _30398_/A VGND VGND VPWR VPWR _35437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20151_ _33216_/Q _32576_/Q _35968_/Q _35904_/Q _20080_/X _20081_/X VGND VGND VPWR
+ VPWR _20151_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32137_ _35815_/CLK _32137_/D VGND VGND VPWR VPWR _32137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32068_ _32518_/CLK _32068_/D VGND VGND VPWR VPWR _32068_/Q sky130_fd_sc_hd__dfxtp_1
X_20082_ _33214_/Q _32574_/Q _35966_/Q _35902_/Q _20080_/X _20081_/X VGND VGND VPWR
+ VPWR _20082_/X sky130_fd_sc_hd__mux4_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31019_ _35732_/Q _29070_/X _31025_/S VGND VGND VPWR VPWR _31020_/A sky130_fd_sc_hd__mux2_1
XTAP_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23910_ _22985_/X _32496_/Q _23920_/S VGND VGND VPWR VPWR _23911_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24890_ _24890_/A VGND VGND VPWR VPWR _32926_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23841_ _22883_/X _32463_/Q _23857_/S VGND VGND VPWR VPWR _23842_/A sky130_fd_sc_hd__mux2_1
XTAP_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35827_ _35827_/CLK _35827_/D VGND VGND VPWR VPWR _35827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26560_ _25004_/X _33682_/Q _26570_/S VGND VGND VPWR VPWR _26561_/A sky130_fd_sc_hd__mux2_1
XANTENNA_508 _17900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20984_ _22557_/A VGND VGND VPWR VPWR _20984_/X sky130_fd_sc_hd__buf_4
X_35758_ _35758_/CLK _35758_/D VGND VGND VPWR VPWR _35758_/Q sky130_fd_sc_hd__dfxtp_1
X_23772_ _22982_/X _32431_/Q _23784_/S VGND VGND VPWR VPWR _23773_/A sky130_fd_sc_hd__mux2_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_519 _17970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25511_ _25511_/A VGND VGND VPWR VPWR _33187_/D sky130_fd_sc_hd__clkbuf_1
X_22723_ _22723_/A _22723_/B _22723_/C _22723_/D VGND VGND VPWR VPWR _22724_/A sky130_fd_sc_hd__or4_4
XFILLER_198_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34709_ _36189_/CLK _34709_/D VGND VGND VPWR VPWR _34709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26491_ _25103_/X _33650_/Q _26497_/S VGND VGND VPWR VPWR _26492_/A sky130_fd_sc_hd__mux2_1
X_35689_ _35815_/CLK _35689_/D VGND VGND VPWR VPWR _35689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28230_ _27008_/X _34442_/Q _28236_/S VGND VGND VPWR VPWR _28231_/A sky130_fd_sc_hd__mux2_1
X_25442_ _25162_/X _33157_/Q _25450_/S VGND VGND VPWR VPWR _25443_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22654_ _20597_/X _22652_/X _22653_/X _20603_/X VGND VGND VPWR VPWR _22654_/X sky130_fd_sc_hd__a22o_1
XFILLER_41_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28161_ _26906_/X _34409_/Q _28165_/S VGND VGND VPWR VPWR _28162_/A sky130_fd_sc_hd__mux2_1
X_21605_ _34792_/Q _34728_/Q _34664_/Q _34600_/Q _21535_/X _21536_/X VGND VGND VPWR
+ VPWR _21605_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22585_ _22369_/X _22583_/X _22584_/X _22373_/X VGND VGND VPWR VPWR _22585_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25373_ _25060_/X _33124_/Q _25387_/S VGND VGND VPWR VPWR _25374_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27112_ _27112_/A VGND VGND VPWR VPWR _33912_/D sky130_fd_sc_hd__clkbuf_1
X_24324_ _32679_/Q _24323_/X _24336_/S VGND VGND VPWR VPWR _24325_/A sky130_fd_sc_hd__mux2_1
X_28092_ _28092_/A VGND VGND VPWR VPWR _34376_/D sky130_fd_sc_hd__clkbuf_1
X_21536_ _22595_/A VGND VGND VPWR VPWR _21536_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_194_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27043_ _27154_/S VGND VGND VPWR VPWR _27062_/S sky130_fd_sc_hd__buf_6
XFILLER_166_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24255_ input34/X VGND VGND VPWR VPWR _24255_/X sky130_fd_sc_hd__buf_6
X_21467_ _21246_/X _21465_/X _21466_/X _21249_/X VGND VGND VPWR VPWR _21467_/X sky130_fd_sc_hd__a22o_1
XFILLER_181_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20418_ _20155_/X _20416_/X _20417_/X _20158_/X VGND VGND VPWR VPWR _20418_/X sky130_fd_sc_hd__a22o_1
X_23206_ _32185_/Q _23145_/X _23206_/S VGND VGND VPWR VPWR _23207_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24186_ _22991_/X _32626_/Q _24192_/S VGND VGND VPWR VPWR _24187_/A sky130_fd_sc_hd__mux2_1
X_21398_ _35298_/Q _35234_/Q _35170_/Q _32290_/Q _21253_/X _21254_/X VGND VGND VPWR
+ VPWR _21398_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20349_ _35846_/Q _32225_/Q _35718_/Q _35654_/Q _18289_/X _18291_/X VGND VGND VPWR
+ VPWR _20349_/X sky130_fd_sc_hd__mux4_1
X_23137_ _32158_/Q _23136_/X _23146_/S VGND VGND VPWR VPWR _23138_/A sky130_fd_sc_hd__mux2_1
XTAP_6101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28994_ _34804_/Q _24363_/X _28996_/S VGND VGND VPWR VPWR _28995_/A sky130_fd_sc_hd__mux2_1
XTAP_6112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27945_ _27945_/A VGND VGND VPWR VPWR _34306_/D sky130_fd_sc_hd__clkbuf_1
X_23068_ input58/X VGND VGND VPWR VPWR _23068_/X sky130_fd_sc_hd__buf_2
XTAP_5400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22019_ _33012_/Q _32948_/Q _32884_/Q _32820_/Q _21942_/X _21943_/X VGND VGND VPWR
+ VPWR _22019_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27876_ _27966_/S VGND VGND VPWR VPWR _27895_/S sky130_fd_sc_hd__buf_4
XTAP_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26827_ _26826_/X _33807_/Q _26851_/S VGND VGND VPWR VPWR _26828_/A sky130_fd_sc_hd__mux2_1
XTAP_5488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29615_ _35067_/Q _29191_/X _29623_/S VGND VGND VPWR VPWR _29616_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_42__f_CLK clkbuf_5_21_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_42__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_63_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ _17554_/X _17559_/X _17481_/X VGND VGND VPWR VPWR _17584_/A sky130_fd_sc_hd__o21ba_1
X_29546_ _35034_/Q _29089_/X _29560_/S VGND VGND VPWR VPWR _29547_/A sky130_fd_sc_hd__mux2_1
XTAP_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26758_ _26758_/A VGND VGND VPWR VPWR _33775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16511_ _16288_/X _16509_/X _16510_/X _16291_/X VGND VGND VPWR VPWR _16511_/X sky130_fd_sc_hd__a22o_1
XFILLER_84_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25709_ _33280_/Q _24400_/X _25727_/S VGND VGND VPWR VPWR _25710_/A sky130_fd_sc_hd__mux2_1
X_29477_ _29477_/A VGND VGND VPWR VPWR _35001_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17491_ _17485_/X _17488_/X _17489_/X _17490_/X VGND VGND VPWR VPWR _17516_/B sky130_fd_sc_hd__o211a_1
X_26689_ _26689_/A VGND VGND VPWR VPWR _33742_/D sky130_fd_sc_hd__clkbuf_1
X_19230_ _18941_/X _19228_/X _19229_/X _18944_/X VGND VGND VPWR VPWR _19230_/X sky130_fd_sc_hd__a22o_1
XFILLER_44_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28428_ _28428_/A VGND VGND VPWR VPWR _34535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16442_ _16437_/X _16440_/X _16441_/X VGND VGND VPWR VPWR _16457_/C sky130_fd_sc_hd__o21ba_1
XFILLER_147_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _35166_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19161_ _19157_/X _19160_/X _19083_/X _19084_/X VGND VGND VPWR VPWR _19178_/B sky130_fd_sc_hd__o211a_1
X_28359_ _34503_/Q _24422_/X _28363_/S VGND VGND VPWR VPWR _28360_/A sky130_fd_sc_hd__mux2_1
X_16373_ _34774_/Q _34710_/Q _34646_/Q _34582_/Q _16229_/X _16230_/X VGND VGND VPWR
+ VPWR _16373_/X sky130_fd_sc_hd__mux4_1
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18112_ _35592_/Q _35528_/Q _35464_/Q _35400_/Q _17956_/X _17957_/X VGND VGND VPWR
+ VPWR _18112_/X sky130_fd_sc_hd__mux4_1
XFILLER_160_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31370_ _31370_/A VGND VGND VPWR VPWR _35898_/D sky130_fd_sc_hd__clkbuf_1
X_19092_ _33186_/Q _32546_/Q _35938_/Q _35874_/Q _19021_/X _19022_/X VGND VGND VPWR
+ VPWR _19092_/X sky130_fd_sc_hd__mux4_1
XFILLER_8_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1099 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30321_ _35402_/Q _29237_/X _30327_/S VGND VGND VPWR VPWR _30322_/A sky130_fd_sc_hd__mux2_1
X_18043_ _33286_/Q _36166_/Q _33158_/Q _33094_/Q _17764_/X _17765_/X VGND VGND VPWR
+ VPWR _18043_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33040_ _36114_/CLK _33040_/D VGND VGND VPWR VPWR _33040_/Q sky130_fd_sc_hd__dfxtp_1
X_30252_ _35369_/Q _29135_/X _30256_/S VGND VGND VPWR VPWR _30253_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30183_ _30183_/A VGND VGND VPWR VPWR _35336_/D sky130_fd_sc_hd__clkbuf_1
X_19994_ _32508_/Q _32380_/Q _32060_/Q _36028_/Q _19929_/X _19717_/X VGND VGND VPWR
+ VPWR _19994_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18945_ _18941_/X _18942_/X _18943_/X _18944_/X VGND VGND VPWR VPWR _18945_/X sky130_fd_sc_hd__a22o_1
X_34991_ _35758_/CLK _34991_/D VGND VGND VPWR VPWR _34991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33942_ _34006_/CLK _33942_/D VGND VGND VPWR VPWR _33942_/Q sky130_fd_sc_hd__dfxtp_1
X_18876_ _35740_/Q _35100_/Q _34460_/Q _33820_/Q _18734_/X _18735_/X VGND VGND VPWR
+ VPWR _18876_/X sky130_fd_sc_hd__mux4_1
XTAP_6690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17827_ _34304_/Q _34240_/Q _34176_/Q _34112_/Q _17795_/X _17796_/X VGND VGND VPWR
+ VPWR _17827_/X sky130_fd_sc_hd__mux4_1
X_33873_ _36228_/CLK _33873_/D VGND VGND VPWR VPWR _33873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35612_ _35803_/CLK _35612_/D VGND VGND VPWR VPWR _35612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32824_ _36025_/CLK _32824_/D VGND VGND VPWR VPWR _32824_/Q sky130_fd_sc_hd__dfxtp_1
X_17758_ _34046_/Q _33982_/Q _33918_/Q _32254_/Q _17726_/X _17727_/X VGND VGND VPWR
+ VPWR _17758_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35543_ _35797_/CLK _35543_/D VGND VGND VPWR VPWR _35543_/Q sky130_fd_sc_hd__dfxtp_1
X_16709_ _16702_/X _16704_/X _16707_/X _16708_/X VGND VGND VPWR VPWR _16709_/X sky130_fd_sc_hd__a22o_1
X_17689_ _17555_/X _17687_/X _17688_/X _17558_/X VGND VGND VPWR VPWR _17689_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32755_ _36018_/CLK _32755_/D VGND VGND VPWR VPWR _32755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31706_ _31706_/A VGND VGND VPWR VPWR _36057_/D sky130_fd_sc_hd__clkbuf_1
X_19428_ _20134_/A VGND VGND VPWR VPWR _19428_/X sky130_fd_sc_hd__clkbuf_4
X_35474_ _35922_/CLK _35474_/D VGND VGND VPWR VPWR _35474_/Q sky130_fd_sc_hd__dfxtp_1
X_32686_ _36078_/CLK _32686_/D VGND VGND VPWR VPWR _32686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34425_ _35577_/CLK _34425_/D VGND VGND VPWR VPWR _34425_/Q sky130_fd_sc_hd__dfxtp_1
X_31637_ _36025_/Q input38/X _31649_/S VGND VGND VPWR VPWR _31638_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19359_ _20070_/A VGND VGND VPWR VPWR _19359_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22370_ _22370_/A VGND VGND VPWR VPWR _22370_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_241_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31568_ _35992_/Q input2/X _31586_/S VGND VGND VPWR VPWR _31569_/A sky130_fd_sc_hd__mux2_1
X_34356_ _35250_/CLK _34356_/D VGND VGND VPWR VPWR _34356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21321_ _22531_/A VGND VGND VPWR VPWR _21321_/X sky130_fd_sc_hd__buf_6
X_33307_ _36194_/CLK _33307_/D VGND VGND VPWR VPWR _33307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30519_ _23220_/X _35495_/Q _30527_/S VGND VGND VPWR VPWR _30520_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34287_ _34288_/CLK _34287_/D VGND VGND VPWR VPWR _34287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31499_ _31499_/A VGND VGND VPWR VPWR _35959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36026_ _36027_/CLK _36026_/D VGND VGND VPWR VPWR _36026_/Q sky130_fd_sc_hd__dfxtp_1
X_33238_ _36119_/CLK _33238_/D VGND VGND VPWR VPWR _33238_/Q sky130_fd_sc_hd__dfxtp_1
X_24040_ _22976_/X _32557_/Q _24056_/S VGND VGND VPWR VPWR _24041_/A sky130_fd_sc_hd__mux2_1
X_21252_ _34782_/Q _34718_/Q _34654_/Q _34590_/Q _21182_/X _21183_/X VGND VGND VPWR
+ VPWR _21252_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20203_ _20203_/A VGND VGND VPWR VPWR _20203_/X sky130_fd_sc_hd__buf_6
XFILLER_190_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33169_ _36112_/CLK _33169_/D VGND VGND VPWR VPWR _33169_/Q sky130_fd_sc_hd__dfxtp_1
X_21183_ _22595_/A VGND VGND VPWR VPWR _21183_/X sky130_fd_sc_hd__buf_4
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20134_ _20134_/A VGND VGND VPWR VPWR _20134_/X sky130_fd_sc_hd__buf_2
X_25991_ _25162_/X _33413_/Q _25999_/S VGND VGND VPWR VPWR _25992_/A sky130_fd_sc_hd__mux2_1
X_27730_ _27730_/A VGND VGND VPWR VPWR _34204_/D sky130_fd_sc_hd__clkbuf_1
X_20065_ _20070_/A VGND VGND VPWR VPWR _20065_/X sky130_fd_sc_hd__clkbuf_4
X_24942_ _23007_/X _32951_/Q _24958_/S VGND VGND VPWR VPWR _24943_/A sky130_fd_sc_hd__mux2_1
XTAP_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27661_ _34172_/Q _24388_/X _27667_/S VGND VGND VPWR VPWR _27662_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24873_ _24873_/A VGND VGND VPWR VPWR _32918_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29400_ _23108_/X _34965_/Q _29404_/S VGND VGND VPWR VPWR _29401_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26612_ _25081_/X _33707_/Q _26612_/S VGND VGND VPWR VPWR _26613_/A sky130_fd_sc_hd__mux2_1
XTAP_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23824_ _23059_/X _32456_/Q _23826_/S VGND VGND VPWR VPWR _23825_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27592_ _34139_/Q _24286_/X _27604_/S VGND VGND VPWR VPWR _27593_/A sky130_fd_sc_hd__mux2_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_305 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_316 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_327 _32141_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29331_ _29331_/A VGND VGND VPWR VPWR _34932_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26543_ _25180_/X _33675_/Q _26547_/S VGND VGND VPWR VPWR _26544_/A sky130_fd_sc_hd__mux2_1
XANTENNA_338 _36205_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23755_ _22957_/X _32423_/Q _23763_/S VGND VGND VPWR VPWR _23756_/A sky130_fd_sc_hd__mux2_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_349 _36205_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20967_ _35542_/Q _35478_/Q _35414_/Q _35350_/Q _20791_/X _20792_/X VGND VGND VPWR
+ VPWR _20967_/X sky130_fd_sc_hd__mux4_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22706_ _33032_/Q _32968_/Q _32904_/Q _32840_/Q _20580_/X _20583_/X VGND VGND VPWR
+ VPWR _22706_/X sky130_fd_sc_hd__mux4_1
X_29262_ _29262_/A VGND VGND VPWR VPWR _34899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26474_ _25078_/X _33642_/Q _26476_/S VGND VGND VPWR VPWR _26475_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23686_ _32392_/Q _23330_/X _23688_/S VGND VGND VPWR VPWR _23687_/A sky130_fd_sc_hd__mux2_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ _20892_/X _20897_/X _20671_/X VGND VGND VPWR VPWR _20908_/C sky130_fd_sc_hd__o21ba_1
X_28213_ _28213_/A VGND VGND VPWR VPWR _34433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25425_ _25137_/X _33149_/Q _25429_/S VGND VGND VPWR VPWR _25426_/A sky130_fd_sc_hd__mux2_1
X_22637_ _22501_/X _22635_/X _22636_/X _22506_/X VGND VGND VPWR VPWR _22637_/X sky130_fd_sc_hd__a22o_1
XFILLER_224_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29193_ _29193_/A VGND VGND VPWR VPWR _34875_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28144_ _26881_/X _34401_/Q _28144_/S VGND VGND VPWR VPWR _28145_/A sky130_fd_sc_hd__mux2_1
X_25356_ _25035_/X _33116_/Q _25366_/S VGND VGND VPWR VPWR _25357_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22568_ _22564_/X _22567_/X _22467_/X VGND VGND VPWR VPWR _22569_/D sky130_fd_sc_hd__o21ba_1
XFILLER_194_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24307_ input13/X VGND VGND VPWR VPWR _24307_/X sky130_fd_sc_hd__buf_4
X_28075_ _26977_/X _34368_/Q _28093_/S VGND VGND VPWR VPWR _28076_/A sky130_fd_sc_hd__mux2_1
X_21519_ _22578_/A VGND VGND VPWR VPWR _21519_/X sky130_fd_sc_hd__buf_6
X_25287_ _25134_/X _33084_/Q _25293_/S VGND VGND VPWR VPWR _25288_/A sky130_fd_sc_hd__mux2_1
X_22499_ _22499_/A _22499_/B _22499_/C _22499_/D VGND VGND VPWR VPWR _22500_/A sky130_fd_sc_hd__or4_4
XFILLER_119_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27026_ _27026_/A VGND VGND VPWR VPWR _33871_/D sky130_fd_sc_hd__clkbuf_1
X_24238_ _23068_/X _32651_/Q _24242_/S VGND VGND VPWR VPWR _24239_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24169_ _22966_/X _32618_/Q _24171_/S VGND VGND VPWR VPWR _24170_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16991_ _33000_/Q _32936_/Q _32872_/Q _32808_/Q _16989_/X _16990_/X VGND VGND VPWR
+ VPWR _16991_/X sky130_fd_sc_hd__mux4_1
XFILLER_205_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28977_ _28998_/A VGND VGND VPWR VPWR _28996_/S sky130_fd_sc_hd__buf_4
XFILLER_122_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18730_ _20142_/A VGND VGND VPWR VPWR _18730_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_77_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27928_ _27928_/A VGND VGND VPWR VPWR _34298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18661_ _20211_/A VGND VGND VPWR VPWR _18661_/X sky130_fd_sc_hd__buf_4
XFILLER_62_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27859_ _27859_/A VGND VGND VPWR VPWR _34265_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17612_ _34553_/Q _32441_/Q _34425_/Q _34361_/Q _17578_/X _17579_/X VGND VGND VPWR
+ VPWR _17612_/X sky130_fd_sc_hd__mux4_1
X_30870_ _31140_/A _30870_/B VGND VGND VPWR VPWR _31003_/S sky130_fd_sc_hd__nor2_8
XTAP_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18592_ _18588_/X _18589_/X _18590_/X _18591_/X VGND VGND VPWR VPWR _18592_/X sky130_fd_sc_hd__a22o_1
XTAP_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17543_ _35063_/Q _34999_/Q _34935_/Q _34871_/Q _17509_/X _17510_/X VGND VGND VPWR
+ VPWR _17543_/X sky130_fd_sc_hd__mux4_1
X_29529_ _35026_/Q _29064_/X _29539_/S VGND VGND VPWR VPWR _29530_/A sky130_fd_sc_hd__mux2_1
XTAP_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_850 _24401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32540_ _35928_/CLK _32540_/D VGND VGND VPWR VPWR _32540_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_861 _24366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_872 _24987_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17474_ _34294_/Q _34230_/Q _34166_/Q _34102_/Q _17442_/X _17443_/X VGND VGND VPWR
+ VPWR _17474_/X sky130_fd_sc_hd__mux4_1
XANTENNA_883 _25084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_894 _25735_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16425_ _33240_/Q _36120_/Q _33112_/Q _33048_/Q _16352_/X _16353_/X VGND VGND VPWR
+ VPWR _16425_/X sky130_fd_sc_hd__mux4_1
X_19213_ _34278_/Q _34214_/Q _34150_/Q _34086_/Q _19036_/X _19037_/X VGND VGND VPWR
+ VPWR _19213_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32471_ _35991_/CLK _32471_/D VGND VGND VPWR VPWR _32471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31422_ _23102_/X _35923_/Q _31430_/S VGND VGND VPWR VPWR _31423_/A sky130_fd_sc_hd__mux2_1
X_19144_ _20203_/A VGND VGND VPWR VPWR _19144_/X sky130_fd_sc_hd__clkbuf_4
X_34210_ _35992_/CLK _34210_/D VGND VGND VPWR VPWR _34210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16356_ _16349_/X _16351_/X _16354_/X _16355_/X VGND VGND VPWR VPWR _16356_/X sky130_fd_sc_hd__a22o_1
X_35190_ _35319_/CLK _35190_/D VGND VGND VPWR VPWR _35190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34141_ _34142_/CLK _34141_/D VGND VGND VPWR VPWR _34141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31353_ _31353_/A VGND VGND VPWR VPWR _35890_/D sky130_fd_sc_hd__clkbuf_1
X_19075_ _20134_/A VGND VGND VPWR VPWR _19075_/X sky130_fd_sc_hd__buf_2
X_16287_ _16281_/X _16286_/X _16040_/X _16042_/X VGND VGND VPWR VPWR _16308_/B sky130_fd_sc_hd__o211a_1
XFILLER_121_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18026_ _34821_/Q _34757_/Q _34693_/Q _34629_/Q _17994_/X _17995_/X VGND VGND VPWR
+ VPWR _18026_/X sky130_fd_sc_hd__mux4_1
X_30304_ _30304_/A VGND VGND VPWR VPWR _35393_/D sky130_fd_sc_hd__clkbuf_1
X_34072_ _34266_/CLK _34072_/D VGND VGND VPWR VPWR _34072_/Q sky130_fd_sc_hd__dfxtp_1
X_31284_ _31284_/A VGND VGND VPWR VPWR _35857_/D sky130_fd_sc_hd__clkbuf_1
X_33023_ _36097_/CLK _33023_/D VGND VGND VPWR VPWR _33023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30235_ _35361_/Q _29110_/X _30235_/S VGND VGND VPWR VPWR _30236_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30166_ _35328_/Q _29206_/X _30184_/S VGND VGND VPWR VPWR _30167_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19977_ _19802_/X _19975_/X _19976_/X _19805_/X VGND VGND VPWR VPWR _19977_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18928_ _33502_/Q _33438_/Q _33374_/Q _33310_/Q _18717_/X _18718_/X VGND VGND VPWR
+ VPWR _18928_/X sky130_fd_sc_hd__mux4_1
X_30097_ _30097_/A VGND VGND VPWR VPWR _35295_/D sky130_fd_sc_hd__clkbuf_1
X_34974_ _35038_/CLK _34974_/D VGND VGND VPWR VPWR _34974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1260 _28506_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1271 _31003_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1282 _17830_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33925_ _34057_/CLK _33925_/D VGND VGND VPWR VPWR _33925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1293 _17932_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18859_ _33756_/Q _33692_/Q _33628_/Q _33564_/Q _18790_/X _18791_/X VGND VGND VPWR
+ VPWR _18859_/X sky130_fd_sc_hd__mux4_1
X_33856_ _35777_/CLK _33856_/D VGND VGND VPWR VPWR _33856_/Q sky130_fd_sc_hd__dfxtp_1
X_21870_ _21802_/X _21868_/X _21869_/X _21805_/X VGND VGND VPWR VPWR _21870_/X sky130_fd_sc_hd__a22o_1
X_20821_ _20816_/X _20820_/X _20640_/X _20642_/X VGND VGND VPWR VPWR _20838_/B sky130_fd_sc_hd__o211a_1
X_32807_ _36007_/CLK _32807_/D VGND VGND VPWR VPWR _32807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30999_ _35723_/Q _29240_/X _31003_/S VGND VGND VPWR VPWR _31000_/A sky130_fd_sc_hd__mux2_1
X_33787_ _33787_/CLK _33787_/D VGND VGND VPWR VPWR _33787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23540_ _23540_/A VGND VGND VPWR VPWR _32323_/D sky130_fd_sc_hd__clkbuf_1
X_35526_ _35975_/CLK _35526_/D VGND VGND VPWR VPWR _35526_/Q sky130_fd_sc_hd__dfxtp_1
X_20752_ _32464_/Q _32336_/Q _32016_/Q _35984_/Q _20628_/X _22463_/A VGND VGND VPWR
+ VPWR _20752_/X sky130_fd_sc_hd__mux4_1
X_32738_ _36067_/CLK _32738_/D VGND VGND VPWR VPWR _32738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35457_ _35585_/CLK _35457_/D VGND VGND VPWR VPWR _35457_/Q sky130_fd_sc_hd__dfxtp_1
X_20683_ _22367_/A VGND VGND VPWR VPWR _21752_/A sky130_fd_sc_hd__buf_12
X_23471_ _23471_/A VGND VGND VPWR VPWR _32290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32669_ _36127_/CLK _32669_/D VGND VGND VPWR VPWR _32669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25210_ _25210_/A VGND VGND VPWR VPWR _33047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22422_ _22107_/X _22420_/X _22421_/X _22112_/X VGND VGND VPWR VPWR _22422_/X sky130_fd_sc_hd__a22o_1
X_34408_ _34922_/CLK _34408_/D VGND VGND VPWR VPWR _34408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26190_ _25057_/X _33507_/Q _26206_/S VGND VGND VPWR VPWR _26191_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35388_ _35517_/CLK _35388_/D VGND VGND VPWR VPWR _35388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25141_ _25140_/X _33022_/Q _25144_/S VGND VGND VPWR VPWR _25142_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22353_ _22353_/A VGND VGND VPWR VPWR _36221_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34339_ _35932_/CLK _34339_/D VGND VGND VPWR VPWR _34339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_6__f_CLK clkbuf_5_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_6__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_21304_ _32736_/Q _32672_/Q _32608_/Q _36064_/Q _21166_/X _21303_/X VGND VGND VPWR
+ VPWR _21304_/X sky130_fd_sc_hd__mux4_1
X_22284_ _33788_/Q _33724_/Q _33660_/Q _33596_/Q _22149_/X _22150_/X VGND VGND VPWR
+ VPWR _22284_/X sky130_fd_sc_hd__mux4_1
X_25072_ input19/X VGND VGND VPWR VPWR _25072_/X sky130_fd_sc_hd__buf_2
X_28900_ _28900_/A VGND VGND VPWR VPWR _34759_/D sky130_fd_sc_hd__clkbuf_1
X_24023_ _22951_/X _32549_/Q _24035_/S VGND VGND VPWR VPWR _24024_/A sky130_fd_sc_hd__mux2_1
X_36009_ _36009_/CLK _36009_/D VGND VGND VPWR VPWR _36009_/Q sky130_fd_sc_hd__dfxtp_1
X_21235_ _32478_/Q _32350_/Q _32030_/Q _35998_/Q _21170_/X _20958_/X VGND VGND VPWR
+ VPWR _21235_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29880_ _29880_/A VGND VGND VPWR VPWR _35192_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28831_ _28831_/A VGND VGND VPWR VPWR _34726_/D sky130_fd_sc_hd__clkbuf_1
X_21166_ _22578_/A VGND VGND VPWR VPWR _21166_/X sky130_fd_sc_hd__buf_6
X_20117_ _34815_/Q _34751_/Q _34687_/Q _34623_/Q _19941_/X _19942_/X VGND VGND VPWR
+ VPWR _20117_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28762_ _26996_/X _34694_/Q _28768_/S VGND VGND VPWR VPWR _28763_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25974_ _25137_/X _33405_/Q _25978_/S VGND VGND VPWR VPWR _25975_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21097_ _33498_/Q _33434_/Q _33370_/Q _33306_/Q _21017_/X _21018_/X VGND VGND VPWR
+ VPWR _21097_/X sky130_fd_sc_hd__mux4_1
XFILLER_115_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27713_ _27713_/A VGND VGND VPWR VPWR _34196_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20048_ _34557_/Q _32445_/Q _34429_/Q _34365_/Q _19878_/X _19879_/X VGND VGND VPWR
+ VPWR _20048_/X sky130_fd_sc_hd__mux4_1
X_24925_ _22982_/X _32943_/Q _24937_/S VGND VGND VPWR VPWR _24926_/A sky130_fd_sc_hd__mux2_1
X_28693_ _26894_/X _34661_/Q _28705_/S VGND VGND VPWR VPWR _28694_/A sky130_fd_sc_hd__mux2_1
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27644_ _34164_/Q _24363_/X _27646_/S VGND VGND VPWR VPWR _27645_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24856_ _22875_/X _32910_/Q _24874_/S VGND VGND VPWR VPWR _24857_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23807_ _23834_/S VGND VGND VPWR VPWR _23826_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_22_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_113 _32129_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27575_ _34131_/Q _24261_/X _27583_/S VGND VGND VPWR VPWR _27576_/A sky130_fd_sc_hd__mux2_1
XANTENNA_124 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24787_ _24787_/A VGND VGND VPWR VPWR _32877_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21999_ _21999_/A _21999_/B _21999_/C _21999_/D VGND VGND VPWR VPWR _22000_/A sky130_fd_sc_hd__or4_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_157 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29314_ _23237_/X _34924_/Q _29332_/S VGND VGND VPWR VPWR _29315_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26526_ _26526_/A VGND VGND VPWR VPWR _33666_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23738_ _22932_/X _32415_/Q _23742_/S VGND VGND VPWR VPWR _23739_/A sky130_fd_sc_hd__mux2_1
XANTENNA_168 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_179 _32134_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29245_ _29245_/A VGND VGND VPWR VPWR _34892_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26457_ _26547_/S VGND VGND VPWR VPWR _26476_/S sky130_fd_sc_hd__buf_4
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23669_ _23696_/S VGND VGND VPWR VPWR _23688_/S sky130_fd_sc_hd__clkbuf_8
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _34002_/Q _33938_/Q _33874_/Q _32146_/Q _16108_/X _16109_/X VGND VGND VPWR
+ VPWR _16210_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25408_ _25112_/X _33141_/Q _25408_/S VGND VGND VPWR VPWR _25409_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29176_ _29247_/S VGND VGND VPWR VPWR _29204_/S sky130_fd_sc_hd__buf_4
X_17190_ _35053_/Q _34989_/Q _34925_/Q _34861_/Q _17156_/X _17157_/X VGND VGND VPWR
+ VPWR _17190_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_1014 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26388_ _25150_/X _33601_/Q _26404_/S VGND VGND VPWR VPWR _26389_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16141_ _17858_/A VGND VGND VPWR VPWR _16141_/X sky130_fd_sc_hd__buf_4
XFILLER_31_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28127_ _28127_/A VGND VGND VPWR VPWR _34392_/D sky130_fd_sc_hd__clkbuf_1
X_25339_ _25010_/X _33108_/Q _25345_/S VGND VGND VPWR VPWR _25340_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16072_ _16055_/X _16069_/X _16071_/X VGND VGND VPWR VPWR _16102_/C sky130_fd_sc_hd__o21ba_1
XFILLER_155_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28058_ _26953_/X _34360_/Q _28072_/S VGND VGND VPWR VPWR _28059_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27009_ _27008_/X _33866_/Q _27018_/S VGND VGND VPWR VPWR _27010_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19900_ _35833_/Q _32211_/Q _35705_/Q _35641_/Q _19613_/X _19614_/X VGND VGND VPWR
+ VPWR _19900_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30020_ _35259_/Q _29191_/X _30028_/S VGND VGND VPWR VPWR _30021_/A sky130_fd_sc_hd__mux2_1
X_19831_ _19827_/X _19830_/X _19789_/X _19790_/X VGND VGND VPWR VPWR _19846_/B sky130_fd_sc_hd__o211a_1
XFILLER_29_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19762_ _19652_/X _19760_/X _19761_/X _19655_/X VGND VGND VPWR VPWR _19762_/X sky130_fd_sc_hd__a22o_1
XFILLER_231_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16974_ _16801_/X _16972_/X _16973_/X _16806_/X VGND VGND VPWR VPWR _16974_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18713_ _18713_/A VGND VGND VPWR VPWR _32087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_209_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31971_ _34970_/CLK _31971_/D VGND VGND VPWR VPWR _31971_/Q sky130_fd_sc_hd__dfxtp_1
X_19693_ _35315_/Q _35251_/Q _35187_/Q _32307_/Q _19659_/X _19660_/X VGND VGND VPWR
+ VPWR _19693_/X sky130_fd_sc_hd__mux4_1
XTAP_5082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 DW[16] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_292_CLK clkbuf_6_57__f_CLK/X VGND VGND VPWR VPWR _36033_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_5093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33710_ _34288_/CLK _33710_/D VGND VGND VPWR VPWR _33710_/Q sky130_fd_sc_hd__dfxtp_1
X_18644_ _18436_/X _18642_/X _18643_/X _18441_/X VGND VGND VPWR VPWR _18644_/X sky130_fd_sc_hd__a22o_1
X_30922_ _35686_/Q _29126_/X _30932_/S VGND VGND VPWR VPWR _30923_/A sky130_fd_sc_hd__mux2_1
X_34690_ _35331_/CLK _34690_/D VGND VGND VPWR VPWR _34690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30853_ _30853_/A VGND VGND VPWR VPWR _35653_/D sky130_fd_sc_hd__clkbuf_1
X_33641_ _34870_/CLK _33641_/D VGND VGND VPWR VPWR _33641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18575_ _33492_/Q _33428_/Q _33364_/Q _33300_/Q _18298_/X _18299_/X VGND VGND VPWR
+ VPWR _18575_/X sky130_fd_sc_hd__mux4_1
XTAP_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17526_ _33271_/Q _36151_/Q _33143_/Q _33079_/Q _17411_/X _17412_/X VGND VGND VPWR
+ VPWR _17526_/X sky130_fd_sc_hd__mux4_1
X_33572_ _33702_/CLK _33572_/D VGND VGND VPWR VPWR _33572_/Q sky130_fd_sc_hd__dfxtp_1
X_30784_ _30784_/A VGND VGND VPWR VPWR _35620_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_680 _22557_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_691 _22595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35311_ _35564_/CLK _35311_/D VGND VGND VPWR VPWR _35311_/Q sky130_fd_sc_hd__dfxtp_1
X_32523_ _36171_/CLK _32523_/D VGND VGND VPWR VPWR _32523_/Q sky130_fd_sc_hd__dfxtp_1
X_17457_ _35829_/Q _32207_/Q _35701_/Q _35637_/Q _17313_/X _17314_/X VGND VGND VPWR
+ VPWR _17457_/X sky130_fd_sc_hd__mux4_1
X_16408_ _34519_/Q _32407_/Q _34391_/Q _34327_/Q _16166_/X _16167_/X VGND VGND VPWR
+ VPWR _16408_/X sky130_fd_sc_hd__mux4_1
XFILLER_242_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35242_ _35242_/CLK _35242_/D VGND VGND VPWR VPWR _35242_/Q sky130_fd_sc_hd__dfxtp_1
X_32454_ _35078_/CLK _32454_/D VGND VGND VPWR VPWR _32454_/Q sky130_fd_sc_hd__dfxtp_1
X_17388_ _35571_/Q _35507_/Q _35443_/Q _35379_/Q _17250_/X _17251_/X VGND VGND VPWR
+ VPWR _17388_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31405_ _31405_/A VGND VGND VPWR VPWR _35915_/D sky130_fd_sc_hd__clkbuf_1
X_16339_ _16335_/X _16338_/X _16100_/X VGND VGND VPWR VPWR _16340_/D sky130_fd_sc_hd__o21ba_1
X_19127_ _35747_/Q _35107_/Q _34467_/Q _33827_/Q _19087_/X _19088_/X VGND VGND VPWR
+ VPWR _19127_/X sky130_fd_sc_hd__mux4_1
X_32385_ _36032_/CLK _32385_/D VGND VGND VPWR VPWR _32385_/Q sky130_fd_sc_hd__dfxtp_1
X_35173_ _36004_/CLK _35173_/D VGND VGND VPWR VPWR _35173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34124_ _34124_/CLK _34124_/D VGND VGND VPWR VPWR _34124_/Q sky130_fd_sc_hd__dfxtp_1
X_31336_ _31336_/A VGND VGND VPWR VPWR _35882_/D sky130_fd_sc_hd__clkbuf_1
X_19058_ _34785_/Q _34721_/Q _34657_/Q _34593_/Q _18882_/X _18883_/X VGND VGND VPWR
+ VPWR _19058_/X sky130_fd_sc_hd__mux4_1
XFILLER_161_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18009_ _34053_/Q _33989_/Q _33925_/Q _32261_/Q _17726_/X _17727_/X VGND VGND VPWR
+ VPWR _18009_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34055_ _34816_/CLK _34055_/D VGND VGND VPWR VPWR _34055_/Q sky130_fd_sc_hd__dfxtp_1
X_31267_ _35850_/Q input57/X _31273_/S VGND VGND VPWR VPWR _31268_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21020_ _34008_/Q _33944_/Q _33880_/Q _32152_/Q _20914_/X _20915_/X VGND VGND VPWR
+ VPWR _21020_/X sky130_fd_sc_hd__mux4_1
XFILLER_236_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33006_ _33007_/CLK _33006_/D VGND VGND VPWR VPWR _33006_/Q sky130_fd_sc_hd__dfxtp_1
X_30218_ _30218_/A VGND VGND VPWR VPWR _35352_/D sky130_fd_sc_hd__clkbuf_1
X_31198_ _35817_/Q input20/X _31202_/S VGND VGND VPWR VPWR _31199_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_1076 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30149_ _35320_/Q _29182_/X _30163_/S VGND VGND VPWR VPWR _30150_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34957_ _35021_/CLK _34957_/D VGND VGND VPWR VPWR _34957_/Q sky130_fd_sc_hd__dfxtp_1
X_22971_ _22971_/A VGND VGND VPWR VPWR _32043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1090 _17232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_283_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _36090_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24710_ _24710_/A VGND VGND VPWR VPWR _32842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_946 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21922_ _34801_/Q _34737_/Q _34673_/Q _34609_/Q _21888_/X _21889_/X VGND VGND VPWR
+ VPWR _21922_/X sky130_fd_sc_hd__mux4_1
X_33908_ _34228_/CLK _33908_/D VGND VGND VPWR VPWR _33908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25690_ _33271_/Q _24373_/X _25706_/S VGND VGND VPWR VPWR _25691_/A sky130_fd_sc_hd__mux2_1
X_34888_ _35080_/CLK _34888_/D VGND VGND VPWR VPWR _34888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24641_ _24641_/A VGND VGND VPWR VPWR _32809_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33839_ _35760_/CLK _33839_/D VGND VGND VPWR VPWR _33839_/Q sky130_fd_sc_hd__dfxtp_1
X_21853_ _33199_/Q _32559_/Q _35951_/Q _35887_/Q _21674_/X _21675_/X VGND VGND VPWR
+ VPWR _21853_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20804_ _20804_/A _20804_/B _20804_/C _20804_/D VGND VGND VPWR VPWR _20805_/A sky130_fd_sc_hd__or4_2
X_27360_ _34030_/Q _24345_/X _27374_/S VGND VGND VPWR VPWR _27361_/A sky130_fd_sc_hd__mux2_1
X_24572_ _24572_/A VGND VGND VPWR VPWR _32778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21784_ _21599_/X _21782_/X _21783_/X _21602_/X VGND VGND VPWR VPWR _21784_/X sky130_fd_sc_hd__a22o_1
XFILLER_224_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26311_ _26311_/A VGND VGND VPWR VPWR _33564_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23523_ _23523_/A VGND VGND VPWR VPWR _32315_/D sky130_fd_sc_hd__clkbuf_1
X_35509_ _35958_/CLK _35509_/D VGND VGND VPWR VPWR _35509_/Q sky130_fd_sc_hd__dfxtp_1
X_27291_ _27833_/A _30600_/B VGND VGND VPWR VPWR _27424_/S sky130_fd_sc_hd__nor2_8
XFILLER_168_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20735_ _20735_/A VGND VGND VPWR VPWR _36175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29030_ _34821_/Q _24416_/X _29038_/S VGND VGND VPWR VPWR _29031_/A sky130_fd_sc_hd__mux2_1
X_26242_ _25134_/X _33532_/Q _26248_/S VGND VGND VPWR VPWR _26243_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23454_ _23454_/A VGND VGND VPWR VPWR _32282_/D sky130_fd_sc_hd__clkbuf_1
X_20666_ _33166_/Q _32526_/Q _35918_/Q _35854_/Q _20663_/X _20665_/X VGND VGND VPWR
+ VPWR _20666_/X sky130_fd_sc_hd__mux4_1
XFILLER_167_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22405_ _22361_/X _22403_/X _22404_/X _22367_/X VGND VGND VPWR VPWR _22405_/X sky130_fd_sc_hd__a22o_1
XFILLER_17_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26173_ _25032_/X _33499_/Q _26185_/S VGND VGND VPWR VPWR _26174_/A sky130_fd_sc_hd__mux2_1
X_20597_ _22460_/A VGND VGND VPWR VPWR _20597_/X sky130_fd_sc_hd__buf_4
X_23385_ _23385_/A VGND VGND VPWR VPWR _32251_/D sky130_fd_sc_hd__clkbuf_1
X_25124_ _25124_/A VGND VGND VPWR VPWR _33016_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22336_ _22016_/X _22334_/X _22335_/X _22020_/X VGND VGND VPWR VPWR _22336_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_1187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29932_ _35217_/Q _29061_/X _29944_/S VGND VGND VPWR VPWR _29933_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25055_ _25053_/X _32994_/Q _25082_/S VGND VGND VPWR VPWR _25056_/A sky130_fd_sc_hd__mux2_1
X_22267_ _22396_/A VGND VGND VPWR VPWR _22267_/X sky130_fd_sc_hd__buf_4
X_24006_ _22926_/X _32541_/Q _24014_/S VGND VGND VPWR VPWR _24007_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21218_ _21043_/X _21216_/X _21217_/X _21046_/X VGND VGND VPWR VPWR _21218_/X sky130_fd_sc_hd__a22o_1
X_22198_ _22016_/X _22196_/X _22197_/X _22020_/X VGND VGND VPWR VPWR _22198_/X sky130_fd_sc_hd__a22o_1
X_29863_ _29863_/A VGND VGND VPWR VPWR _35184_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28814_ _28814_/A VGND VGND VPWR VPWR _34718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21149_ _21143_/X _21148_/X _21041_/X VGND VGND VPWR VPWR _21157_/C sky130_fd_sc_hd__o21ba_2
X_29794_ _29794_/A VGND VGND VPWR VPWR _35151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28745_ _26971_/X _34686_/Q _28747_/S VGND VGND VPWR VPWR _28746_/A sky130_fd_sc_hd__mux2_1
X_25957_ _25112_/X _33397_/Q _25957_/S VGND VGND VPWR VPWR _25958_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_274_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _34044_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_46_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24908_ _22957_/X _32935_/Q _24916_/S VGND VGND VPWR VPWR _24909_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16690_ _35039_/Q _34975_/Q _34911_/Q _34847_/Q _16450_/X _16451_/X VGND VGND VPWR
+ VPWR _16690_/X sky130_fd_sc_hd__mux4_1
X_28676_ _26869_/X _34653_/Q _28684_/S VGND VGND VPWR VPWR _28677_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25888_ _25010_/X _33364_/Q _25894_/S VGND VGND VPWR VPWR _25889_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24839_ _24839_/A VGND VGND VPWR VPWR _32902_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_30_0_CLK clkbuf_2_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_30_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_34_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27627_ _27696_/S VGND VGND VPWR VPWR _27646_/S sky130_fd_sc_hd__buf_6
XFILLER_46_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _20147_/A VGND VGND VPWR VPWR _18360_/X sky130_fd_sc_hd__buf_6
XFILLER_215_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27558_ _27558_/A VGND VGND VPWR VPWR _34124_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _17063_/X _17309_/X _17310_/X _17067_/X VGND VGND VPWR VPWR _17311_/X sky130_fd_sc_hd__a22o_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26509_ _26509_/A VGND VGND VPWR VPWR _33658_/D sky130_fd_sc_hd__clkbuf_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18291_ _20096_/A VGND VGND VPWR VPWR _18291_/X sky130_fd_sc_hd__buf_4
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27489_ _27489_/A VGND VGND VPWR VPWR _34091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_226_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17055_/X _17240_/X _17241_/X _17061_/X VGND VGND VPWR VPWR _17242_/X sky130_fd_sc_hd__a22o_1
X_29228_ input53/X VGND VGND VPWR VPWR _29228_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29159_ _29159_/A VGND VGND VPWR VPWR _34864_/D sky130_fd_sc_hd__clkbuf_1
X_17173_ _33261_/Q _36141_/Q _33133_/Q _33069_/Q _17058_/X _17059_/X VGND VGND VPWR
+ VPWR _17173_/X sky130_fd_sc_hd__mux4_1
X_16124_ _33167_/Q _32527_/Q _35919_/Q _35855_/Q _16063_/X _16065_/X VGND VGND VPWR
+ VPWR _16124_/X sky130_fd_sc_hd__mux4_1
X_32170_ _35671_/CLK _32170_/D VGND VGND VPWR VPWR _32170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31121_ _31121_/A VGND VGND VPWR VPWR _35780_/D sky130_fd_sc_hd__clkbuf_1
X_16055_ _16044_/X _16047_/X _16052_/X _16054_/X VGND VGND VPWR VPWR _16055_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31052_ _31052_/A VGND VGND VPWR VPWR _35747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30003_ _35251_/Q _29166_/X _30007_/S VGND VGND VPWR VPWR _30004_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19814_ _20167_/A VGND VGND VPWR VPWR _19814_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35860_ _36117_/CLK _35860_/D VGND VGND VPWR VPWR _35860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34811_ _34811_/CLK _34811_/D VGND VGND VPWR VPWR _34811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19745_ _19495_/X _19741_/X _19744_/X _19500_/X VGND VGND VPWR VPWR _19745_/X sky130_fd_sc_hd__a22o_1
X_35791_ _35791_/CLK _35791_/D VGND VGND VPWR VPWR _35791_/Q sky130_fd_sc_hd__dfxtp_1
X_16957_ _32999_/Q _32935_/Q _32871_/Q _32807_/Q _16636_/X _16637_/X VGND VGND VPWR
+ VPWR _16957_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_265_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _34046_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34742_ _34745_/CLK _34742_/D VGND VGND VPWR VPWR _34742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31954_ _34973_/CLK _31954_/D VGND VGND VPWR VPWR _31954_/Q sky130_fd_sc_hd__dfxtp_1
X_19676_ _19502_/X _19672_/X _19675_/X _19505_/X VGND VGND VPWR VPWR _19676_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16888_ _33253_/Q _36133_/Q _33125_/Q _33061_/Q _16705_/X _16706_/X VGND VGND VPWR
+ VPWR _16888_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18627_ _35733_/Q _35093_/Q _34453_/Q _33813_/Q _18349_/X _18351_/X VGND VGND VPWR
+ VPWR _18627_/X sky130_fd_sc_hd__mux4_1
X_30905_ _35678_/Q _29101_/X _30911_/S VGND VGND VPWR VPWR _30906_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34673_ _34932_/CLK _34673_/D VGND VGND VPWR VPWR _34673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31885_ _31885_/A VGND VGND VPWR VPWR _36142_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33624_ _35284_/CLK _33624_/D VGND VGND VPWR VPWR _33624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18558_ _18344_/X _18556_/X _18557_/X _18354_/X VGND VGND VPWR VPWR _18558_/X sky130_fd_sc_hd__a22o_1
X_30836_ _30836_/A VGND VGND VPWR VPWR _35645_/D sky130_fd_sc_hd__clkbuf_1
X_17509_ _17862_/A VGND VGND VPWR VPWR _17509_/X sky130_fd_sc_hd__buf_4
XFILLER_33_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33555_ _33685_/CLK _33555_/D VGND VGND VPWR VPWR _33555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18489_ _35729_/Q _35089_/Q _34449_/Q _33809_/Q _18349_/X _18351_/X VGND VGND VPWR
+ VPWR _18489_/X sky130_fd_sc_hd__mux4_1
X_30767_ _30767_/A VGND VGND VPWR VPWR _35612_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_13 _32115_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20520_ _18326_/X _20518_/X _20519_/X _18337_/X VGND VGND VPWR VPWR _20520_/X sky130_fd_sc_hd__a22o_1
X_32506_ _36027_/CLK _32506_/D VGND VGND VPWR VPWR _32506_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_24 _32116_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33486_ _33490_/CLK _33486_/D VGND VGND VPWR VPWR _33486_/Q sky130_fd_sc_hd__dfxtp_1
X_30698_ _35580_/Q _29194_/X _30704_/S VGND VGND VPWR VPWR _30699_/A sky130_fd_sc_hd__mux2_1
XANTENNA_35 _32117_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 _32119_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 _32126_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20451_ _20160_/X _20449_/X _20450_/X _20165_/X VGND VGND VPWR VPWR _20451_/X sky130_fd_sc_hd__a22o_1
XFILLER_140_1332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35225_ _36201_/CLK _35225_/D VGND VGND VPWR VPWR _35225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_19__f_CLK clkbuf_5_9_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_80_CLK/A sky130_fd_sc_hd__clkbuf_16
XANTENNA_68 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32437_ _34805_/CLK _32437_/D VGND VGND VPWR VPWR _32437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_79 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20382_ _35591_/Q _35527_/Q _35463_/Q _35399_/Q _20256_/X _20257_/X VGND VGND VPWR
+ VPWR _20382_/X sky130_fd_sc_hd__mux4_1
X_23170_ _23170_/A VGND VGND VPWR VPWR _32168_/D sky130_fd_sc_hd__clkbuf_1
X_35156_ _36191_/CLK _35156_/D VGND VGND VPWR VPWR _35156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32368_ _36077_/CLK _32368_/D VGND VGND VPWR VPWR _32368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34107_ _36154_/CLK _34107_/D VGND VGND VPWR VPWR _34107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22121_ _33527_/Q _33463_/Q _33399_/Q _33335_/Q _22076_/X _22077_/X VGND VGND VPWR
+ VPWR _22121_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31319_ _35874_/Q input13/X _31337_/S VGND VGND VPWR VPWR _31320_/A sky130_fd_sc_hd__mux2_1
X_35087_ _35279_/CLK _35087_/D VGND VGND VPWR VPWR _35087_/Q sky130_fd_sc_hd__dfxtp_1
X_32299_ _35179_/CLK _32299_/D VGND VGND VPWR VPWR _32299_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput120 _31987_/Q VGND VGND VPWR VPWR D1[37] sky130_fd_sc_hd__buf_2
Xoutput131 _31997_/Q VGND VGND VPWR VPWR D1[47] sky130_fd_sc_hd__buf_2
Xoutput142 _32007_/Q VGND VGND VPWR VPWR D1[57] sky130_fd_sc_hd__buf_2
XTAP_6508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22052_ _22008_/X _22050_/X _22051_/X _22014_/X VGND VGND VPWR VPWR _22052_/X sky130_fd_sc_hd__a22o_1
XTAP_6519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput153 _31959_/Q VGND VGND VPWR VPWR D1[9] sky130_fd_sc_hd__buf_2
XFILLER_88_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34038_ _34039_/CLK _34038_/D VGND VGND VPWR VPWR _34038_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput164 _36193_/Q VGND VGND VPWR VPWR D2[19] sky130_fd_sc_hd__buf_2
XFILLER_102_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput175 _36203_/Q VGND VGND VPWR VPWR D2[29] sky130_fd_sc_hd__buf_2
Xoutput186 _36213_/Q VGND VGND VPWR VPWR D2[39] sky130_fd_sc_hd__buf_2
Xoutput197 _36223_/Q VGND VGND VPWR VPWR D2[49] sky130_fd_sc_hd__buf_2
XTAP_5807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21003_ _20893_/X _21001_/X _21002_/X _20896_/X VGND VGND VPWR VPWR _21003_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26860_ input4/X VGND VGND VPWR VPWR _26860_/X sky130_fd_sc_hd__buf_4
XFILLER_102_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25811_ _25811_/A VGND VGND VPWR VPWR _33327_/D sky130_fd_sc_hd__clkbuf_1
X_26791_ _26791_/A VGND VGND VPWR VPWR _33791_/D sky130_fd_sc_hd__clkbuf_1
X_35989_ _35989_/CLK _35989_/D VGND VGND VPWR VPWR _35989_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_256_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _36166_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28530_ _28641_/S VGND VGND VPWR VPWR _28549_/S sky130_fd_sc_hd__buf_4
X_25742_ _25742_/A VGND VGND VPWR VPWR _33294_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22954_ input17/X VGND VGND VPWR VPWR _22954_/X sky130_fd_sc_hd__buf_2
XFILLER_112_1467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28461_ _26950_/X _34551_/Q _28477_/S VGND VGND VPWR VPWR _28462_/A sky130_fd_sc_hd__mux2_1
X_21905_ _21901_/X _21904_/X _21728_/X VGND VGND VPWR VPWR _21929_/A sky130_fd_sc_hd__o21ba_1
X_25673_ _33263_/Q _24348_/X _25685_/S VGND VGND VPWR VPWR _25674_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22885_ _22885_/A VGND VGND VPWR VPWR _32015_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27412_ _34055_/Q _24422_/X _27416_/S VGND VGND VPWR VPWR _27413_/A sky130_fd_sc_hd__mux2_1
X_24624_ _24624_/A VGND VGND VPWR VPWR _32801_/D sky130_fd_sc_hd__clkbuf_1
X_28392_ _28392_/A VGND VGND VPWR VPWR _34518_/D sky130_fd_sc_hd__clkbuf_1
X_21836_ _33519_/Q _33455_/Q _33391_/Q _33327_/Q _21723_/X _21724_/X VGND VGND VPWR
+ VPWR _21836_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_1240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27343_ _34022_/Q _24320_/X _27353_/S VGND VGND VPWR VPWR _27344_/A sky130_fd_sc_hd__mux2_1
X_24555_ _23041_/X _32770_/Q _24569_/S VGND VGND VPWR VPWR _24556_/A sky130_fd_sc_hd__mux2_1
X_21767_ _21442_/X _21765_/X _21766_/X _21447_/X VGND VGND VPWR VPWR _21767_/X sky130_fd_sc_hd__a22o_1
XFILLER_51_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23506_ _23506_/A VGND VGND VPWR VPWR _32307_/D sky130_fd_sc_hd__clkbuf_1
X_27274_ _27274_/A VGND VGND VPWR VPWR _33989_/D sky130_fd_sc_hd__clkbuf_1
X_20718_ _20626_/X _20716_/X _20717_/X _20637_/X VGND VGND VPWR VPWR _20718_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24486_ _24486_/A VGND VGND VPWR VPWR _32737_/D sky130_fd_sc_hd__clkbuf_1
X_21698_ _33259_/Q _36139_/Q _33131_/Q _33067_/Q _21658_/X _21659_/X VGND VGND VPWR
+ VPWR _21698_/X sky130_fd_sc_hd__mux4_1
X_29013_ _34813_/Q _24391_/X _29017_/S VGND VGND VPWR VPWR _29014_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26225_ _25109_/X _33524_/Q _26227_/S VGND VGND VPWR VPWR _26226_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23437_ _23437_/A VGND VGND VPWR VPWR _32274_/D sky130_fd_sc_hd__clkbuf_1
X_20649_ _22594_/A VGND VGND VPWR VPWR _20649_/X sky130_fd_sc_hd__buf_6
XFILLER_109_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26156_ _25007_/X _33491_/Q _26164_/S VGND VGND VPWR VPWR _26157_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23368_ _23368_/A VGND VGND VPWR VPWR _32243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25107_ _25106_/X _33011_/Q _25113_/S VGND VGND VPWR VPWR _25108_/A sky130_fd_sc_hd__mux2_1
X_22319_ _22315_/X _22318_/X _22114_/X VGND VGND VPWR VPWR _22320_/D sky130_fd_sc_hd__o21ba_1
X_26087_ _26087_/A VGND VGND VPWR VPWR _33458_/D sky130_fd_sc_hd__clkbuf_1
X_23299_ _23299_/A VGND VGND VPWR VPWR _32217_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29915_ _29915_/A VGND VGND VPWR VPWR _35209_/D sky130_fd_sc_hd__clkbuf_1
X_25038_ input7/X VGND VGND VPWR VPWR _25038_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_117_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_495_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _35038_/CLK sky130_fd_sc_hd__clkbuf_16
X_17860_ _17860_/A VGND VGND VPWR VPWR _17860_/X sky130_fd_sc_hd__buf_4
X_29846_ _29846_/A VGND VGND VPWR VPWR _35176_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16811_ _16811_/A VGND VGND VPWR VPWR _31970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29777_ _35144_/Q _29231_/X _29779_/S VGND VGND VPWR VPWR _29778_/A sky130_fd_sc_hd__mux2_1
X_17791_ _17787_/X _17790_/X _17514_/X VGND VGND VPWR VPWR _17792_/D sky130_fd_sc_hd__o21ba_1
XFILLER_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26989_ _26989_/A VGND VGND VPWR VPWR _33859_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_247_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _33544_/CLK sky130_fd_sc_hd__clkbuf_16
X_19530_ _19524_/X _19529_/X _19461_/X VGND VGND VPWR VPWR _19531_/D sky130_fd_sc_hd__o21ba_1
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28728_ _28776_/S VGND VGND VPWR VPWR _28747_/S sky130_fd_sc_hd__buf_4
X_16742_ _16496_/X _16740_/X _16741_/X _16499_/X VGND VGND VPWR VPWR _16742_/X sky130_fd_sc_hd__a22o_1
XFILLER_247_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19461_ _20167_/A VGND VGND VPWR VPWR _19461_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_62_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16673_ _33247_/Q _36127_/Q _33119_/Q _33055_/Q _16352_/X _16353_/X VGND VGND VPWR
+ VPWR _16673_/X sky130_fd_sc_hd__mux4_1
X_28659_ _26844_/X _34645_/Q _28663_/S VGND VGND VPWR VPWR _28660_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18412_ _18406_/X _18411_/X _18311_/X VGND VGND VPWR VPWR _18434_/A sky130_fd_sc_hd__o21ba_1
XFILLER_59_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31670_ _36041_/Q input55/X _31670_/S VGND VGND VPWR VPWR _31671_/A sky130_fd_sc_hd__mux2_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ _19142_/X _19388_/X _19391_/X _19147_/X VGND VGND VPWR VPWR _19392_/X sky130_fd_sc_hd__a22o_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18343_ _18324_/X _18338_/X _18340_/X _18342_/X VGND VGND VPWR VPWR _18402_/B sky130_fd_sc_hd__o211a_1
X_30621_ _30621_/A VGND VGND VPWR VPWR _35543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33340_ _34044_/CLK _33340_/D VGND VGND VPWR VPWR _33340_/Q sky130_fd_sc_hd__dfxtp_1
X_18274_ _18274_/A VGND VGND VPWR VPWR _32013_/D sky130_fd_sc_hd__clkbuf_1
X_30552_ _30552_/A VGND VGND VPWR VPWR _35510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17225_ _17931_/A VGND VGND VPWR VPWR _17225_/X sky130_fd_sc_hd__buf_6
X_30483_ _23111_/X _35478_/Q _30485_/S VGND VGND VPWR VPWR _30484_/A sky130_fd_sc_hd__mux2_1
Xinput11 DW[19] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__buf_8
X_33271_ _36150_/CLK _33271_/D VGND VGND VPWR VPWR _33271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput22 DW[29] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__buf_4
X_35010_ _35075_/CLK _35010_/D VGND VGND VPWR VPWR _35010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput33 DW[39] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__buf_4
X_32222_ _35843_/CLK _32222_/D VGND VGND VPWR VPWR _32222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput44 DW[49] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__buf_6
X_17156_ _17862_/A VGND VGND VPWR VPWR _17156_/X sky130_fd_sc_hd__buf_4
Xinput55 DW[59] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__buf_8
Xinput66 R1[1] VGND VGND VPWR VPWR input66/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput77 R3[0] VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__clkbuf_1
X_16107_ _33487_/Q _33423_/Q _33359_/Q _33295_/Q _15998_/X _15999_/X VGND VGND VPWR
+ VPWR _16107_/X sky130_fd_sc_hd__mux4_2
XFILLER_239_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput88 RW[5] VGND VGND VPWR VPWR input88/X sky130_fd_sc_hd__clkbuf_4
X_32153_ _35284_/CLK _32153_/D VGND VGND VPWR VPWR _32153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17087_ _17087_/A VGND VGND VPWR VPWR _31978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31104_ _31104_/A VGND VGND VPWR VPWR _35772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16038_ _16026_/X _16031_/X _16036_/X _16037_/X VGND VGND VPWR VPWR _16038_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32084_ _35040_/CLK _32084_/D VGND VGND VPWR VPWR _32084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_486_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _35937_/CLK sky130_fd_sc_hd__clkbuf_16
X_35912_ _35977_/CLK _35912_/D VGND VGND VPWR VPWR _35912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31035_ _31035_/A VGND VGND VPWR VPWR _35739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35843_ _35843_/CLK _35843_/D VGND VGND VPWR VPWR _35843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17989_ _17700_/X _17987_/X _17988_/X _17703_/X VGND VGND VPWR VPWR _17989_/X sky130_fd_sc_hd__a22o_1
XFILLER_111_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_238_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _35331_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19728_ _20232_/A VGND VGND VPWR VPWR _19728_/X sky130_fd_sc_hd__buf_4
X_35774_ _35837_/CLK _35774_/D VGND VGND VPWR VPWR _35774_/Q sky130_fd_sc_hd__dfxtp_1
X_32986_ _33244_/CLK _32986_/D VGND VGND VPWR VPWR _32986_/Q sky130_fd_sc_hd__dfxtp_1
X_34725_ _36003_/CLK _34725_/D VGND VGND VPWR VPWR _34725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31937_ _31937_/A VGND VGND VPWR VPWR _36167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19659_ _20012_/A VGND VGND VPWR VPWR _19659_/X sky130_fd_sc_hd__buf_6
XFILLER_20_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22670_ _22508_/X _22668_/X _22669_/X _22511_/X VGND VGND VPWR VPWR _22670_/X sky130_fd_sc_hd__a22o_1
X_34656_ _34782_/CLK _34656_/D VGND VGND VPWR VPWR _34656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31868_ _31868_/A VGND VGND VPWR VPWR _36134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33607_ _34819_/CLK _33607_/D VGND VGND VPWR VPWR _33607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_1421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21621_ _22447_/A VGND VGND VPWR VPWR _21621_/X sky130_fd_sc_hd__buf_6
XFILLER_179_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30819_ _30819_/A VGND VGND VPWR VPWR _35637_/D sky130_fd_sc_hd__clkbuf_1
X_34587_ _36201_/CLK _34587_/D VGND VGND VPWR VPWR _34587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31799_ _36102_/Q input52/X _31805_/S VGND VGND VPWR VPWR _31800_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_410_CLK clkbuf_6_33__f_CLK/X VGND VGND VPWR VPWR _34986_/CLK sky130_fd_sc_hd__clkbuf_16
X_24340_ _32684_/Q _24338_/X _24367_/S VGND VGND VPWR VPWR _24341_/A sky130_fd_sc_hd__mux2_1
X_33538_ _34050_/CLK _33538_/D VGND VGND VPWR VPWR _33538_/Q sky130_fd_sc_hd__dfxtp_1
X_21552_ _21548_/X _21551_/X _21375_/X VGND VGND VPWR VPWR _21576_/A sky130_fd_sc_hd__o21ba_1
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20503_ _33227_/Q _32587_/Q _35979_/Q _35915_/Q _18375_/X _18376_/X VGND VGND VPWR
+ VPWR _20503_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24271_ _32662_/Q _24270_/X _24274_/S VGND VGND VPWR VPWR _24272_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33469_ _33789_/CLK _33469_/D VGND VGND VPWR VPWR _33469_/Q sky130_fd_sc_hd__dfxtp_1
X_21483_ _33509_/Q _33445_/Q _33381_/Q _33317_/Q _21370_/X _21371_/X VGND VGND VPWR
+ VPWR _21483_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26010_ _26142_/S VGND VGND VPWR VPWR _26029_/S sky130_fd_sc_hd__buf_4
XFILLER_20_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35208_ _35334_/CLK _35208_/D VGND VGND VPWR VPWR _35208_/Q sky130_fd_sc_hd__dfxtp_1
X_23222_ _23222_/A VGND VGND VPWR VPWR _32191_/D sky130_fd_sc_hd__clkbuf_1
X_20434_ _19449_/A _20432_/X _20433_/X _19452_/A VGND VGND VPWR VPWR _20434_/X sky130_fd_sc_hd__a22o_1
XFILLER_181_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36188_ _36189_/CLK _36188_/D VGND VGND VPWR VPWR _36188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35139_ _35780_/CLK _35139_/D VGND VGND VPWR VPWR _35139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23153_ _32163_/Q _23152_/X _23350_/S VGND VGND VPWR VPWR _23154_/A sky130_fd_sc_hd__mux2_1
XTAP_7006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20365_ _33799_/Q _33735_/Q _33671_/Q _33607_/Q _20202_/X _20203_/X VGND VGND VPWR
+ VPWR _20365_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22104_ _35318_/Q _35254_/Q _35190_/Q _32310_/Q _21959_/X _21960_/X VGND VGND VPWR
+ VPWR _22104_/X sky130_fd_sc_hd__mux4_1
XTAP_7039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20296_ _34820_/Q _34756_/Q _34692_/Q _34628_/Q _20294_/X _20295_/X VGND VGND VPWR
+ VPWR _20296_/X sky130_fd_sc_hd__mux4_1
XTAP_6305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27961_ _27961_/A VGND VGND VPWR VPWR _34314_/D sky130_fd_sc_hd__clkbuf_1
X_23084_ _31545_/A _26549_/C VGND VGND VPWR VPWR _23085_/A sky130_fd_sc_hd__or2_1
XTAP_6316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29700_ _35107_/Q _29117_/X _29716_/S VGND VGND VPWR VPWR _29701_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_477_CLK clkbuf_6_9__f_CLK/X VGND VGND VPWR VPWR _35298_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_5604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22035_ _34548_/Q _32436_/Q _34420_/Q _34356_/Q _21825_/X _21826_/X VGND VGND VPWR
+ VPWR _22035_/X sky130_fd_sc_hd__mux4_1
X_26912_ input22/X VGND VGND VPWR VPWR _26912_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27892_ _27892_/A VGND VGND VPWR VPWR _34281_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29631_ _29631_/A VGND VGND VPWR VPWR _35074_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26843_ _26843_/A VGND VGND VPWR VPWR _33812_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_229_CLK clkbuf_6_54__f_CLK/X VGND VGND VPWR VPWR _36037_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29562_ _29652_/S VGND VGND VPWR VPWR _29581_/S sky130_fd_sc_hd__buf_4
X_26774_ _33783_/Q _24373_/X _26790_/S VGND VGND VPWR VPWR _26775_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23986_ _23986_/A VGND VGND VPWR VPWR _32531_/D sky130_fd_sc_hd__clkbuf_1
X_28513_ _28513_/A VGND VGND VPWR VPWR _34575_/D sky130_fd_sc_hd__clkbuf_1
X_25725_ _33288_/Q _24425_/X _25727_/S VGND VGND VPWR VPWR _25726_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22937_ _22937_/A VGND VGND VPWR VPWR _32032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29493_ _23307_/X _35009_/Q _29509_/S VGND VGND VPWR VPWR _29494_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28444_ _26925_/X _34543_/Q _28456_/S VGND VGND VPWR VPWR _28445_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25656_ _33255_/Q _24323_/X _25664_/S VGND VGND VPWR VPWR _25657_/A sky130_fd_sc_hd__mux2_1
X_22868_ _20644_/X _22866_/X _22867_/X _20654_/X VGND VGND VPWR VPWR _22868_/X sky130_fd_sc_hd__a22o_1
XFILLER_243_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24607_ _22914_/X _32793_/Q _24623_/S VGND VGND VPWR VPWR _24608_/A sky130_fd_sc_hd__mux2_1
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28375_ _26821_/X _34510_/Q _28393_/S VGND VGND VPWR VPWR _28376_/A sky130_fd_sc_hd__mux2_1
X_21819_ _33198_/Q _32558_/Q _35950_/Q _35886_/Q _21674_/X _21675_/X VGND VGND VPWR
+ VPWR _21819_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_1070 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25587_ _33224_/Q _24425_/X _25589_/S VGND VGND VPWR VPWR _25588_/A sky130_fd_sc_hd__mux2_1
X_22799_ _35851_/Q _32231_/Q _35723_/Q _35659_/Q _20589_/X _20591_/X VGND VGND VPWR
+ VPWR _22799_/X sky130_fd_sc_hd__mux4_1
XPHY_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_401_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _35562_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27326_ _34014_/Q _24295_/X _27332_/S VGND VGND VPWR VPWR _27327_/A sky130_fd_sc_hd__mux2_1
XPHY_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24538_ _23016_/X _32762_/Q _24548_/S VGND VGND VPWR VPWR _24539_/A sky130_fd_sc_hd__mux2_1
XPHY_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27257_ _27257_/A VGND VGND VPWR VPWR _33981_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24469_ _22914_/X _32729_/Q _24485_/S VGND VGND VPWR VPWR _24470_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17010_ _34536_/Q _32424_/Q _34408_/Q _34344_/Q _16872_/X _16873_/X VGND VGND VPWR
+ VPWR _17010_/X sky130_fd_sc_hd__mux4_1
XFILLER_8_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26208_ _26277_/S VGND VGND VPWR VPWR _26227_/S sky130_fd_sc_hd__buf_4
XFILLER_184_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27188_ _27188_/A VGND VGND VPWR VPWR _33948_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26139_ _26139_/A VGND VGND VPWR VPWR _33483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18961_ _18961_/A _18961_/B _18961_/C _18961_/D VGND VGND VPWR VPWR _18962_/A sky130_fd_sc_hd__or4_1
XFILLER_234_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_468_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _35941_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17912_ _17908_/X _17909_/X _17910_/X _17911_/X VGND VGND VPWR VPWR _17912_/X sky130_fd_sc_hd__a22o_1
XFILLER_156_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18892_ _18892_/A VGND VGND VPWR VPWR _32092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17843_ _17843_/A VGND VGND VPWR VPWR _17843_/X sky130_fd_sc_hd__buf_4
X_29829_ _29829_/A VGND VGND VPWR VPWR _35168_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32840_ _36107_/CLK _32840_/D VGND VGND VPWR VPWR _32840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17774_ _17769_/X _17771_/X _17772_/X _17773_/X VGND VGND VPWR VPWR _17774_/X sky130_fd_sc_hd__a22o_1
XFILLER_19_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19513_ _19363_/X _19511_/X _19512_/X _19367_/X VGND VGND VPWR VPWR _19513_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16725_ _16719_/X _16724_/X _16441_/X VGND VGND VPWR VPWR _16733_/C sky130_fd_sc_hd__o21ba_1
X_32771_ _33026_/CLK _32771_/D VGND VGND VPWR VPWR _32771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34510_ _35728_/CLK _34510_/D VGND VGND VPWR VPWR _34510_/Q sky130_fd_sc_hd__dfxtp_1
X_19444_ _35564_/Q _35500_/Q _35436_/Q _35372_/Q _19197_/X _19198_/X VGND VGND VPWR
+ VPWR _19444_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31722_ _31722_/A VGND VGND VPWR VPWR _36065_/D sky130_fd_sc_hd__clkbuf_1
X_35490_ _35940_/CLK _35490_/D VGND VGND VPWR VPWR _35490_/Q sky130_fd_sc_hd__dfxtp_1
X_16656_ _16443_/X _16652_/X _16655_/X _16446_/X VGND VGND VPWR VPWR _16656_/X sky130_fd_sc_hd__a22o_1
XFILLER_16_960 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34441_ _35337_/CLK _34441_/D VGND VGND VPWR VPWR _34441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31653_ _31653_/A VGND VGND VPWR VPWR _36032_/D sky130_fd_sc_hd__clkbuf_1
X_19375_ _20232_/A VGND VGND VPWR VPWR _19375_/X sky130_fd_sc_hd__buf_4
X_16587_ _34524_/Q _32412_/Q _34396_/Q _34332_/Q _16519_/X _16520_/X VGND VGND VPWR
+ VPWR _16587_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30604_ _35535_/Q _29055_/X _30620_/S VGND VGND VPWR VPWR _30605_/A sky130_fd_sc_hd__mux2_1
X_18326_ _20208_/A VGND VGND VPWR VPWR _18326_/X sky130_fd_sc_hd__clkbuf_4
X_34372_ _35332_/CLK _34372_/D VGND VGND VPWR VPWR _34372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31584_ _36000_/Q input10/X _31586_/S VGND VGND VPWR VPWR _31585_/A sky130_fd_sc_hd__mux2_1
X_36111_ _36112_/CLK _36111_/D VGND VGND VPWR VPWR _36111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33323_ _33512_/CLK _33323_/D VGND VGND VPWR VPWR _33323_/Q sky130_fd_sc_hd__dfxtp_1
X_18257_ _17154_/A _18255_/X _18256_/X _17159_/A VGND VGND VPWR VPWR _18257_/X sky130_fd_sc_hd__a22o_1
X_30535_ _30535_/A VGND VGND VPWR VPWR _35502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36042_ _36170_/CLK _36042_/D VGND VGND VPWR VPWR _36042_/Q sky130_fd_sc_hd__dfxtp_1
X_17208_ _32750_/Q _32686_/Q _32622_/Q _36078_/Q _16919_/X _17056_/X VGND VGND VPWR
+ VPWR _17208_/X sky130_fd_sc_hd__mux4_1
X_30466_ _30598_/S VGND VGND VPWR VPWR _30485_/S sky130_fd_sc_hd__buf_4
X_33254_ _36135_/CLK _33254_/D VGND VGND VPWR VPWR _33254_/Q sky130_fd_sc_hd__dfxtp_1
X_18188_ _33547_/Q _33483_/Q _33419_/Q _33355_/Q _16033_/X _16035_/X VGND VGND VPWR
+ VPWR _18188_/X sky130_fd_sc_hd__mux4_2
XFILLER_11_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32205_ _35827_/CLK _32205_/D VGND VGND VPWR VPWR _32205_/Q sky130_fd_sc_hd__dfxtp_1
X_17139_ _35820_/Q _32197_/Q _35692_/Q _35628_/Q _16960_/X _16961_/X VGND VGND VPWR
+ VPWR _17139_/X sky130_fd_sc_hd__mux4_1
X_30397_ _23241_/X _35437_/Q _30413_/S VGND VGND VPWR VPWR _30398_/A sky130_fd_sc_hd__mux2_1
X_33185_ _35938_/CLK _33185_/D VGND VGND VPWR VPWR _33185_/Q sky130_fd_sc_hd__dfxtp_1
X_20150_ _35584_/Q _35520_/Q _35456_/Q _35392_/Q _19903_/X _19904_/X VGND VGND VPWR
+ VPWR _20150_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32136_ _35815_/CLK _32136_/D VGND VGND VPWR VPWR _32136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_459_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _35302_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_48_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20081_ _20232_/A VGND VGND VPWR VPWR _20081_/X sky130_fd_sc_hd__buf_4
XFILLER_170_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32067_ _36034_/CLK _32067_/D VGND VGND VPWR VPWR _32067_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31018_ _31018_/A VGND VGND VPWR VPWR _35731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23840_ _23840_/A VGND VGND VPWR VPWR _32462_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35826_ _35826_/CLK _35826_/D VGND VGND VPWR VPWR _35826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23771_ _23771_/A VGND VGND VPWR VPWR _32430_/D sky130_fd_sc_hd__clkbuf_1
X_35757_ _35757_/CLK _35757_/D VGND VGND VPWR VPWR _35757_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_509 _17900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32969_ _36107_/CLK _32969_/D VGND VGND VPWR VPWR _32969_/Q sky130_fd_sc_hd__dfxtp_1
X_20983_ _22556_/A VGND VGND VPWR VPWR _20983_/X sky130_fd_sc_hd__buf_6
XFILLER_26_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25510_ _33187_/Q _24311_/X _25526_/S VGND VGND VPWR VPWR _25511_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22722_ _22718_/X _22721_/X _22467_/X VGND VGND VPWR VPWR _22723_/D sky130_fd_sc_hd__o21ba_1
X_34708_ _35286_/CLK _34708_/D VGND VGND VPWR VPWR _34708_/Q sky130_fd_sc_hd__dfxtp_1
X_26490_ _26490_/A VGND VGND VPWR VPWR _33649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35688_ _35879_/CLK _35688_/D VGND VGND VPWR VPWR _35688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25441_ _25441_/A VGND VGND VPWR VPWR _33156_/D sky130_fd_sc_hd__clkbuf_1
X_34639_ _35215_/CLK _34639_/D VGND VGND VPWR VPWR _34639_/Q sky130_fd_sc_hd__dfxtp_1
X_22653_ _33222_/Q _32582_/Q _35974_/Q _35910_/Q _22380_/X _22381_/X VGND VGND VPWR
+ VPWR _22653_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21604_ _21598_/X _21603_/X _21394_/X VGND VGND VPWR VPWR _21614_/C sky130_fd_sc_hd__o21ba_1
X_28160_ _28160_/A VGND VGND VPWR VPWR _34408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25372_ _25372_/A VGND VGND VPWR VPWR _33123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22584_ _33028_/Q _32964_/Q _32900_/Q _32836_/Q _22295_/X _22296_/X VGND VGND VPWR
+ VPWR _22584_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27111_ _26953_/X _33912_/Q _27125_/S VGND VGND VPWR VPWR _27112_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24323_ input18/X VGND VGND VPWR VPWR _24323_/X sky130_fd_sc_hd__clkbuf_4
X_28091_ _27002_/X _34376_/Q _28093_/S VGND VGND VPWR VPWR _28092_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21535_ _22594_/A VGND VGND VPWR VPWR _21535_/X sky130_fd_sc_hd__buf_6
XFILLER_194_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27042_ _27042_/A VGND VGND VPWR VPWR _33879_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24254_ _24254_/A VGND VGND VPWR VPWR _32656_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21466_ _33188_/Q _32548_/Q _35940_/Q _35876_/Q _21321_/X _21322_/X VGND VGND VPWR
+ VPWR _21466_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1090 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23205_ _23205_/A VGND VGND VPWR VPWR _32184_/D sky130_fd_sc_hd__clkbuf_1
X_20417_ _35336_/Q _35272_/Q _35208_/Q _32328_/Q _18388_/X _18390_/X VGND VGND VPWR
+ VPWR _20417_/X sky130_fd_sc_hd__mux4_1
XFILLER_134_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24185_ _24185_/A VGND VGND VPWR VPWR _32625_/D sky130_fd_sc_hd__clkbuf_1
X_21397_ _34786_/Q _34722_/Q _34658_/Q _34594_/Q _21182_/X _21183_/X VGND VGND VPWR
+ VPWR _21397_/X sky130_fd_sc_hd__mux4_1
XFILLER_218_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23136_ input8/X VGND VGND VPWR VPWR _23136_/X sky130_fd_sc_hd__buf_4
XFILLER_107_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20348_ _20344_/X _20347_/X _20142_/X _20143_/X VGND VGND VPWR VPWR _20363_/B sky130_fd_sc_hd__o211a_1
XTAP_6102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28993_ _28993_/A VGND VGND VPWR VPWR _34803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_930 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27944_ _34306_/Q _24407_/X _27958_/S VGND VGND VPWR VPWR _27945_/A sky130_fd_sc_hd__mux2_1
XTAP_6135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23067_ _23067_/A VGND VGND VPWR VPWR _32074_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20279_ _32772_/Q _32708_/Q _32644_/Q _36100_/Q _20278_/X _20062_/X VGND VGND VPWR
+ VPWR _20279_/X sky130_fd_sc_hd__mux4_1
XTAP_5401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22018_ _32500_/Q _32372_/Q _32052_/Q _36020_/Q _21876_/X _22017_/X VGND VGND VPWR
+ VPWR _22018_/X sky130_fd_sc_hd__mux4_1
XFILLER_216_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27875_ _27875_/A VGND VGND VPWR VPWR _34273_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29614_ _29614_/A VGND VGND VPWR VPWR _35066_/D sky130_fd_sc_hd__clkbuf_1
X_26826_ input12/X VGND VGND VPWR VPWR _26826_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29545_ _29545_/A VGND VGND VPWR VPWR _35033_/D sky130_fd_sc_hd__clkbuf_1
X_23969_ _23969_/A VGND VGND VPWR VPWR _32524_/D sky130_fd_sc_hd__clkbuf_1
X_26757_ _33775_/Q _24348_/X _26769_/S VGND VGND VPWR VPWR _26758_/A sky130_fd_sc_hd__mux2_1
XTAP_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16510_ _35738_/Q _35098_/Q _34458_/Q _33818_/Q _16434_/X _16435_/X VGND VGND VPWR
+ VPWR _16510_/X sky130_fd_sc_hd__mux4_1
XFILLER_205_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25708_ _25735_/S VGND VGND VPWR VPWR _25727_/S sky130_fd_sc_hd__buf_6
XFILLER_229_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26688_ _33742_/Q _24244_/X _26706_/S VGND VGND VPWR VPWR _26689_/A sky130_fd_sc_hd__mux2_1
X_17490_ _17843_/A VGND VGND VPWR VPWR _17490_/X sky130_fd_sc_hd__clkbuf_4
X_29476_ _23280_/X _35001_/Q _29488_/S VGND VGND VPWR VPWR _29477_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_1479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16441_ _17853_/A VGND VGND VPWR VPWR _16441_/X sky130_fd_sc_hd__buf_2
X_28427_ _26900_/X _34535_/Q _28435_/S VGND VGND VPWR VPWR _28428_/A sky130_fd_sc_hd__mux2_1
X_25639_ _33247_/Q _24298_/X _25643_/S VGND VGND VPWR VPWR _25640_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16372_ _16366_/X _16371_/X _16071_/X VGND VGND VPWR VPWR _16380_/C sky130_fd_sc_hd__o21ba_1
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19160_ _19010_/X _19158_/X _19159_/X _19014_/X VGND VGND VPWR VPWR _19160_/X sky130_fd_sc_hd__a22o_1
X_28358_ _28358_/A VGND VGND VPWR VPWR _34502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18111_ _15977_/X _18109_/X _18110_/X _15987_/X VGND VGND VPWR VPWR _18111_/X sky130_fd_sc_hd__a22o_1
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27309_ _34006_/Q _24270_/X _27311_/S VGND VGND VPWR VPWR _27310_/A sky130_fd_sc_hd__mux2_1
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19091_ _35554_/Q _35490_/Q _35426_/Q _35362_/Q _18844_/X _18845_/X VGND VGND VPWR
+ VPWR _19091_/X sky130_fd_sc_hd__mux4_1
X_28289_ _28289_/A VGND VGND VPWR VPWR _34469_/D sky130_fd_sc_hd__clkbuf_1
X_30320_ _30320_/A VGND VGND VPWR VPWR _35401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18042_ _32774_/Q _32710_/Q _32646_/Q _36102_/Q _17978_/X _17762_/X VGND VGND VPWR
+ VPWR _18042_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30251_ _30251_/A VGND VGND VPWR VPWR _35368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30182_ _35336_/Q _29231_/X _30184_/S VGND VGND VPWR VPWR _30183_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19993_ _19708_/X _19991_/X _19992_/X _19714_/X VGND VGND VPWR VPWR _19993_/X sky130_fd_sc_hd__a22o_1
XFILLER_154_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18944_ _20158_/A VGND VGND VPWR VPWR _18944_/X sky130_fd_sc_hd__clkbuf_4
X_34990_ _35054_/CLK _34990_/D VGND VGND VPWR VPWR _34990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33941_ _34001_/CLK _33941_/D VGND VGND VPWR VPWR _33941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18875_ _35804_/Q _32179_/Q _35676_/Q _35612_/Q _18554_/X _18555_/X VGND VGND VPWR
+ VPWR _18875_/X sky130_fd_sc_hd__mux4_1
XTAP_6680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17826_ _33792_/Q _33728_/Q _33664_/Q _33600_/Q _17549_/X _17550_/X VGND VGND VPWR
+ VPWR _17826_/X sky130_fd_sc_hd__mux4_1
X_33872_ _34001_/CLK _33872_/D VGND VGND VPWR VPWR _33872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35611_ _35803_/CLK _35611_/D VGND VGND VPWR VPWR _35611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32823_ _36024_/CLK _32823_/D VGND VGND VPWR VPWR _32823_/Q sky130_fd_sc_hd__dfxtp_1
X_17757_ _33534_/Q _33470_/Q _33406_/Q _33342_/Q _17476_/X _17477_/X VGND VGND VPWR
+ VPWR _17757_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35542_ _35927_/CLK _35542_/D VGND VGND VPWR VPWR _35542_/Q sky130_fd_sc_hd__dfxtp_1
X_16708_ _17906_/A VGND VGND VPWR VPWR _16708_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_35_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32754_ _36141_/CLK _32754_/D VGND VGND VPWR VPWR _32754_/Q sky130_fd_sc_hd__dfxtp_1
X_17688_ _34044_/Q _33980_/Q _33916_/Q _32252_/Q _17373_/X _17374_/X VGND VGND VPWR
+ VPWR _17688_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31705_ _36057_/Q input3/X _31721_/S VGND VGND VPWR VPWR _31706_/A sky130_fd_sc_hd__mux2_1
X_19427_ _19149_/X _19425_/X _19426_/X _19152_/X VGND VGND VPWR VPWR _19427_/X sky130_fd_sc_hd__a22o_1
X_35473_ _35921_/CLK _35473_/D VGND VGND VPWR VPWR _35473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16639_ _16357_/X _16635_/X _16638_/X _16361_/X VGND VGND VPWR VPWR _16639_/X sky130_fd_sc_hd__a22o_1
X_32685_ _36076_/CLK _32685_/D VGND VGND VPWR VPWR _32685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34424_ _35319_/CLK _34424_/D VGND VGND VPWR VPWR _34424_/Q sky130_fd_sc_hd__dfxtp_1
X_31636_ _31636_/A VGND VGND VPWR VPWR _36024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19358_ _20282_/A VGND VGND VPWR VPWR _19358_/X sky130_fd_sc_hd__buf_6
XFILLER_241_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18309_ _18297_/X _18300_/X _18303_/X _18308_/X VGND VGND VPWR VPWR _18309_/X sky130_fd_sc_hd__a22o_1
XFILLER_200_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34355_ _34805_/CLK _34355_/D VGND VGND VPWR VPWR _34355_/Q sky130_fd_sc_hd__dfxtp_1
X_19289_ _20129_/A VGND VGND VPWR VPWR _19289_/X sky130_fd_sc_hd__buf_6
X_31567_ _31678_/S VGND VGND VPWR VPWR _31586_/S sky130_fd_sc_hd__buf_4
X_33306_ _34202_/CLK _33306_/D VGND VGND VPWR VPWR _33306_/Q sky130_fd_sc_hd__dfxtp_1
X_21320_ _35552_/Q _35488_/Q _35424_/Q _35360_/Q _21144_/X _21145_/X VGND VGND VPWR
+ VPWR _21320_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30518_ _30518_/A VGND VGND VPWR VPWR _35494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34286_ _34286_/CLK _34286_/D VGND VGND VPWR VPWR _34286_/Q sky130_fd_sc_hd__dfxtp_1
X_31498_ _23274_/X _35959_/Q _31514_/S VGND VGND VPWR VPWR _31499_/A sky130_fd_sc_hd__mux2_1
X_36025_ _36025_/CLK _36025_/D VGND VGND VPWR VPWR _36025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33237_ _36117_/CLK _33237_/D VGND VGND VPWR VPWR _33237_/Q sky130_fd_sc_hd__dfxtp_1
X_21251_ _21245_/X _21250_/X _21041_/X VGND VGND VPWR VPWR _21261_/C sky130_fd_sc_hd__o21ba_2
XFILLER_50_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30449_ _23322_/X _35462_/Q _30455_/S VGND VGND VPWR VPWR _30450_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_1331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20202_ _20202_/A VGND VGND VPWR VPWR _20202_/X sky130_fd_sc_hd__buf_6
XFILLER_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33168_ _34317_/CLK _33168_/D VGND VGND VPWR VPWR _33168_/Q sky130_fd_sc_hd__dfxtp_1
X_21182_ _22594_/A VGND VGND VPWR VPWR _21182_/X sky130_fd_sc_hd__buf_6
XFILLER_145_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20133_ _19855_/X _20131_/X _20132_/X _19858_/X VGND VGND VPWR VPWR _20133_/X sky130_fd_sc_hd__a22o_1
X_32119_ _35811_/CLK _32119_/D VGND VGND VPWR VPWR _32119_/Q sky130_fd_sc_hd__dfxtp_1
X_25990_ _25990_/A VGND VGND VPWR VPWR _33412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33099_ _33548_/CLK _33099_/D VGND VGND VPWR VPWR _33099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20064_ _20282_/A VGND VGND VPWR VPWR _20064_/X sky130_fd_sc_hd__buf_4
X_24941_ _24941_/A VGND VGND VPWR VPWR _32950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27660_ _27660_/A VGND VGND VPWR VPWR _34171_/D sky130_fd_sc_hd__clkbuf_1
X_24872_ _22904_/X _32918_/Q _24874_/S VGND VGND VPWR VPWR _24873_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23823_ _23823_/A VGND VGND VPWR VPWR _32455_/D sky130_fd_sc_hd__clkbuf_1
X_26611_ _26611_/A VGND VGND VPWR VPWR _33706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35809_ _35809_/CLK _35809_/D VGND VGND VPWR VPWR _35809_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27591_ _27591_/A VGND VGND VPWR VPWR _34138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_306 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26542_ _26542_/A VGND VGND VPWR VPWR _33674_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_317 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29330_ _23264_/X _34932_/Q _29332_/S VGND VGND VPWR VPWR _29331_/A sky130_fd_sc_hd__mux2_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_328 _32141_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23754_ _23754_/A VGND VGND VPWR VPWR _32422_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20966_ _20888_/X _20964_/X _20965_/X _20891_/X VGND VGND VPWR VPWR _20966_/X sky130_fd_sc_hd__a22o_1
XANTENNA_339 _36205_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_213_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22705_ _32520_/Q _32392_/Q _32072_/Q _36040_/Q _22582_/X _21607_/A VGND VGND VPWR
+ VPWR _22705_/X sky130_fd_sc_hd__mux4_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29261_ _23102_/X _34899_/Q _29269_/S VGND VGND VPWR VPWR _29262_/A sky130_fd_sc_hd__mux2_1
X_26473_ _26473_/A VGND VGND VPWR VPWR _33641_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23685_ _23685_/A VGND VGND VPWR VPWR _32391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20897_ _20893_/X _20894_/X _20895_/X _20896_/X VGND VGND VPWR VPWR _20897_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28212_ _26981_/X _34433_/Q _28228_/S VGND VGND VPWR VPWR _28213_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25424_ _25424_/A VGND VGND VPWR VPWR _33148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22636_ _34310_/Q _34246_/Q _34182_/Q _34118_/Q _22395_/X _22396_/X VGND VGND VPWR
+ VPWR _22636_/X sky130_fd_sc_hd__mux4_1
X_29192_ _34875_/Q _29191_/X _29204_/S VGND VGND VPWR VPWR _29193_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25355_ _25355_/A VGND VGND VPWR VPWR _33115_/D sky130_fd_sc_hd__clkbuf_1
X_28143_ _28143_/A VGND VGND VPWR VPWR _34400_/D sky130_fd_sc_hd__clkbuf_1
X_22567_ _22460_/X _22565_/X _22566_/X _22465_/X VGND VGND VPWR VPWR _22567_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24306_ _24306_/A VGND VGND VPWR VPWR _32673_/D sky130_fd_sc_hd__clkbuf_1
X_28074_ _28101_/S VGND VGND VPWR VPWR _28093_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_194_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21518_ _21514_/X _21517_/X _21375_/X VGND VGND VPWR VPWR _21544_/A sky130_fd_sc_hd__o21ba_1
X_25286_ _25286_/A VGND VGND VPWR VPWR _33083_/D sky130_fd_sc_hd__clkbuf_1
X_22498_ _22494_/X _22497_/X _22467_/X VGND VGND VPWR VPWR _22499_/D sky130_fd_sc_hd__o21ba_1
XFILLER_182_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27025_ _26826_/X _33871_/Q _27041_/S VGND VGND VPWR VPWR _27026_/A sky130_fd_sc_hd__mux2_1
X_24237_ _24237_/A VGND VGND VPWR VPWR _32650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21449_ _22508_/A VGND VGND VPWR VPWR _21449_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_135_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24168_ _24168_/A VGND VGND VPWR VPWR _32617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23119_ _32152_/Q _23117_/X _23146_/S VGND VGND VPWR VPWR _23120_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24099_ _24099_/A VGND VGND VPWR VPWR _32585_/D sky130_fd_sc_hd__clkbuf_1
X_28976_ _28976_/A VGND VGND VPWR VPWR _34795_/D sky130_fd_sc_hd__clkbuf_1
X_16990_ _17830_/A VGND VGND VPWR VPWR _16990_/X sky130_fd_sc_hd__buf_6
XFILLER_110_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27927_ _34298_/Q _24382_/X _27937_/S VGND VGND VPWR VPWR _27928_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18660_ _32982_/Q _32918_/Q _32854_/Q _32790_/Q _18583_/X _18584_/X VGND VGND VPWR
+ VPWR _18660_/X sky130_fd_sc_hd__mux4_1
XTAP_5275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27858_ _34265_/Q _24280_/X _27874_/S VGND VGND VPWR VPWR _27859_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17611_ _17502_/X _17609_/X _17610_/X _17505_/X VGND VGND VPWR VPWR _17611_/X sky130_fd_sc_hd__a22o_1
X_26809_ _33800_/Q _24425_/X _26811_/S VGND VGND VPWR VPWR _26810_/A sky130_fd_sc_hd__mux2_1
XTAP_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18591_ _20158_/A VGND VGND VPWR VPWR _18591_/X sky130_fd_sc_hd__buf_4
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27789_ _27789_/A VGND VGND VPWR VPWR _34232_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29528_ _29528_/A VGND VGND VPWR VPWR _35025_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ _34551_/Q _32439_/Q _34423_/Q _34359_/Q _17225_/X _17226_/X VGND VGND VPWR
+ VPWR _17542_/X sky130_fd_sc_hd__mux4_1
XFILLER_217_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_840 _23322_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_851 _24401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_862 _24407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29459_ _23253_/X _34993_/Q _29467_/S VGND VGND VPWR VPWR _29460_/A sky130_fd_sc_hd__mux2_1
X_17473_ _33782_/Q _33718_/Q _33654_/Q _33590_/Q _17196_/X _17197_/X VGND VGND VPWR
+ VPWR _17473_/X sky130_fd_sc_hd__mux4_1
XANTENNA_873 _24987_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_884 _25088_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_895 _25735_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19212_ _33766_/Q _33702_/Q _33638_/Q _33574_/Q _19143_/X _19144_/X VGND VGND VPWR
+ VPWR _19212_/X sky130_fd_sc_hd__mux4_1
X_16424_ _32728_/Q _32664_/Q _32600_/Q _36056_/Q _16213_/X _16350_/X VGND VGND VPWR
+ VPWR _16424_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32470_ _33507_/CLK _32470_/D VGND VGND VPWR VPWR _32470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31421_ _31421_/A VGND VGND VPWR VPWR _35922_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19143_ _20202_/A VGND VGND VPWR VPWR _19143_/X sky130_fd_sc_hd__buf_4
X_16355_ _17906_/A VGND VGND VPWR VPWR _16355_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_34_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34140_ _34777_/CLK _34140_/D VGND VGND VPWR VPWR _34140_/Q sky130_fd_sc_hd__dfxtp_1
X_16286_ _16026_/X _16282_/X _16285_/X _16037_/X VGND VGND VPWR VPWR _16286_/X sky130_fd_sc_hd__a22o_1
X_31352_ _35890_/Q input30/X _31358_/S VGND VGND VPWR VPWR _31353_/A sky130_fd_sc_hd__mux2_1
X_19074_ _18796_/X _19072_/X _19073_/X _18799_/X VGND VGND VPWR VPWR _19074_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18025_ _18021_/X _18024_/X _17853_/X VGND VGND VPWR VPWR _18033_/C sky130_fd_sc_hd__o21ba_1
XFILLER_201_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30303_ _35393_/Q _29210_/X _30319_/S VGND VGND VPWR VPWR _30304_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34071_ _35730_/CLK _34071_/D VGND VGND VPWR VPWR _34071_/Q sky130_fd_sc_hd__dfxtp_1
X_31283_ _35857_/Q input34/X _31295_/S VGND VGND VPWR VPWR _31284_/A sky130_fd_sc_hd__mux2_1
X_33022_ _36097_/CLK _33022_/D VGND VGND VPWR VPWR _33022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30234_ _30234_/A VGND VGND VPWR VPWR _35360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30165_ _30192_/S VGND VGND VPWR VPWR _30184_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_99_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19976_ _35323_/Q _35259_/Q _35195_/Q _32315_/Q _19659_/X _19660_/X VGND VGND VPWR
+ VPWR _19976_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18927_ _18789_/X _18925_/X _18926_/X _18794_/X VGND VGND VPWR VPWR _18927_/X sky130_fd_sc_hd__a22o_1
X_30096_ _35295_/Q _29104_/X _30100_/S VGND VGND VPWR VPWR _30097_/A sky130_fd_sc_hd__mux2_1
X_34973_ _34973_/CLK _34973_/D VGND VGND VPWR VPWR _34973_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1250 _26683_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1261 _29046_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1272 _31138_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33924_ _34306_/CLK _33924_/D VGND VGND VPWR VPWR _33924_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1283 _17842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18858_ _18858_/A VGND VGND VPWR VPWR _32091_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_1294 _17853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17809_ _17805_/X _17808_/X _17489_/X _17490_/X VGND VGND VPWR VPWR _17824_/B sky130_fd_sc_hd__o211a_1
XFILLER_83_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33855_ _35903_/CLK _33855_/D VGND VGND VPWR VPWR _33855_/Q sky130_fd_sc_hd__dfxtp_1
X_18789_ _20201_/A VGND VGND VPWR VPWR _18789_/X sky130_fd_sc_hd__buf_4
XFILLER_227_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20820_ _20626_/X _20818_/X _20819_/X _20637_/X VGND VGND VPWR VPWR _20820_/X sky130_fd_sc_hd__a22o_1
X_32806_ _36007_/CLK _32806_/D VGND VGND VPWR VPWR _32806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33786_ _34298_/CLK _33786_/D VGND VGND VPWR VPWR _33786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30998_ _30998_/A VGND VGND VPWR VPWR _35722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35525_ _36168_/CLK _35525_/D VGND VGND VPWR VPWR _35525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20751_ _20614_/X _20749_/X _20750_/X _20623_/X VGND VGND VPWR VPWR _20751_/X sky130_fd_sc_hd__a22o_1
X_32737_ _36065_/CLK _32737_/D VGND VGND VPWR VPWR _32737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35456_ _35585_/CLK _35456_/D VGND VGND VPWR VPWR _35456_/Q sky130_fd_sc_hd__dfxtp_1
X_23470_ _22941_/X _32290_/Q _23488_/S VGND VGND VPWR VPWR _23471_/A sky130_fd_sc_hd__mux2_1
X_20682_ _35278_/Q _35214_/Q _35150_/Q _32270_/Q _20679_/X _20681_/X VGND VGND VPWR
+ VPWR _20682_/X sky130_fd_sc_hd__mux4_1
XFILLER_126_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32668_ _36127_/CLK _32668_/D VGND VGND VPWR VPWR _32668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22421_ _35071_/Q _35007_/Q _34943_/Q _34879_/Q _22109_/X _22110_/X VGND VGND VPWR
+ VPWR _22421_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34407_ _35302_/CLK _34407_/D VGND VGND VPWR VPWR _34407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31619_ _31619_/A VGND VGND VPWR VPWR _36016_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35387_ _35579_/CLK _35387_/D VGND VGND VPWR VPWR _35387_/Q sky130_fd_sc_hd__dfxtp_1
X_32599_ _36055_/CLK _32599_/D VGND VGND VPWR VPWR _32599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25140_ input43/X VGND VGND VPWR VPWR _25140_/X sky130_fd_sc_hd__buf_2
X_22352_ _22352_/A _22352_/B _22352_/C _22352_/D VGND VGND VPWR VPWR _22353_/A sky130_fd_sc_hd__or4_4
XFILLER_143_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34338_ _35932_/CLK _34338_/D VGND VGND VPWR VPWR _34338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21303_ _22362_/A VGND VGND VPWR VPWR _21303_/X sky130_fd_sc_hd__clkbuf_4
X_25071_ _25071_/A VGND VGND VPWR VPWR _32999_/D sky130_fd_sc_hd__clkbuf_1
X_22283_ _22283_/A VGND VGND VPWR VPWR _36219_/D sky130_fd_sc_hd__clkbuf_1
X_34269_ _34779_/CLK _34269_/D VGND VGND VPWR VPWR _34269_/Q sky130_fd_sc_hd__dfxtp_1
X_24022_ _24022_/A VGND VGND VPWR VPWR _32548_/D sky130_fd_sc_hd__clkbuf_1
X_36008_ _36072_/CLK _36008_/D VGND VGND VPWR VPWR _36008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21234_ _20949_/X _21232_/X _21233_/X _20955_/X VGND VGND VPWR VPWR _21234_/X sky130_fd_sc_hd__a22o_1
X_28830_ _26897_/X _34726_/Q _28840_/S VGND VGND VPWR VPWR _28831_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21165_ _21161_/X _21164_/X _21022_/X VGND VGND VPWR VPWR _21191_/A sky130_fd_sc_hd__o21ba_1
XFILLER_236_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20116_ _20112_/X _20115_/X _19800_/X VGND VGND VPWR VPWR _20124_/C sky130_fd_sc_hd__o21ba_1
XFILLER_131_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28761_ _28761_/A VGND VGND VPWR VPWR _34693_/D sky130_fd_sc_hd__clkbuf_1
X_25973_ _25973_/A VGND VGND VPWR VPWR _33404_/D sky130_fd_sc_hd__clkbuf_1
X_21096_ _22508_/A VGND VGND VPWR VPWR _21096_/X sky130_fd_sc_hd__buf_4
XFILLER_219_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27712_ _34196_/Q _24264_/X _27718_/S VGND VGND VPWR VPWR _27713_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20047_ _19802_/X _20045_/X _20046_/X _19805_/X VGND VGND VPWR VPWR _20047_/X sky130_fd_sc_hd__a22o_1
X_24924_ _24924_/A VGND VGND VPWR VPWR _32942_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28692_ _28692_/A VGND VGND VPWR VPWR _34660_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27643_ _27643_/A VGND VGND VPWR VPWR _34163_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24855_ _24987_/S VGND VGND VPWR VPWR _24874_/S sky130_fd_sc_hd__buf_4
XFILLER_73_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_103 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23806_ _23806_/A VGND VGND VPWR VPWR _32447_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_114 _32129_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27574_ _27574_/A VGND VGND VPWR VPWR _34130_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_125 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24786_ _22976_/X _32877_/Q _24802_/S VGND VGND VPWR VPWR _24787_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21998_ _21994_/X _21997_/X _21761_/X VGND VGND VPWR VPWR _21999_/D sky130_fd_sc_hd__o21ba_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_136 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29313_ _29382_/S VGND VGND VPWR VPWR _29332_/S sky130_fd_sc_hd__buf_4
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26525_ _25153_/X _33666_/Q _26539_/S VGND VGND VPWR VPWR _26526_/A sky130_fd_sc_hd__mux2_1
X_23737_ _23737_/A VGND VGND VPWR VPWR _32414_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_158 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20949_ _22501_/A VGND VGND VPWR VPWR _20949_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_169 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29244_ _34892_/Q _29243_/X _29247_/S VGND VGND VPWR VPWR _29245_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23668_ _23668_/A VGND VGND VPWR VPWR _32383_/D sky130_fd_sc_hd__clkbuf_1
X_26456_ _26456_/A VGND VGND VPWR VPWR _33633_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22619_ _35845_/Q _32224_/Q _35717_/Q _35653_/Q _20589_/X _20591_/X VGND VGND VPWR
+ VPWR _22619_/X sky130_fd_sc_hd__mux4_1
X_25407_ _25407_/A VGND VGND VPWR VPWR _33140_/D sky130_fd_sc_hd__clkbuf_1
X_26387_ _26387_/A VGND VGND VPWR VPWR _33600_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29175_ input35/X VGND VGND VPWR VPWR _29175_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_224_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23599_ _23599_/A VGND VGND VPWR VPWR _32350_/D sky130_fd_sc_hd__clkbuf_1
X_16140_ _34256_/Q _34192_/Q _34128_/Q _34064_/Q _16005_/X _16007_/X VGND VGND VPWR
+ VPWR _16140_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25338_ _25338_/A VGND VGND VPWR VPWR _33107_/D sky130_fd_sc_hd__clkbuf_1
X_28126_ _26853_/X _34392_/Q _28144_/S VGND VGND VPWR VPWR _28127_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16071_ _17853_/A VGND VGND VPWR VPWR _16071_/X sky130_fd_sc_hd__buf_2
XFILLER_202_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28057_ _28057_/A VGND VGND VPWR VPWR _34359_/D sky130_fd_sc_hd__clkbuf_1
X_25269_ _25269_/A VGND VGND VPWR VPWR _33075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27008_ input57/X VGND VGND VPWR VPWR _27008_/X sky130_fd_sc_hd__buf_2
XFILLER_6_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19830_ _19716_/X _19828_/X _19829_/X _19720_/X VGND VGND VPWR VPWR _19830_/X sky130_fd_sc_hd__a22o_1
XFILLER_233_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19761_ _33205_/Q _32565_/Q _35957_/Q _35893_/Q _19727_/X _19728_/X VGND VGND VPWR
+ VPWR _19761_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16973_ _35047_/Q _34983_/Q _34919_/Q _34855_/Q _16803_/X _16804_/X VGND VGND VPWR
+ VPWR _16973_/X sky130_fd_sc_hd__mux4_1
X_28959_ _34787_/Q _24311_/X _28975_/S VGND VGND VPWR VPWR _28960_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18712_ _18712_/A _18712_/B _18712_/C _18712_/D VGND VGND VPWR VPWR _18713_/A sky130_fd_sc_hd__or4_4
XTAP_5050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31970_ _34970_/CLK _31970_/D VGND VGND VPWR VPWR _31970_/Q sky130_fd_sc_hd__dfxtp_1
X_19692_ _34803_/Q _34739_/Q _34675_/Q _34611_/Q _19588_/X _19589_/X VGND VGND VPWR
+ VPWR _19692_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 DW[17] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__buf_6
X_18643_ _34262_/Q _34198_/Q _34134_/Q _34070_/Q _18305_/X _18307_/X VGND VGND VPWR
+ VPWR _18643_/X sky130_fd_sc_hd__mux4_1
XTAP_5094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30921_ _30921_/A VGND VGND VPWR VPWR _35685_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33640_ _34279_/CLK _33640_/D VGND VGND VPWR VPWR _33640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18574_ _18436_/X _18572_/X _18573_/X _18441_/X VGND VGND VPWR VPWR _18574_/X sky130_fd_sc_hd__a22o_1
X_30852_ _23319_/X _35653_/Q _30860_/S VGND VGND VPWR VPWR _30853_/A sky130_fd_sc_hd__mux2_1
XTAP_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17525_ _32759_/Q _32695_/Q _32631_/Q _36087_/Q _17272_/X _17409_/X VGND VGND VPWR
+ VPWR _17525_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33571_ _33635_/CLK _33571_/D VGND VGND VPWR VPWR _33571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30783_ _23175_/X _35620_/Q _30797_/S VGND VGND VPWR VPWR _30784_/A sky130_fd_sc_hd__mux2_1
XFILLER_233_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_670 _22460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35310_ _35564_/CLK _35310_/D VGND VGND VPWR VPWR _35310_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32522_ _36170_/CLK _32522_/D VGND VGND VPWR VPWR _32522_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_681 _22557_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_692 _22595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17456_ _17452_/X _17455_/X _17136_/X _17137_/X VGND VGND VPWR VPWR _17471_/B sky130_fd_sc_hd__o211a_1
XFILLER_20_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16407_ _16074_/X _16405_/X _16406_/X _16084_/X VGND VGND VPWR VPWR _16407_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35241_ _35307_/CLK _35241_/D VGND VGND VPWR VPWR _35241_/Q sky130_fd_sc_hd__dfxtp_1
X_32453_ _35779_/CLK _32453_/D VGND VGND VPWR VPWR _32453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17387_ _17347_/X _17385_/X _17386_/X _17350_/X VGND VGND VPWR VPWR _17387_/X sky130_fd_sc_hd__a22o_1
XFILLER_220_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31404_ _35915_/Q input58/X _31408_/S VGND VGND VPWR VPWR _31405_/A sky130_fd_sc_hd__mux2_1
X_19126_ _35811_/Q _32187_/Q _35683_/Q _35619_/Q _18907_/X _18908_/X VGND VGND VPWR
+ VPWR _19126_/X sky130_fd_sc_hd__mux4_1
X_16338_ _16087_/X _16336_/X _16337_/X _16097_/X VGND VGND VPWR VPWR _16338_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35172_ _36003_/CLK _35172_/D VGND VGND VPWR VPWR _35172_/Q sky130_fd_sc_hd__dfxtp_1
X_32384_ _36032_/CLK _32384_/D VGND VGND VPWR VPWR _32384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34123_ _35273_/CLK _34123_/D VGND VGND VPWR VPWR _34123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19057_ _19053_/X _19056_/X _18741_/X VGND VGND VPWR VPWR _19065_/C sky130_fd_sc_hd__o21ba_1
X_31335_ _35882_/Q input21/X _31337_/S VGND VGND VPWR VPWR _31336_/A sky130_fd_sc_hd__mux2_1
X_16269_ _16265_/X _16268_/X _16100_/X VGND VGND VPWR VPWR _16270_/D sky130_fd_sc_hd__o21ba_1
X_18008_ _33541_/Q _33477_/Q _33413_/Q _33349_/Q _17829_/X _17830_/X VGND VGND VPWR
+ VPWR _18008_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34054_ _34057_/CLK _34054_/D VGND VGND VPWR VPWR _34054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31266_ _31266_/A VGND VGND VPWR VPWR _35849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33005_ _33007_/CLK _33005_/D VGND VGND VPWR VPWR _33005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30217_ _35352_/Q _29082_/X _30235_/S VGND VGND VPWR VPWR _30218_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31197_ _31197_/A VGND VGND VPWR VPWR _35816_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19959_ _32763_/Q _32699_/Q _32635_/Q _36091_/Q _19925_/X _19709_/X VGND VGND VPWR
+ VPWR _19959_/X sky130_fd_sc_hd__mux4_1
X_30148_ _30148_/A VGND VGND VPWR VPWR _35319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34956_ _35853_/CLK _34956_/D VGND VGND VPWR VPWR _34956_/Q sky130_fd_sc_hd__dfxtp_1
X_22970_ _22969_/X _32043_/Q _22970_/S VGND VGND VPWR VPWR _22971_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30079_ _35287_/Q _29079_/X _30079_/S VGND VGND VPWR VPWR _30080_/A sky130_fd_sc_hd__mux2_1
XANTENNA_1080 _17194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1091 _17264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21921_ _21917_/X _21920_/X _21747_/X VGND VGND VPWR VPWR _21929_/C sky130_fd_sc_hd__o21ba_1
XFILLER_110_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33907_ _34228_/CLK _33907_/D VGND VGND VPWR VPWR _33907_/Q sky130_fd_sc_hd__dfxtp_1
X_34887_ _35079_/CLK _34887_/D VGND VGND VPWR VPWR _34887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24640_ _22963_/X _32809_/Q _24644_/S VGND VGND VPWR VPWR _24641_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33838_ _35758_/CLK _33838_/D VGND VGND VPWR VPWR _33838_/Q sky130_fd_sc_hd__dfxtp_1
X_21852_ _35567_/Q _35503_/Q _35439_/Q _35375_/Q _21850_/X _21851_/X VGND VGND VPWR
+ VPWR _21852_/X sky130_fd_sc_hd__mux4_1
XFILLER_167_1138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20803_ _20799_/X _20802_/X _20700_/X VGND VGND VPWR VPWR _20804_/D sky130_fd_sc_hd__o21ba_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24571_ _23065_/X _32778_/Q _24577_/S VGND VGND VPWR VPWR _24572_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21783_ _33197_/Q _32557_/Q _35949_/Q _35885_/Q _21674_/X _21675_/X VGND VGND VPWR
+ VPWR _21783_/X sky130_fd_sc_hd__mux4_1
X_33769_ _34154_/CLK _33769_/D VGND VGND VPWR VPWR _33769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23522_ _23019_/X _32315_/Q _23530_/S VGND VGND VPWR VPWR _23523_/A sky130_fd_sc_hd__mux2_1
X_26310_ _25035_/X _33564_/Q _26320_/S VGND VGND VPWR VPWR _26311_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20734_ _20734_/A _20734_/B _20734_/C _20734_/D VGND VGND VPWR VPWR _20735_/A sky130_fd_sc_hd__or4_4
X_27290_ _27290_/A VGND VGND VPWR VPWR _33997_/D sky130_fd_sc_hd__clkbuf_1
X_35508_ _35956_/CLK _35508_/D VGND VGND VPWR VPWR _35508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26241_ _26241_/A VGND VGND VPWR VPWR _33531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35439_ _35951_/CLK _35439_/D VGND VGND VPWR VPWR _35439_/Q sky130_fd_sc_hd__dfxtp_1
X_23453_ _22917_/X _32282_/Q _23467_/S VGND VGND VPWR VPWR _23454_/A sky130_fd_sc_hd__mux2_1
X_20665_ _22532_/A VGND VGND VPWR VPWR _20665_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_50_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22404_ _33279_/Q _36159_/Q _33151_/Q _33087_/Q _22364_/X _22365_/X VGND VGND VPWR
+ VPWR _22404_/X sky130_fd_sc_hd__mux4_1
XFILLER_167_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26172_ _26172_/A VGND VGND VPWR VPWR _33498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23384_ _32251_/Q _23286_/X _23392_/S VGND VGND VPWR VPWR _23385_/A sky130_fd_sc_hd__mux2_1
X_20596_ _22369_/A VGND VGND VPWR VPWR _22460_/A sky130_fd_sc_hd__buf_12
XFILLER_137_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25123_ _25122_/X _33016_/Q _25144_/S VGND VGND VPWR VPWR _25124_/A sky130_fd_sc_hd__mux2_1
X_22335_ _33021_/Q _32957_/Q _32893_/Q _32829_/Q _22295_/X _22296_/X VGND VGND VPWR
+ VPWR _22335_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29931_ _29931_/A VGND VGND VPWR VPWR _35216_/D sky130_fd_sc_hd__clkbuf_1
X_25054_ _25187_/S VGND VGND VPWR VPWR _25082_/S sky130_fd_sc_hd__buf_4
X_22266_ _22395_/A VGND VGND VPWR VPWR _22266_/X sky130_fd_sc_hd__buf_6
XFILLER_191_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24005_ _24005_/A VGND VGND VPWR VPWR _32540_/D sky130_fd_sc_hd__clkbuf_1
X_21217_ _35293_/Q _35229_/Q _35165_/Q _32285_/Q _20900_/X _20901_/X VGND VGND VPWR
+ VPWR _21217_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29862_ _35184_/Q _29157_/X _29872_/S VGND VGND VPWR VPWR _29863_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22197_ _33017_/Q _32953_/Q _32889_/Q _32825_/Q _21942_/X _21943_/X VGND VGND VPWR
+ VPWR _22197_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28813_ _26872_/X _34718_/Q _28819_/S VGND VGND VPWR VPWR _28814_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21148_ _20893_/X _21146_/X _21147_/X _20896_/X VGND VGND VPWR VPWR _21148_/X sky130_fd_sc_hd__a22o_1
X_29793_ _35151_/Q _29055_/X _29809_/S VGND VGND VPWR VPWR _29794_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28744_ _28744_/A VGND VGND VPWR VPWR _34685_/D sky130_fd_sc_hd__clkbuf_1
X_21079_ _21075_/X _21078_/X _21041_/X VGND VGND VPWR VPWR _21087_/C sky130_fd_sc_hd__o21ba_2
X_25956_ _25956_/A VGND VGND VPWR VPWR _33396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24907_ _24907_/A VGND VGND VPWR VPWR _32934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28675_ _28675_/A VGND VGND VPWR VPWR _34652_/D sky130_fd_sc_hd__clkbuf_1
X_25887_ _25887_/A VGND VGND VPWR VPWR _33363_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27626_ _27626_/A VGND VGND VPWR VPWR _34155_/D sky130_fd_sc_hd__clkbuf_1
X_24838_ _23053_/X _32902_/Q _24844_/S VGND VGND VPWR VPWR _24839_/A sky130_fd_sc_hd__mux2_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27557_ _27014_/X _34124_/Q _27559_/S VGND VGND VPWR VPWR _27558_/A sky130_fd_sc_hd__mux2_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24769_ _22951_/X _32869_/Q _24781_/S VGND VGND VPWR VPWR _24770_/A sky130_fd_sc_hd__mux2_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17310_ _33009_/Q _32945_/Q _32881_/Q _32817_/Q _16989_/X _16990_/X VGND VGND VPWR
+ VPWR _17310_/X sky130_fd_sc_hd__mux4_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26508_ _25128_/X _33658_/Q _26518_/S VGND VGND VPWR VPWR _26509_/A sky130_fd_sc_hd__mux2_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18290_ _18359_/A VGND VGND VPWR VPWR _20096_/A sky130_fd_sc_hd__buf_12
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27488_ _26912_/X _34091_/Q _27488_/S VGND VGND VPWR VPWR _27489_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29227_ _29227_/A VGND VGND VPWR VPWR _34886_/D sky130_fd_sc_hd__clkbuf_1
X_17241_ _33263_/Q _36143_/Q _33135_/Q _33071_/Q _17058_/X _17059_/X VGND VGND VPWR
+ VPWR _17241_/X sky130_fd_sc_hd__mux4_1
XFILLER_230_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26439_ _25026_/X _33625_/Q _26455_/S VGND VGND VPWR VPWR _26440_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29158_ _34864_/Q _29157_/X _29173_/S VGND VGND VPWR VPWR _29159_/A sky130_fd_sc_hd__mux2_1
X_17172_ _32749_/Q _32685_/Q _32621_/Q _36077_/Q _16919_/X _17056_/X VGND VGND VPWR
+ VPWR _17172_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16123_ _35535_/Q _35471_/Q _35407_/Q _35343_/Q _16058_/X _16060_/X VGND VGND VPWR
+ VPWR _16123_/X sky130_fd_sc_hd__mux4_1
X_28109_ _26829_/X _34384_/Q _28123_/S VGND VGND VPWR VPWR _28110_/A sky130_fd_sc_hd__mux2_1
X_29089_ input4/X VGND VGND VPWR VPWR _29089_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_182_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31120_ _35780_/Q _29219_/X _31130_/S VGND VGND VPWR VPWR _31121_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16054_ _17858_/A VGND VGND VPWR VPWR _16054_/X sky130_fd_sc_hd__buf_4
XFILLER_51_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31051_ _35747_/Q _29117_/X _31067_/S VGND VGND VPWR VPWR _31052_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19813_ _19807_/X _19808_/X _19811_/X _19812_/X VGND VGND VPWR VPWR _19813_/X sky130_fd_sc_hd__a22o_1
X_30002_ _30002_/A VGND VGND VPWR VPWR _35250_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_1239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34810_ _35771_/CLK _34810_/D VGND VGND VPWR VPWR _34810_/Q sky130_fd_sc_hd__dfxtp_1
X_19744_ _34293_/Q _34229_/Q _34165_/Q _34101_/Q _19742_/X _19743_/X VGND VGND VPWR
+ VPWR _19744_/X sky130_fd_sc_hd__mux4_1
X_35790_ _35793_/CLK _35790_/D VGND VGND VPWR VPWR _35790_/Q sky130_fd_sc_hd__dfxtp_1
X_16956_ _32487_/Q _32359_/Q _32039_/Q _36007_/Q _16923_/X _16711_/X VGND VGND VPWR
+ VPWR _16956_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34741_ _35250_/CLK _34741_/D VGND VGND VPWR VPWR _34741_/Q sky130_fd_sc_hd__dfxtp_1
X_31953_ _34973_/CLK _31953_/D VGND VGND VPWR VPWR _31953_/Q sky130_fd_sc_hd__dfxtp_1
X_19675_ _34035_/Q _33971_/Q _33907_/Q _32243_/Q _19673_/X _19674_/X VGND VGND VPWR
+ VPWR _19675_/X sky130_fd_sc_hd__mux4_1
X_16887_ _32741_/Q _32677_/Q _32613_/Q _36069_/Q _16566_/X _16703_/X VGND VGND VPWR
+ VPWR _16887_/X sky130_fd_sc_hd__mux4_1
X_18626_ _35797_/Q _32172_/Q _35669_/Q _35605_/Q _18554_/X _18555_/X VGND VGND VPWR
+ VPWR _18626_/X sky130_fd_sc_hd__mux4_1
X_30904_ _30904_/A VGND VGND VPWR VPWR _35677_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34672_ _34797_/CLK _34672_/D VGND VGND VPWR VPWR _34672_/Q sky130_fd_sc_hd__dfxtp_1
X_31884_ _23244_/X _36142_/Q _31898_/S VGND VGND VPWR VPWR _31885_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33623_ _35215_/CLK _33623_/D VGND VGND VPWR VPWR _33623_/Q sky130_fd_sc_hd__dfxtp_1
X_18557_ _35731_/Q _35091_/Q _34451_/Q _33811_/Q _18349_/X _18351_/X VGND VGND VPWR
+ VPWR _18557_/X sky130_fd_sc_hd__mux4_1
X_30835_ _23294_/X _35645_/Q _30839_/S VGND VGND VPWR VPWR _30836_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17508_ _34550_/Q _32438_/Q _34422_/Q _34358_/Q _17225_/X _17226_/X VGND VGND VPWR
+ VPWR _17508_/X sky130_fd_sc_hd__mux4_1
X_33554_ _34194_/CLK _33554_/D VGND VGND VPWR VPWR _33554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18488_ _35793_/Q _32167_/Q _35665_/Q _35601_/Q _18345_/X _18346_/X VGND VGND VPWR
+ VPWR _18488_/X sky130_fd_sc_hd__mux4_1
X_30766_ _23130_/X _35612_/Q _30776_/S VGND VGND VPWR VPWR _30767_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32505_ _36025_/CLK _32505_/D VGND VGND VPWR VPWR _32505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_14 _32115_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17439_ _17439_/A _17439_/B _17439_/C _17439_/D VGND VGND VPWR VPWR _17440_/A sky130_fd_sc_hd__or4_4
X_33485_ _35984_/CLK _33485_/D VGND VGND VPWR VPWR _33485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_25 _32116_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_221_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30697_ _30697_/A VGND VGND VPWR VPWR _35579_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_36 _32117_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_47 _32119_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35224_ _35226_/CLK _35224_/D VGND VGND VPWR VPWR _35224_/Q sky130_fd_sc_hd__dfxtp_1
X_20450_ _35081_/Q _35017_/Q _34953_/Q _34889_/Q _20162_/X _20163_/X VGND VGND VPWR
+ VPWR _20450_/X sky130_fd_sc_hd__mux4_1
XANTENNA_58 _32126_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32436_ _34805_/CLK _32436_/D VGND VGND VPWR VPWR _32436_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_69 _32127_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19109_ _19100_/X _19107_/X _19108_/X VGND VGND VPWR VPWR _19110_/D sky130_fd_sc_hd__o21ba_1
X_35155_ _36216_/CLK _35155_/D VGND VGND VPWR VPWR _35155_/Q sky130_fd_sc_hd__dfxtp_1
X_20381_ _18277_/X _20379_/X _20380_/X _18287_/X VGND VGND VPWR VPWR _20381_/X sky130_fd_sc_hd__a22o_1
X_32367_ _36015_/CLK _32367_/D VGND VGND VPWR VPWR _32367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34106_ _36154_/CLK _34106_/D VGND VGND VPWR VPWR _34106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1060 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22120_ _21795_/X _22118_/X _22119_/X _21800_/X VGND VGND VPWR VPWR _22120_/X sky130_fd_sc_hd__a22o_1
X_31318_ _31408_/S VGND VGND VPWR VPWR _31337_/S sky130_fd_sc_hd__buf_4
X_35086_ _35728_/CLK _35086_/D VGND VGND VPWR VPWR _35086_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput110 _31978_/Q VGND VGND VPWR VPWR D1[28] sky130_fd_sc_hd__buf_2
X_32298_ _34794_/CLK _32298_/D VGND VGND VPWR VPWR _32298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput121 _31988_/Q VGND VGND VPWR VPWR D1[38] sky130_fd_sc_hd__buf_2
XFILLER_217_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput132 _31998_/Q VGND VGND VPWR VPWR D1[48] sky130_fd_sc_hd__buf_2
Xoutput143 _32008_/Q VGND VGND VPWR VPWR D1[58] sky130_fd_sc_hd__buf_2
X_34037_ _34229_/CLK _34037_/D VGND VGND VPWR VPWR _34037_/Q sky130_fd_sc_hd__dfxtp_1
X_22051_ _33269_/Q _36149_/Q _33141_/Q _33077_/Q _22011_/X _22012_/X VGND VGND VPWR
+ VPWR _22051_/X sky130_fd_sc_hd__mux4_1
XTAP_6509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31249_ _35841_/Q input47/X _31265_/S VGND VGND VPWR VPWR _31250_/A sky130_fd_sc_hd__mux2_1
Xoutput154 _36174_/Q VGND VGND VPWR VPWR D2[0] sky130_fd_sc_hd__buf_2
Xoutput165 _36175_/Q VGND VGND VPWR VPWR D2[1] sky130_fd_sc_hd__buf_2
XFILLER_88_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21002_ _33175_/Q _32535_/Q _35927_/Q _35863_/Q _20968_/X _20969_/X VGND VGND VPWR
+ VPWR _21002_/X sky130_fd_sc_hd__mux4_1
Xoutput176 _36176_/Q VGND VGND VPWR VPWR D2[2] sky130_fd_sc_hd__buf_2
Xoutput187 _36177_/Q VGND VGND VPWR VPWR D2[3] sky130_fd_sc_hd__buf_2
XFILLER_87_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput198 _36178_/Q VGND VGND VPWR VPWR D2[4] sky130_fd_sc_hd__buf_2
XTAP_5819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25810_ _25094_/X _33327_/Q _25822_/S VGND VGND VPWR VPWR _25811_/A sky130_fd_sc_hd__mux2_1
X_26790_ _33791_/Q _24397_/X _26790_/S VGND VGND VPWR VPWR _26791_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35988_ _35989_/CLK _35988_/D VGND VGND VPWR VPWR _35988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25741_ _24989_/X _33294_/Q _25759_/S VGND VGND VPWR VPWR _25742_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22953_ _22953_/A VGND VGND VPWR VPWR _32037_/D sky130_fd_sc_hd__clkbuf_1
X_34939_ _35515_/CLK _34939_/D VGND VGND VPWR VPWR _34939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21904_ _21802_/X _21902_/X _21903_/X _21805_/X VGND VGND VPWR VPWR _21904_/X sky130_fd_sc_hd__a22o_1
XFILLER_56_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28460_ _28460_/A VGND VGND VPWR VPWR _34550_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22884_ _22883_/X _32015_/Q _22908_/S VGND VGND VPWR VPWR _22885_/A sky130_fd_sc_hd__mux2_1
X_25672_ _25672_/A VGND VGND VPWR VPWR _33262_/D sky130_fd_sc_hd__clkbuf_1
X_27411_ _27411_/A VGND VGND VPWR VPWR _34054_/D sky130_fd_sc_hd__clkbuf_1
X_21835_ _21795_/X _21833_/X _21834_/X _21800_/X VGND VGND VPWR VPWR _21835_/X sky130_fd_sc_hd__a22o_1
X_24623_ _22938_/X _32801_/Q _24623_/S VGND VGND VPWR VPWR _24624_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28391_ _26847_/X _34518_/Q _28393_/S VGND VGND VPWR VPWR _28392_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24554_ _24554_/A VGND VGND VPWR VPWR _32769_/D sky130_fd_sc_hd__clkbuf_1
X_27342_ _27342_/A VGND VGND VPWR VPWR _34021_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21766_ _34285_/Q _34221_/Q _34157_/Q _34093_/Q _21689_/X _21690_/X VGND VGND VPWR
+ VPWR _21766_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20717_ _32975_/Q _32911_/Q _32847_/Q _32783_/Q _20633_/X _20635_/X VGND VGND VPWR
+ VPWR _20717_/X sky130_fd_sc_hd__mux4_1
X_23505_ _22994_/X _32307_/Q _23509_/S VGND VGND VPWR VPWR _23506_/A sky130_fd_sc_hd__mux2_1
X_27273_ _26993_/X _33989_/Q _27281_/S VGND VGND VPWR VPWR _27274_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24485_ _22938_/X _32737_/Q _24485_/S VGND VGND VPWR VPWR _24486_/A sky130_fd_sc_hd__mux2_1
X_21697_ _32747_/Q _32683_/Q _32619_/Q _36075_/Q _21519_/X _21656_/X VGND VGND VPWR
+ VPWR _21697_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29012_ _29012_/A VGND VGND VPWR VPWR _34812_/D sky130_fd_sc_hd__clkbuf_1
X_23436_ _22892_/X _32274_/Q _23446_/S VGND VGND VPWR VPWR _23437_/A sky130_fd_sc_hd__mux2_1
X_26224_ _26224_/A VGND VGND VPWR VPWR _33523_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20648_ _22578_/A VGND VGND VPWR VPWR _22594_/A sky130_fd_sc_hd__buf_12
X_26155_ _26155_/A VGND VGND VPWR VPWR _33490_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_192_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _35326_/CLK sky130_fd_sc_hd__clkbuf_16
X_23367_ _32243_/Q _23261_/X _23371_/S VGND VGND VPWR VPWR _23368_/A sky130_fd_sc_hd__mux2_1
X_20579_ _20657_/A VGND VGND VPWR VPWR _22502_/A sky130_fd_sc_hd__buf_12
XFILLER_165_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1064 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22318_ _22107_/X _22316_/X _22317_/X _22112_/X VGND VGND VPWR VPWR _22318_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_1160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25106_ input31/X VGND VGND VPWR VPWR _25106_/X sky130_fd_sc_hd__clkbuf_4
X_26086_ _25103_/X _33458_/Q _26092_/S VGND VGND VPWR VPWR _26087_/A sky130_fd_sc_hd__mux2_1
X_23298_ _32217_/Q _23297_/X _23301_/S VGND VGND VPWR VPWR _23299_/A sky130_fd_sc_hd__mux2_1
X_29914_ _35209_/Q _29234_/X _29914_/S VGND VGND VPWR VPWR _29915_/A sky130_fd_sc_hd__mux2_1
X_25037_ _25037_/A VGND VGND VPWR VPWR _32988_/D sky130_fd_sc_hd__clkbuf_1
X_22249_ _22245_/X _22248_/X _22114_/X VGND VGND VPWR VPWR _22250_/D sky130_fd_sc_hd__o21ba_1
XFILLER_124_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_1351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29845_ _35176_/Q _29132_/X _29851_/S VGND VGND VPWR VPWR _29846_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16810_ _16810_/A _16810_/B _16810_/C _16810_/D VGND VGND VPWR VPWR _16811_/A sky130_fd_sc_hd__or4_4
X_29776_ _29776_/A VGND VGND VPWR VPWR _35143_/D sky130_fd_sc_hd__clkbuf_1
X_17790_ _17507_/X _17788_/X _17789_/X _17512_/X VGND VGND VPWR VPWR _17790_/X sky130_fd_sc_hd__a22o_1
X_26988_ _26987_/X _33859_/Q _27006_/S VGND VGND VPWR VPWR _26989_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28727_ _28727_/A VGND VGND VPWR VPWR _34677_/D sky130_fd_sc_hd__clkbuf_1
X_16741_ _34017_/Q _33953_/Q _33889_/Q _32161_/Q _16667_/X _16668_/X VGND VGND VPWR
+ VPWR _16741_/X sky130_fd_sc_hd__mux4_1
XFILLER_207_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25939_ _25084_/X _33388_/Q _25957_/S VGND VGND VPWR VPWR _25940_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19460_ _19454_/X _19455_/X _19458_/X _19459_/X VGND VGND VPWR VPWR _19460_/X sky130_fd_sc_hd__a22o_1
X_28658_ _28658_/A VGND VGND VPWR VPWR _34644_/D sky130_fd_sc_hd__clkbuf_1
X_16672_ _32735_/Q _32671_/Q _32607_/Q _36063_/Q _16566_/X _16350_/X VGND VGND VPWR
+ VPWR _16672_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_6_25__f_CLK clkbuf_5_12_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_76_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_62_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18411_ _18297_/X _18407_/X _18410_/X _18303_/X VGND VGND VPWR VPWR _18411_/X sky130_fd_sc_hd__a22o_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27609_ _34147_/Q _24311_/X _27625_/S VGND VGND VPWR VPWR _27610_/A sky130_fd_sc_hd__mux2_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19391_ _34283_/Q _34219_/Q _34155_/Q _34091_/Q _19389_/X _19390_/X VGND VGND VPWR
+ VPWR _19391_/X sky130_fd_sc_hd__mux4_1
X_28589_ _26940_/X _34612_/Q _28591_/S VGND VGND VPWR VPWR _28590_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_1303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30620_ _35543_/Q _29079_/X _30620_/S VGND VGND VPWR VPWR _30621_/A sky130_fd_sc_hd__mux2_1
X_18342_ _20143_/A VGND VGND VPWR VPWR _18342_/X sky130_fd_sc_hd__buf_2
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18273_ _18273_/A _18273_/B _18273_/C _18273_/D VGND VGND VPWR VPWR _18274_/A sky130_fd_sc_hd__or4_4
XFILLER_30_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30551_ _23270_/X _35510_/Q _30569_/S VGND VGND VPWR VPWR _30552_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17224_ _17149_/X _17222_/X _17223_/X _17152_/X VGND VGND VPWR VPWR _17224_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33270_ _36150_/CLK _33270_/D VGND VGND VPWR VPWR _33270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30482_ _30482_/A VGND VGND VPWR VPWR _35477_/D sky130_fd_sc_hd__clkbuf_1
Xinput12 DW[1] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__buf_8
Xinput23 DW[2] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__buf_8
X_32221_ _35843_/CLK _32221_/D VGND VGND VPWR VPWR _32221_/Q sky130_fd_sc_hd__dfxtp_1
Xinput34 DW[3] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__buf_8
Xinput45 DW[4] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__buf_6
X_17155_ _34540_/Q _32428_/Q _34412_/Q _34348_/Q _16872_/X _16873_/X VGND VGND VPWR
+ VPWR _17155_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_183_CLK clkbuf_leaf_66_CLK/A VGND VGND VPWR VPWR _35986_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput56 DW[5] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__buf_8
Xinput67 R1[2] VGND VGND VPWR VPWR input67/X sky130_fd_sc_hd__buf_6
XFILLER_183_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput78 R3[1] VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__clkbuf_2
XFILLER_239_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16106_ _15977_/X _16104_/X _16105_/X _15987_/X VGND VGND VPWR VPWR _16106_/X sky130_fd_sc_hd__a22o_1
Xinput89 WE VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__buf_6
XFILLER_183_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32152_ _34267_/CLK _32152_/D VGND VGND VPWR VPWR _32152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17086_ _17086_/A _17086_/B _17086_/C _17086_/D VGND VGND VPWR VPWR _17087_/A sky130_fd_sc_hd__or4_4
XFILLER_66_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31103_ _35772_/Q _29194_/X _31109_/S VGND VGND VPWR VPWR _31104_/A sky130_fd_sc_hd__mux2_1
X_16037_ _17911_/A VGND VGND VPWR VPWR _16037_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32083_ _35038_/CLK _32083_/D VGND VGND VPWR VPWR _32083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35911_ _36168_/CLK _35911_/D VGND VGND VPWR VPWR _35911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31034_ _35739_/Q _29092_/X _31046_/S VGND VGND VPWR VPWR _31035_/A sky130_fd_sc_hd__mux2_1
XFILLER_233_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35842_ _36038_/CLK _35842_/D VGND VGND VPWR VPWR _35842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17988_ _35780_/Q _35140_/Q _34500_/Q _33860_/Q _17846_/X _17847_/X VGND VGND VPWR
+ VPWR _17988_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19727_ _20231_/A VGND VGND VPWR VPWR _19727_/X sky130_fd_sc_hd__buf_6
XFILLER_211_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16939_ _16796_/X _16937_/X _16938_/X _16799_/X VGND VGND VPWR VPWR _16939_/X sky130_fd_sc_hd__a22o_1
X_35773_ _35837_/CLK _35773_/D VGND VGND VPWR VPWR _35773_/Q sky130_fd_sc_hd__dfxtp_1
X_32985_ _36119_/CLK _32985_/D VGND VGND VPWR VPWR _32985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31936_ _23327_/X _36167_/Q _31940_/S VGND VGND VPWR VPWR _31937_/A sky130_fd_sc_hd__mux2_1
X_34724_ _35928_/CLK _34724_/D VGND VGND VPWR VPWR _34724_/Q sky130_fd_sc_hd__dfxtp_1
X_19658_ _34802_/Q _34738_/Q _34674_/Q _34610_/Q _19588_/X _19589_/X VGND VGND VPWR
+ VPWR _19658_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18609_ _18609_/A VGND VGND VPWR VPWR _32084_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34655_ _34782_/CLK _34655_/D VGND VGND VPWR VPWR _34655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19589_ _20295_/A VGND VGND VPWR VPWR _19589_/X sky130_fd_sc_hd__buf_4
X_31867_ _23217_/X _36134_/Q _31877_/S VGND VGND VPWR VPWR _31868_/A sky130_fd_sc_hd__mux2_1
XFILLER_209_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33606_ _34312_/CLK _33606_/D VGND VGND VPWR VPWR _33606_/Q sky130_fd_sc_hd__dfxtp_1
X_21620_ _22446_/A VGND VGND VPWR VPWR _21620_/X sky130_fd_sc_hd__buf_6
X_30818_ _23267_/X _35637_/Q _30818_/S VGND VGND VPWR VPWR _30819_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34586_ _36201_/CLK _34586_/D VGND VGND VPWR VPWR _34586_/Q sky130_fd_sc_hd__dfxtp_1
X_31798_ _31798_/A VGND VGND VPWR VPWR _36101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33537_ _34305_/CLK _33537_/D VGND VGND VPWR VPWR _33537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21551_ _21449_/X _21549_/X _21550_/X _21452_/X VGND VGND VPWR VPWR _21551_/X sky130_fd_sc_hd__a22o_1
X_30749_ _23105_/X _35604_/Q _30755_/S VGND VGND VPWR VPWR _30750_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20502_ _35595_/Q _35531_/Q _35467_/Q _35403_/Q _20256_/X _20257_/X VGND VGND VPWR
+ VPWR _20502_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24270_ input63/X VGND VGND VPWR VPWR _24270_/X sky130_fd_sc_hd__buf_6
X_33468_ _33723_/CLK _33468_/D VGND VGND VPWR VPWR _33468_/Q sky130_fd_sc_hd__dfxtp_1
X_21482_ _21442_/X _21480_/X _21481_/X _21447_/X VGND VGND VPWR VPWR _21482_/X sky130_fd_sc_hd__a22o_1
XFILLER_222_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35207_ _35339_/CLK _35207_/D VGND VGND VPWR VPWR _35207_/Q sky130_fd_sc_hd__dfxtp_1
X_23221_ _32191_/Q _23220_/X _23235_/S VGND VGND VPWR VPWR _23222_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20433_ _33289_/Q _36169_/Q _33161_/Q _33097_/Q _18328_/X _19457_/A VGND VGND VPWR
+ VPWR _20433_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32419_ _35298_/CLK _32419_/D VGND VGND VPWR VPWR _32419_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_174_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _36049_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_147_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36187_ _36202_/CLK _36187_/D VGND VGND VPWR VPWR _36187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33399_ _34297_/CLK _33399_/D VGND VGND VPWR VPWR _33399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35138_ _35779_/CLK _35138_/D VGND VGND VPWR VPWR _35138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23152_ input14/X VGND VGND VPWR VPWR _23152_/X sky130_fd_sc_hd__buf_4
X_20364_ _20364_/A VGND VGND VPWR VPWR _32134_/D sky130_fd_sc_hd__buf_4
XFILLER_31_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22103_ _34806_/Q _34742_/Q _34678_/Q _34614_/Q _21888_/X _21889_/X VGND VGND VPWR
+ VPWR _22103_/X sky130_fd_sc_hd__mux4_1
XTAP_7029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27960_ _34314_/Q _24431_/X _27966_/S VGND VGND VPWR VPWR _27961_/A sky130_fd_sc_hd__mux2_1
X_23083_ input83/X input89/X VGND VGND VPWR VPWR _26549_/C sky130_fd_sc_hd__nand2_8
X_35069_ _35989_/CLK _35069_/D VGND VGND VPWR VPWR _35069_/Q sky130_fd_sc_hd__dfxtp_1
X_20295_ _20295_/A VGND VGND VPWR VPWR _20295_/X sky130_fd_sc_hd__buf_4
XTAP_6306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26911_ _26911_/A VGND VGND VPWR VPWR _33834_/D sky130_fd_sc_hd__clkbuf_1
X_22034_ _21749_/X _22032_/X _22033_/X _21752_/X VGND VGND VPWR VPWR _22034_/X sky130_fd_sc_hd__a22o_1
XTAP_6339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27891_ _34281_/Q _24329_/X _27895_/S VGND VGND VPWR VPWR _27892_/A sky130_fd_sc_hd__mux2_1
XTAP_5616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29630_ _35074_/Q _29213_/X _29644_/S VGND VGND VPWR VPWR _29631_/A sky130_fd_sc_hd__mux2_1
XTAP_5627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26842_ _26841_/X _33812_/Q _26851_/S VGND VGND VPWR VPWR _26843_/A sky130_fd_sc_hd__mux2_1
XTAP_5649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29561_ _29561_/A VGND VGND VPWR VPWR _35041_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26773_ _26773_/A VGND VGND VPWR VPWR _33782_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23985_ _22895_/X _32531_/Q _23993_/S VGND VGND VPWR VPWR _23986_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28512_ _26826_/X _34575_/Q _28528_/S VGND VGND VPWR VPWR _28513_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25724_ _25724_/A VGND VGND VPWR VPWR _33287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_917 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29492_ _29492_/A VGND VGND VPWR VPWR _35008_/D sky130_fd_sc_hd__clkbuf_1
X_22936_ _22935_/X _32032_/Q _22939_/S VGND VGND VPWR VPWR _22937_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28443_ _28443_/A VGND VGND VPWR VPWR _34542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25655_ _25655_/A VGND VGND VPWR VPWR _33254_/D sky130_fd_sc_hd__clkbuf_1
X_22867_ _35341_/Q _35277_/Q _35213_/Q _32333_/Q _20688_/X _20690_/X VGND VGND VPWR
+ VPWR _22867_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24606_ _24606_/A VGND VGND VPWR VPWR _32792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28374_ _28506_/S VGND VGND VPWR VPWR _28393_/S sky130_fd_sc_hd__buf_6
X_21818_ _35566_/Q _35502_/Q _35438_/Q _35374_/Q _21497_/X _21498_/X VGND VGND VPWR
+ VPWR _21818_/X sky130_fd_sc_hd__mux4_1
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22798_ _22794_/X _22797_/X _22442_/A _22443_/A VGND VGND VPWR VPWR _22813_/B sky130_fd_sc_hd__o211a_1
X_25586_ _25586_/A VGND VGND VPWR VPWR _33223_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1030 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27325_ _27325_/A VGND VGND VPWR VPWR _34013_/D sky130_fd_sc_hd__clkbuf_1
XPHY_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24537_ _24537_/A VGND VGND VPWR VPWR _32761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21749_ _21749_/A VGND VGND VPWR VPWR _21749_/X sky130_fd_sc_hd__clkbuf_4
XPHY_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27256_ _26968_/X _33981_/Q _27260_/S VGND VGND VPWR VPWR _27257_/A sky130_fd_sc_hd__mux2_1
X_24468_ _24468_/A VGND VGND VPWR VPWR _32728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26207_ _26207_/A VGND VGND VPWR VPWR _33515_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_165_CLK clkbuf_6_30__f_CLK/X VGND VGND VPWR VPWR _35979_/CLK sky130_fd_sc_hd__clkbuf_16
X_23419_ _32268_/Q _23342_/X _23421_/S VGND VGND VPWR VPWR _23420_/A sky130_fd_sc_hd__mux2_1
X_24399_ _24399_/A VGND VGND VPWR VPWR _32703_/D sky130_fd_sc_hd__clkbuf_1
X_27187_ _26866_/X _33948_/Q _27197_/S VGND VGND VPWR VPWR _27188_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26138_ _25180_/X _33483_/Q _26142_/S VGND VGND VPWR VPWR _26139_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18960_ _18956_/X _18959_/X _18755_/X VGND VGND VPWR VPWR _18961_/D sky130_fd_sc_hd__o21ba_1
XFILLER_152_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26069_ _25078_/X _33450_/Q _26071_/S VGND VGND VPWR VPWR _26070_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17911_ _17911_/A VGND VGND VPWR VPWR _17911_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_3_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18891_ _18891_/A _18891_/B _18891_/C _18891_/D VGND VGND VPWR VPWR _18892_/A sky130_fd_sc_hd__or4_2
XTAP_6840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17842_ _17842_/A VGND VGND VPWR VPWR _17842_/X sky130_fd_sc_hd__buf_4
X_29828_ _35168_/Q _29107_/X _29830_/S VGND VGND VPWR VPWR _29829_/A sky130_fd_sc_hd__mux2_1
XTAP_6873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17773_ _17773_/A VGND VGND VPWR VPWR _17773_/X sky130_fd_sc_hd__clkbuf_4
X_29759_ _29759_/A VGND VGND VPWR VPWR _35135_/D sky130_fd_sc_hd__clkbuf_1
X_19512_ _33006_/Q _32942_/Q _32878_/Q _32814_/Q _19289_/X _19290_/X VGND VGND VPWR
+ VPWR _19512_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16724_ _16646_/X _16720_/X _16723_/X _16649_/X VGND VGND VPWR VPWR _16724_/X sky130_fd_sc_hd__a22o_1
X_32770_ _33026_/CLK _32770_/D VGND VGND VPWR VPWR _32770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19443_ _19294_/X _19439_/X _19442_/X _19297_/X VGND VGND VPWR VPWR _19443_/X sky130_fd_sc_hd__a22o_1
X_31721_ _36065_/Q input11/X _31721_/S VGND VGND VPWR VPWR _31722_/A sky130_fd_sc_hd__mux2_1
X_16655_ _35294_/Q _35230_/Q _35166_/Q _32286_/Q _16653_/X _16654_/X VGND VGND VPWR
+ VPWR _16655_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34440_ _35078_/CLK _34440_/D VGND VGND VPWR VPWR _34440_/Q sky130_fd_sc_hd__dfxtp_1
X_31652_ _36032_/Q input46/X _31670_/S VGND VGND VPWR VPWR _31653_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19374_ _20231_/A VGND VGND VPWR VPWR _19374_/X sky130_fd_sc_hd__buf_6
X_16586_ _16443_/X _16584_/X _16585_/X _16446_/X VGND VGND VPWR VPWR _16586_/X sky130_fd_sc_hd__a22o_1
X_18325_ _20069_/A VGND VGND VPWR VPWR _20208_/A sky130_fd_sc_hd__buf_12
X_30603_ _30603_/A VGND VGND VPWR VPWR _35534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34371_ _34562_/CLK _34371_/D VGND VGND VPWR VPWR _34371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31583_ _31583_/A VGND VGND VPWR VPWR _35999_/D sky130_fd_sc_hd__clkbuf_1
X_36110_ _36114_/CLK _36110_/D VGND VGND VPWR VPWR _36110_/Q sky130_fd_sc_hd__dfxtp_1
X_33322_ _33512_/CLK _33322_/D VGND VGND VPWR VPWR _33322_/Q sky130_fd_sc_hd__dfxtp_1
X_18256_ _33037_/Q _32973_/Q _32909_/Q _32845_/Q _15980_/X _15983_/X VGND VGND VPWR
+ VPWR _18256_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30534_ _23244_/X _35502_/Q _30548_/S VGND VGND VPWR VPWR _30535_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36041_ _36041_/CLK _36041_/D VGND VGND VPWR VPWR _36041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17207_ _17201_/X _17206_/X _17128_/X VGND VGND VPWR VPWR _17231_/A sky130_fd_sc_hd__o21ba_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33253_ _36135_/CLK _33253_/D VGND VGND VPWR VPWR _33253_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_156_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _35848_/CLK sky130_fd_sc_hd__clkbuf_16
X_18187_ _17901_/X _18185_/X _18186_/X _17906_/X VGND VGND VPWR VPWR _18187_/X sky130_fd_sc_hd__a22o_1
X_30465_ _30735_/A _30465_/B VGND VGND VPWR VPWR _30598_/S sky130_fd_sc_hd__nand2_8
XFILLER_8_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32204_ _36135_/CLK _32204_/D VGND VGND VPWR VPWR _32204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17138_ _17132_/X _17135_/X _17136_/X _17137_/X VGND VGND VPWR VPWR _17163_/B sky130_fd_sc_hd__o211a_1
X_33184_ _35938_/CLK _33184_/D VGND VGND VPWR VPWR _33184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30396_ _30396_/A VGND VGND VPWR VPWR _35436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32135_ _35750_/CLK _32135_/D VGND VGND VPWR VPWR _32135_/Q sky130_fd_sc_hd__dfxtp_1
X_17069_ _17062_/X _17068_/X _16783_/X _16784_/X VGND VGND VPWR VPWR _17086_/B sky130_fd_sc_hd__o211a_1
XFILLER_171_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32066_ _36034_/CLK _32066_/D VGND VGND VPWR VPWR _32066_/Q sky130_fd_sc_hd__dfxtp_1
X_20080_ _20231_/A VGND VGND VPWR VPWR _20080_/X sky130_fd_sc_hd__buf_6
XFILLER_134_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31017_ _35731_/Q _29067_/X _31025_/S VGND VGND VPWR VPWR _31018_/A sky130_fd_sc_hd__mux2_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35825_ _35954_/CLK _35825_/D VGND VGND VPWR VPWR _35825_/Q sky130_fd_sc_hd__dfxtp_1
X_23770_ _22979_/X _32430_/Q _23784_/S VGND VGND VPWR VPWR _23771_/A sky130_fd_sc_hd__mux2_1
X_20982_ _33751_/Q _33687_/Q _33623_/Q _33559_/Q _20737_/X _20738_/X VGND VGND VPWR
+ VPWR _20982_/X sky130_fd_sc_hd__mux4_1
X_32968_ _36107_/CLK _32968_/D VGND VGND VPWR VPWR _32968_/Q sky130_fd_sc_hd__dfxtp_1
X_35756_ _35758_/CLK _35756_/D VGND VGND VPWR VPWR _35756_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22721_ _22460_/X _22719_/X _22720_/X _22465_/X VGND VGND VPWR VPWR _22721_/X sky130_fd_sc_hd__a22o_1
X_34707_ _36196_/CLK _34707_/D VGND VGND VPWR VPWR _34707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31919_ _23300_/X _36159_/Q _31919_/S VGND VGND VPWR VPWR _31920_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32899_ _32965_/CLK _32899_/D VGND VGND VPWR VPWR _32899_/Q sky130_fd_sc_hd__dfxtp_1
X_35687_ _35815_/CLK _35687_/D VGND VGND VPWR VPWR _35687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25440_ _25159_/X _33156_/Q _25450_/S VGND VGND VPWR VPWR _25441_/A sky130_fd_sc_hd__mux2_1
X_22652_ _35590_/Q _35526_/Q _35462_/Q _35398_/Q _22556_/X _22557_/X VGND VGND VPWR
+ VPWR _22652_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34638_ _34638_/CLK _34638_/D VGND VGND VPWR VPWR _34638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21603_ _21599_/X _21600_/X _21601_/X _21602_/X VGND VGND VPWR VPWR _21603_/X sky130_fd_sc_hd__a22o_1
XFILLER_94_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34569_ _35080_/CLK _34569_/D VGND VGND VPWR VPWR _34569_/Q sky130_fd_sc_hd__dfxtp_1
X_22583_ _32516_/Q _32388_/Q _32068_/Q _36036_/Q _22582_/X _22370_/X VGND VGND VPWR
+ VPWR _22583_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_395_CLK clkbuf_6_34__f_CLK/X VGND VGND VPWR VPWR _35950_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25371_ _25057_/X _33123_/Q _25387_/S VGND VGND VPWR VPWR _25372_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27110_ _27110_/A VGND VGND VPWR VPWR _33911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21534_ _21530_/X _21533_/X _21394_/X VGND VGND VPWR VPWR _21544_/C sky130_fd_sc_hd__o21ba_1
X_24322_ _24322_/A VGND VGND VPWR VPWR _32678_/D sky130_fd_sc_hd__clkbuf_1
X_28090_ _28090_/A VGND VGND VPWR VPWR _34375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27041_ _26850_/X _33879_/Q _27041_/S VGND VGND VPWR VPWR _27042_/A sky130_fd_sc_hd__mux2_1
X_24253_ _32656_/Q _24252_/X _24274_/S VGND VGND VPWR VPWR _24254_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_147_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _35340_/CLK sky130_fd_sc_hd__clkbuf_16
X_21465_ _35556_/Q _35492_/Q _35428_/Q _35364_/Q _21144_/X _21145_/X VGND VGND VPWR
+ VPWR _21465_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23204_ _32184_/Q _23142_/X _23206_/S VGND VGND VPWR VPWR _23205_/A sky130_fd_sc_hd__mux2_1
X_20416_ _34824_/Q _34760_/Q _34696_/Q _34632_/Q _20294_/X _20295_/X VGND VGND VPWR
+ VPWR _20416_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24184_ _22988_/X _32625_/Q _24192_/S VGND VGND VPWR VPWR _24185_/A sky130_fd_sc_hd__mux2_1
X_21396_ _21749_/A VGND VGND VPWR VPWR _21396_/X sky130_fd_sc_hd__clkbuf_4
X_23135_ _23135_/A VGND VGND VPWR VPWR _32157_/D sky130_fd_sc_hd__clkbuf_1
X_20347_ _20069_/X _20345_/X _20346_/X _20073_/X VGND VGND VPWR VPWR _20347_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28992_ _34803_/Q _24360_/X _28996_/S VGND VGND VPWR VPWR _28993_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23066_ _23065_/X _32074_/Q _23075_/S VGND VGND VPWR VPWR _23067_/A sky130_fd_sc_hd__mux2_1
X_27943_ _27943_/A VGND VGND VPWR VPWR _34305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20278_ _20278_/A VGND VGND VPWR VPWR _20278_/X sky130_fd_sc_hd__buf_8
XFILLER_161_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22017_ _22370_/A VGND VGND VPWR VPWR _22017_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_89_975 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27874_ _34273_/Q _24304_/X _27874_/S VGND VGND VPWR VPWR _27875_/A sky130_fd_sc_hd__mux2_1
XTAP_5446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29613_ _35066_/Q _29188_/X _29623_/S VGND VGND VPWR VPWR _29614_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26825_ _26825_/A VGND VGND VPWR VPWR _33806_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29544_ _35033_/Q _29086_/X _29560_/S VGND VGND VPWR VPWR _29545_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26756_ _26756_/A VGND VGND VPWR VPWR _33774_/D sky130_fd_sc_hd__clkbuf_1
X_23968_ _23071_/X _32524_/Q _23970_/S VGND VGND VPWR VPWR _23969_/A sky130_fd_sc_hd__mux2_1
XTAP_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25707_ _25707_/A VGND VGND VPWR VPWR _33279_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29475_ _29475_/A VGND VGND VPWR VPWR _35000_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22919_ _22919_/A VGND VGND VPWR VPWR _32026_/D sky130_fd_sc_hd__clkbuf_1
X_26687_ _26819_/S VGND VGND VPWR VPWR _26706_/S sky130_fd_sc_hd__buf_4
XFILLER_232_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23899_ _22969_/X _32491_/Q _23899_/S VGND VGND VPWR VPWR _23900_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28426_ _28426_/A VGND VGND VPWR VPWR _34534_/D sky130_fd_sc_hd__clkbuf_1
X_16440_ _16293_/X _16438_/X _16439_/X _16296_/X VGND VGND VPWR VPWR _16440_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25638_ _25638_/A VGND VGND VPWR VPWR _33246_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28357_ _34502_/Q _24419_/X _28363_/S VGND VGND VPWR VPWR _28358_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16371_ _16293_/X _16367_/X _16370_/X _16296_/X VGND VGND VPWR VPWR _16371_/X sky130_fd_sc_hd__a22o_1
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25569_ _25569_/A VGND VGND VPWR VPWR _33215_/D sky130_fd_sc_hd__clkbuf_1
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_386_CLK clkbuf_6_41__f_CLK/X VGND VGND VPWR VPWR _35826_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_185_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18110_ _35784_/Q _35144_/Q _34504_/Q _33864_/Q _17846_/X _17847_/X VGND VGND VPWR
+ VPWR _18110_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27308_ _27308_/A VGND VGND VPWR VPWR _34005_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19090_ _18941_/X _19086_/X _19089_/X _18944_/X VGND VGND VPWR VPWR _19090_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28288_ _34469_/Q _24317_/X _28300_/S VGND VGND VPWR VPWR _28289_/A sky130_fd_sc_hd__mux2_1
X_18041_ _18037_/X _18040_/X _17834_/X VGND VGND VPWR VPWR _18063_/A sky130_fd_sc_hd__o21ba_2
XFILLER_240_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_138_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _35919_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27239_ _26943_/X _33973_/Q _27239_/S VGND VGND VPWR VPWR _27240_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30250_ _35368_/Q _29132_/X _30256_/S VGND VGND VPWR VPWR _30251_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30181_ _30181_/A VGND VGND VPWR VPWR _35335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19992_ _33276_/Q _36156_/Q _33148_/Q _33084_/Q _19711_/X _19712_/X VGND VGND VPWR
+ VPWR _19992_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18943_ _35742_/Q _35102_/Q _34462_/Q _33822_/Q _18734_/X _18735_/X VGND VGND VPWR
+ VPWR _18943_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33940_ _33940_/CLK _33940_/D VGND VGND VPWR VPWR _33940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_310_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _35320_/CLK sky130_fd_sc_hd__clkbuf_16
X_18874_ _18869_/X _18873_/X _18730_/X _18731_/X VGND VGND VPWR VPWR _18891_/B sky130_fd_sc_hd__o211a_2
XFILLER_234_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17825_ _17825_/A VGND VGND VPWR VPWR _31999_/D sky130_fd_sc_hd__clkbuf_4
X_33871_ _34262_/CLK _33871_/D VGND VGND VPWR VPWR _33871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35610_ _35675_/CLK _35610_/D VGND VGND VPWR VPWR _35610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32822_ _36022_/CLK _32822_/D VGND VGND VPWR VPWR _32822_/Q sky130_fd_sc_hd__dfxtp_1
X_17756_ _17548_/X _17754_/X _17755_/X _17553_/X VGND VGND VPWR VPWR _17756_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16707_ _33248_/Q _36128_/Q _33120_/Q _33056_/Q _16705_/X _16706_/X VGND VGND VPWR
+ VPWR _16707_/X sky130_fd_sc_hd__mux4_1
XFILLER_207_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35541_ _35925_/CLK _35541_/D VGND VGND VPWR VPWR _35541_/Q sky130_fd_sc_hd__dfxtp_1
X_32753_ _36081_/CLK _32753_/D VGND VGND VPWR VPWR _32753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17687_ _33532_/Q _33468_/Q _33404_/Q _33340_/Q _17476_/X _17477_/X VGND VGND VPWR
+ VPWR _17687_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31704_ _31704_/A VGND VGND VPWR VPWR _36056_/D sky130_fd_sc_hd__clkbuf_1
X_19426_ _34028_/Q _33964_/Q _33900_/Q _32236_/Q _19320_/X _19321_/X VGND VGND VPWR
+ VPWR _19426_/X sky130_fd_sc_hd__mux4_1
X_35472_ _35793_/CLK _35472_/D VGND VGND VPWR VPWR _35472_/Q sky130_fd_sc_hd__dfxtp_1
X_16638_ _32990_/Q _32926_/Q _32862_/Q _32798_/Q _16636_/X _16637_/X VGND VGND VPWR
+ VPWR _16638_/X sky130_fd_sc_hd__mux4_1
X_32684_ _36076_/CLK _32684_/D VGND VGND VPWR VPWR _32684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34423_ _35319_/CLK _34423_/D VGND VGND VPWR VPWR _34423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31635_ _36024_/Q input37/X _31649_/S VGND VGND VPWR VPWR _31636_/A sky130_fd_sc_hd__mux2_1
X_19357_ _32746_/Q _32682_/Q _32618_/Q _36074_/Q _19219_/X _19356_/X VGND VGND VPWR
+ VPWR _19357_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_377_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _36013_/CLK sky130_fd_sc_hd__clkbuf_16
X_16569_ _16349_/X _16567_/X _16568_/X _16355_/X VGND VGND VPWR VPWR _16569_/X sky130_fd_sc_hd__a22o_1
X_18308_ _33998_/Q _33934_/Q _33870_/Q _32142_/Q _18305_/X _18307_/X VGND VGND VPWR
+ VPWR _18308_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34354_ _34866_/CLK _34354_/D VGND VGND VPWR VPWR _34354_/Q sky130_fd_sc_hd__dfxtp_1
X_31566_ _31566_/A VGND VGND VPWR VPWR _35991_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19288_ _32488_/Q _32360_/Q _32040_/Q _36008_/Q _19223_/X _19011_/X VGND VGND VPWR
+ VPWR _19288_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33305_ _34267_/CLK _33305_/D VGND VGND VPWR VPWR _33305_/Q sky130_fd_sc_hd__dfxtp_1
X_18239_ _34572_/Q _32460_/Q _34444_/Q _34380_/Q _16063_/X _16065_/X VGND VGND VPWR
+ VPWR _18239_/X sky130_fd_sc_hd__mux4_1
X_30517_ _23217_/X _35494_/Q _30527_/S VGND VGND VPWR VPWR _30518_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_129_CLK clkbuf_6_23__f_CLK/X VGND VGND VPWR VPWR _34259_/CLK sky130_fd_sc_hd__clkbuf_16
X_34285_ _35575_/CLK _34285_/D VGND VGND VPWR VPWR _34285_/Q sky130_fd_sc_hd__dfxtp_1
X_31497_ _31497_/A VGND VGND VPWR VPWR _35958_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33236_ _36116_/CLK _33236_/D VGND VGND VPWR VPWR _33236_/Q sky130_fd_sc_hd__dfxtp_1
X_36024_ _36024_/CLK _36024_/D VGND VGND VPWR VPWR _36024_/Q sky130_fd_sc_hd__dfxtp_1
X_21250_ _21246_/X _21247_/X _21248_/X _21249_/X VGND VGND VPWR VPWR _21250_/X sky130_fd_sc_hd__a22o_1
X_30448_ _30448_/A VGND VGND VPWR VPWR _35461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20201_ _20201_/A VGND VGND VPWR VPWR _20201_/X sky130_fd_sc_hd__buf_4
XFILLER_176_1343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33167_ _35919_/CLK _33167_/D VGND VGND VPWR VPWR _33167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21181_ _21177_/X _21180_/X _21041_/X VGND VGND VPWR VPWR _21191_/C sky130_fd_sc_hd__o21ba_2
X_30379_ _30379_/A VGND VGND VPWR VPWR _35428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20132_ _34048_/Q _33984_/Q _33920_/Q _32256_/Q _20026_/X _20027_/X VGND VGND VPWR
+ VPWR _20132_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32118_ _35811_/CLK _32118_/D VGND VGND VPWR VPWR _32118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33098_ _33548_/CLK _33098_/D VGND VGND VPWR VPWR _33098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20063_ _32766_/Q _32702_/Q _32638_/Q _36094_/Q _19925_/X _20062_/X VGND VGND VPWR
+ VPWR _20063_/X sky130_fd_sc_hd__mux4_1
X_32049_ _36076_/CLK _32049_/D VGND VGND VPWR VPWR _32049_/Q sky130_fd_sc_hd__dfxtp_1
X_24940_ _23003_/X _32950_/Q _24958_/S VGND VGND VPWR VPWR _24941_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_301_CLK clkbuf_6_50__f_CLK/X VGND VGND VPWR VPWR _35834_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24871_ _24871_/A VGND VGND VPWR VPWR _32917_/D sky130_fd_sc_hd__clkbuf_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26610_ _25078_/X _33706_/Q _26612_/S VGND VGND VPWR VPWR _26611_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23822_ _23056_/X _32455_/Q _23826_/S VGND VGND VPWR VPWR _23823_/A sky130_fd_sc_hd__mux2_1
X_35808_ _35808_/CLK _35808_/D VGND VGND VPWR VPWR _35808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27590_ _34138_/Q _24283_/X _27604_/S VGND VGND VPWR VPWR _27591_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_307 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26541_ _25177_/X _33674_/Q _26547_/S VGND VGND VPWR VPWR _26542_/A sky130_fd_sc_hd__mux2_1
XANTENNA_318 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_329 _32141_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20965_ _35734_/Q _35094_/Q _34454_/Q _33814_/Q _20649_/X _20651_/X VGND VGND VPWR
+ VPWR _20965_/X sky130_fd_sc_hd__mux4_1
X_23753_ _22954_/X _32422_/Q _23763_/S VGND VGND VPWR VPWR _23754_/A sky130_fd_sc_hd__mux2_1
X_35739_ _35933_/CLK _35739_/D VGND VGND VPWR VPWR _35739_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22704_ _21749_/A _22702_/X _22703_/X _21752_/A VGND VGND VPWR VPWR _22704_/X sky130_fd_sc_hd__a22o_1
X_29260_ _29260_/A VGND VGND VPWR VPWR _34898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26472_ _25075_/X _33641_/Q _26476_/S VGND VGND VPWR VPWR _26473_/A sky130_fd_sc_hd__mux2_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23684_ _32391_/Q _23327_/X _23688_/S VGND VGND VPWR VPWR _23685_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20896_ _22465_/A VGND VGND VPWR VPWR _20896_/X sky130_fd_sc_hd__buf_4
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28211_ _28211_/A VGND VGND VPWR VPWR _34432_/D sky130_fd_sc_hd__clkbuf_1
X_25423_ _25134_/X _33148_/Q _25429_/S VGND VGND VPWR VPWR _25424_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22635_ _33798_/Q _33734_/Q _33670_/Q _33606_/Q _22502_/X _22503_/X VGND VGND VPWR
+ VPWR _22635_/X sky130_fd_sc_hd__mux4_1
X_29191_ input40/X VGND VGND VPWR VPWR _29191_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_368_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _33262_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_201_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28142_ _26878_/X _34400_/Q _28144_/S VGND VGND VPWR VPWR _28143_/A sky130_fd_sc_hd__mux2_1
X_22566_ _35075_/Q _35011_/Q _34947_/Q _34883_/Q _22462_/X _22463_/X VGND VGND VPWR
+ VPWR _22566_/X sky130_fd_sc_hd__mux4_1
X_25354_ _25032_/X _33115_/Q _25366_/S VGND VGND VPWR VPWR _25355_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1069 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24305_ _32673_/Q _24304_/X _24305_/S VGND VGND VPWR VPWR _24306_/A sky130_fd_sc_hd__mux2_1
X_21517_ _21449_/X _21515_/X _21516_/X _21452_/X VGND VGND VPWR VPWR _21517_/X sky130_fd_sc_hd__a22o_1
XFILLER_210_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28073_ _28073_/A VGND VGND VPWR VPWR _34367_/D sky130_fd_sc_hd__clkbuf_1
X_22497_ _22460_/X _22495_/X _22496_/X _22465_/X VGND VGND VPWR VPWR _22497_/X sky130_fd_sc_hd__a22o_1
X_25285_ _25131_/X _33083_/Q _25293_/S VGND VGND VPWR VPWR _25286_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27024_ _27024_/A VGND VGND VPWR VPWR _33870_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24236_ _23065_/X _32650_/Q _24242_/S VGND VGND VPWR VPWR _24237_/A sky130_fd_sc_hd__mux2_1
X_21448_ _21442_/X _21445_/X _21446_/X _21447_/X VGND VGND VPWR VPWR _21448_/X sky130_fd_sc_hd__a22o_1
XFILLER_181_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24167_ _22963_/X _32617_/Q _24171_/S VGND VGND VPWR VPWR _24168_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21379_ _21302_/X _21377_/X _21378_/X _21308_/X VGND VGND VPWR VPWR _21379_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23118_ _23421_/S VGND VGND VPWR VPWR _23146_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_1_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24098_ _23062_/X _32585_/Q _24098_/S VGND VGND VPWR VPWR _24099_/A sky130_fd_sc_hd__mux2_1
X_28975_ _34795_/Q _24335_/X _28975_/S VGND VGND VPWR VPWR _28976_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23049_ _23049_/A VGND VGND VPWR VPWR _32068_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27926_ _27926_/A VGND VGND VPWR VPWR _34297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27857_ _27857_/A VGND VGND VPWR VPWR _34264_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ _35321_/Q _35257_/Q _35193_/Q _32313_/Q _17359_/X _17360_/X VGND VGND VPWR
+ VPWR _17610_/X sky130_fd_sc_hd__mux4_1
X_26808_ _26808_/A VGND VGND VPWR VPWR _33799_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ _35732_/Q _35092_/Q _34452_/Q _33812_/Q _18349_/X _18351_/X VGND VGND VPWR
+ VPWR _18590_/X sky130_fd_sc_hd__mux4_1
XTAP_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27788_ _34232_/Q _24376_/X _27802_/S VGND VGND VPWR VPWR _27789_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29527_ _35025_/Q _29061_/X _29539_/S VGND VGND VPWR VPWR _29528_/A sky130_fd_sc_hd__mux2_1
XTAP_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ _17502_/X _17539_/X _17540_/X _17505_/X VGND VGND VPWR VPWR _17541_/X sky130_fd_sc_hd__a22o_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26739_ _26739_/A VGND VGND VPWR VPWR _33766_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_830 _23130_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_841 _23322_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_852 _24255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29458_ _29458_/A VGND VGND VPWR VPWR _34992_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17472_ _17472_/A VGND VGND VPWR VPWR _31989_/D sky130_fd_sc_hd__buf_4
XANTENNA_863 _24410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_874 _24979_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19211_ _19211_/A VGND VGND VPWR VPWR _32101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_885 _25171_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16423_ _16416_/X _16421_/X _16422_/X VGND VGND VPWR VPWR _16457_/A sky130_fd_sc_hd__o21ba_1
X_28409_ _28409_/A VGND VGND VPWR VPWR _34526_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_896 _26007_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29389_ _29389_/A VGND VGND VPWR VPWR _34959_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_359_CLK clkbuf_6_41__f_CLK/X VGND VGND VPWR VPWR _36018_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_73_1141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31420_ _23099_/X _35922_/Q _31430_/S VGND VGND VPWR VPWR _31421_/A sky130_fd_sc_hd__mux2_1
X_19142_ _20201_/A VGND VGND VPWR VPWR _19142_/X sky130_fd_sc_hd__clkbuf_4
X_16354_ _33238_/Q _36118_/Q _33110_/Q _33046_/Q _16352_/X _16353_/X VGND VGND VPWR
+ VPWR _16354_/X sky130_fd_sc_hd__mux4_1
XFILLER_242_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31351_ _31351_/A VGND VGND VPWR VPWR _35889_/D sky130_fd_sc_hd__clkbuf_1
X_19073_ _34018_/Q _33954_/Q _33890_/Q _32162_/Q _18967_/X _18968_/X VGND VGND VPWR
+ VPWR _19073_/X sky130_fd_sc_hd__mux4_1
XFILLER_199_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16285_ _32980_/Q _32916_/Q _32852_/Q _32788_/Q _16283_/X _16284_/X VGND VGND VPWR
+ VPWR _16285_/X sky130_fd_sc_hd__mux4_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18024_ _17705_/X _18022_/X _18023_/X _17708_/X VGND VGND VPWR VPWR _18024_/X sky130_fd_sc_hd__a22o_1
X_30302_ _30302_/A VGND VGND VPWR VPWR _35392_/D sky130_fd_sc_hd__clkbuf_1
X_34070_ _34197_/CLK _34070_/D VGND VGND VPWR VPWR _34070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31282_ _31282_/A VGND VGND VPWR VPWR _35856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33021_ _36095_/CLK _33021_/D VGND VGND VPWR VPWR _33021_/Q sky130_fd_sc_hd__dfxtp_1
X_30233_ _35360_/Q _29107_/X _30235_/S VGND VGND VPWR VPWR _30234_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30164_ _30164_/A VGND VGND VPWR VPWR _35327_/D sky130_fd_sc_hd__clkbuf_1
X_19975_ _34811_/Q _34747_/Q _34683_/Q _34619_/Q _19941_/X _19942_/X VGND VGND VPWR
+ VPWR _19975_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18926_ _34270_/Q _34206_/Q _34142_/Q _34078_/Q _18683_/X _18684_/X VGND VGND VPWR
+ VPWR _18926_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30095_ _30095_/A VGND VGND VPWR VPWR _35294_/D sky130_fd_sc_hd__clkbuf_1
X_34972_ _35036_/CLK _34972_/D VGND VGND VPWR VPWR _34972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1240 _25727_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_945 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1251 _26769_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1262 _29247_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33923_ _34057_/CLK _33923_/D VGND VGND VPWR VPWR _33923_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1273 _31408_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18857_ _18857_/A _18857_/B _18857_/C _18857_/D VGND VGND VPWR VPWR _18858_/A sky130_fd_sc_hd__or4_2
XANTENNA_1284 _17843_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1295 _17152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17808_ _17769_/X _17806_/X _17807_/X _17773_/X VGND VGND VPWR VPWR _17808_/X sky130_fd_sc_hd__a22o_1
XFILLER_132_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33854_ _35711_/CLK _33854_/D VGND VGND VPWR VPWR _33854_/Q sky130_fd_sc_hd__dfxtp_1
X_18788_ _18788_/A VGND VGND VPWR VPWR _32089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17739_ _35773_/Q _35133_/Q _34493_/Q _33853_/Q _17493_/X _17494_/X VGND VGND VPWR
+ VPWR _17739_/X sky130_fd_sc_hd__mux4_1
X_32805_ _36069_/CLK _32805_/D VGND VGND VPWR VPWR _32805_/Q sky130_fd_sc_hd__dfxtp_1
X_30997_ _35722_/Q _29237_/X _31003_/S VGND VGND VPWR VPWR _30998_/A sky130_fd_sc_hd__mux2_1
X_33785_ _34298_/CLK _33785_/D VGND VGND VPWR VPWR _33785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35524_ _35973_/CLK _35524_/D VGND VGND VPWR VPWR _35524_/Q sky130_fd_sc_hd__dfxtp_1
X_20750_ _33232_/Q _36112_/Q _33104_/Q _33040_/Q _20620_/X _20621_/X VGND VGND VPWR
+ VPWR _20750_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32736_ _36065_/CLK _32736_/D VGND VGND VPWR VPWR _32736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19409_ _19299_/X _19407_/X _19408_/X _19302_/X VGND VGND VPWR VPWR _19409_/X sky130_fd_sc_hd__a22o_1
X_20681_ _21607_/A VGND VGND VPWR VPWR _20681_/X sky130_fd_sc_hd__buf_4
X_35455_ _36105_/CLK _35455_/D VGND VGND VPWR VPWR _35455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32667_ _35799_/CLK _32667_/D VGND VGND VPWR VPWR _32667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22420_ _34559_/Q _32447_/Q _34431_/Q _34367_/Q _22178_/X _22179_/X VGND VGND VPWR
+ VPWR _22420_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31618_ _36016_/Q input28/X _31628_/S VGND VGND VPWR VPWR _31619_/A sky130_fd_sc_hd__mux2_1
X_34406_ _35942_/CLK _34406_/D VGND VGND VPWR VPWR _34406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35386_ _35386_/CLK _35386_/D VGND VGND VPWR VPWR _35386_/Q sky130_fd_sc_hd__dfxtp_1
X_32598_ _36055_/CLK _32598_/D VGND VGND VPWR VPWR _32598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22351_ _22347_/X _22350_/X _22114_/X VGND VGND VPWR VPWR _22352_/D sky130_fd_sc_hd__o21ba_1
XFILLER_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31549_ _35983_/Q input12/X _31565_/S VGND VGND VPWR VPWR _31550_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34337_ _35039_/CLK _34337_/D VGND VGND VPWR VPWR _34337_/Q sky130_fd_sc_hd__dfxtp_1
X_21302_ _22501_/A VGND VGND VPWR VPWR _21302_/X sky130_fd_sc_hd__clkbuf_4
X_25070_ _25069_/X _32999_/Q _25082_/S VGND VGND VPWR VPWR _25071_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22282_ _22282_/A _22282_/B _22282_/C _22282_/D VGND VGND VPWR VPWR _22283_/A sky130_fd_sc_hd__or4_4
X_34268_ _34777_/CLK _34268_/D VGND VGND VPWR VPWR _34268_/Q sky130_fd_sc_hd__dfxtp_1
X_24021_ _22948_/X _32548_/Q _24035_/S VGND VGND VPWR VPWR _24022_/A sky130_fd_sc_hd__mux2_1
X_33219_ _36034_/CLK _33219_/D VGND VGND VPWR VPWR _33219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36007_ _36007_/CLK _36007_/D VGND VGND VPWR VPWR _36007_/Q sky130_fd_sc_hd__dfxtp_1
X_21233_ _33246_/Q _36126_/Q _33118_/Q _33054_/Q _20952_/X _20953_/X VGND VGND VPWR
+ VPWR _21233_/X sky130_fd_sc_hd__mux4_1
X_34199_ _35667_/CLK _34199_/D VGND VGND VPWR VPWR _34199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21164_ _21096_/X _21162_/X _21163_/X _21099_/X VGND VGND VPWR VPWR _21164_/X sky130_fd_sc_hd__a22o_1
XFILLER_172_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20115_ _20005_/X _20113_/X _20114_/X _20008_/X VGND VGND VPWR VPWR _20115_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28760_ _26993_/X _34693_/Q _28768_/S VGND VGND VPWR VPWR _28761_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25972_ _25134_/X _33404_/Q _25978_/S VGND VGND VPWR VPWR _25973_/A sky130_fd_sc_hd__mux2_1
X_21095_ _21089_/X _21092_/X _21093_/X _21094_/X VGND VGND VPWR VPWR _21095_/X sky130_fd_sc_hd__a22o_1
XFILLER_154_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27711_ _27711_/A VGND VGND VPWR VPWR _34195_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20046_ _35325_/Q _35261_/Q _35197_/Q _32317_/Q _20012_/X _20013_/X VGND VGND VPWR
+ VPWR _20046_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24923_ _22979_/X _32942_/Q _24937_/S VGND VGND VPWR VPWR _24924_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28691_ _26891_/X _34660_/Q _28705_/S VGND VGND VPWR VPWR _28692_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27642_ _34163_/Q _24360_/X _27646_/S VGND VGND VPWR VPWR _27643_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24854_ _30465_/B _31815_/B VGND VGND VPWR VPWR _24987_/S sky130_fd_sc_hd__nand2_8
XFILLER_248_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23805_ _23031_/X _32447_/Q _23805_/S VGND VGND VPWR VPWR _23806_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27573_ _34130_/Q _24258_/X _27583_/S VGND VGND VPWR VPWR _27574_/A sky130_fd_sc_hd__mux2_1
XANTENNA_104 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_115 _32130_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24785_ _24785_/A VGND VGND VPWR VPWR _32876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ _21754_/X _21995_/X _21996_/X _21759_/X VGND VGND VPWR VPWR _21997_/X sky130_fd_sc_hd__a22o_1
XANTENNA_137 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29312_ _29312_/A VGND VGND VPWR VPWR _34923_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26524_ _26524_/A VGND VGND VPWR VPWR _33665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_148 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23736_ _22929_/X _32414_/Q _23742_/S VGND VGND VPWR VPWR _23737_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ _20944_/X _20947_/X _20611_/X VGND VGND VPWR VPWR _20980_/A sky130_fd_sc_hd__o21ba_1
XANTENNA_159 _32133_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29243_ input59/X VGND VGND VPWR VPWR _29243_/X sky130_fd_sc_hd__buf_2
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26455_ _25050_/X _33633_/Q _26455_/S VGND VGND VPWR VPWR _26456_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23667_ _32383_/Q _23300_/X _23667_/S VGND VGND VPWR VPWR _23668_/A sky130_fd_sc_hd__mux2_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20879_ _32724_/Q _32660_/Q _32596_/Q _36052_/Q _20813_/X _22313_/A VGND VGND VPWR
+ VPWR _20879_/X sky130_fd_sc_hd__mux4_1
XFILLER_230_968 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25406_ _25109_/X _33140_/Q _25408_/S VGND VGND VPWR VPWR _25407_/A sky130_fd_sc_hd__mux2_1
X_22618_ _22614_/X _22617_/X _22442_/X _22443_/X VGND VGND VPWR VPWR _22633_/B sky130_fd_sc_hd__o211a_1
X_29174_ _29174_/A VGND VGND VPWR VPWR _34869_/D sky130_fd_sc_hd__clkbuf_1
X_26386_ _25146_/X _33600_/Q _26404_/S VGND VGND VPWR VPWR _26387_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23598_ _32350_/Q _23136_/X _23604_/S VGND VGND VPWR VPWR _23599_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28125_ _28236_/S VGND VGND VPWR VPWR _28144_/S sky130_fd_sc_hd__buf_4
X_25337_ _25007_/X _33107_/Q _25345_/S VGND VGND VPWR VPWR _25338_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22549_ _32515_/Q _32387_/Q _32067_/Q _36035_/Q _22229_/X _22370_/X VGND VGND VPWR
+ VPWR _22549_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16070_ input69/X input70/X VGND VGND VPWR VPWR _17853_/A sky130_fd_sc_hd__or2_4
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28056_ _26950_/X _34359_/Q _28072_/S VGND VGND VPWR VPWR _28057_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25268_ _25106_/X _33075_/Q _25272_/S VGND VGND VPWR VPWR _25269_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27007_ _27007_/A VGND VGND VPWR VPWR _33865_/D sky130_fd_sc_hd__clkbuf_1
X_24219_ _24219_/A VGND VGND VPWR VPWR _32641_/D sky130_fd_sc_hd__clkbuf_1
X_25199_ _25004_/X _33042_/Q _25209_/S VGND VGND VPWR VPWR _25200_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16972_ _34535_/Q _32423_/Q _34407_/Q _34343_/Q _16872_/X _16873_/X VGND VGND VPWR
+ VPWR _16972_/X sky130_fd_sc_hd__mux4_1
X_19760_ _35573_/Q _35509_/Q _35445_/Q _35381_/Q _19550_/X _19551_/X VGND VGND VPWR
+ VPWR _19760_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28958_ _28958_/A VGND VGND VPWR VPWR _34786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18711_ _18707_/X _18710_/X _18400_/X VGND VGND VPWR VPWR _18712_/D sky130_fd_sc_hd__o21ba_1
XTAP_5040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19691_ _19687_/X _19690_/X _19447_/X VGND VGND VPWR VPWR _19699_/C sky130_fd_sc_hd__o21ba_1
X_27909_ _27909_/A VGND VGND VPWR VPWR _34289_/D sky130_fd_sc_hd__clkbuf_1
X_28889_ _26984_/X _34754_/Q _28903_/S VGND VGND VPWR VPWR _28890_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18642_ _33750_/Q _33686_/Q _33622_/Q _33558_/Q _18437_/X _18438_/X VGND VGND VPWR
+ VPWR _18642_/X sky130_fd_sc_hd__mux4_1
XTAP_5084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30920_ _35685_/Q _29123_/X _30932_/S VGND VGND VPWR VPWR _30921_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ _34260_/Q _34196_/Q _34132_/Q _34068_/Q _18305_/X _18307_/X VGND VGND VPWR
+ VPWR _18573_/X sky130_fd_sc_hd__mux4_1
X_30851_ _30851_/A VGND VGND VPWR VPWR _35652_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17524_ _17520_/X _17523_/X _17481_/X VGND VGND VPWR VPWR _17546_/A sky130_fd_sc_hd__o21ba_1
XTAP_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33570_ _33635_/CLK _33570_/D VGND VGND VPWR VPWR _33570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30782_ _30782_/A VGND VGND VPWR VPWR _35619_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_660 _20423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_671 _22460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32521_ _36105_/CLK _32521_/D VGND VGND VPWR VPWR _32521_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_682 _22434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17455_ _17416_/X _17453_/X _17454_/X _17420_/X VGND VGND VPWR VPWR _17455_/X sky130_fd_sc_hd__a22o_1
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_693 _22595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_221_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16406_ _35287_/Q _35223_/Q _35159_/Q _32279_/Q _16300_/X _16301_/X VGND VGND VPWR
+ VPWR _16406_/X sky130_fd_sc_hd__mux4_1
X_32452_ _34947_/CLK _32452_/D VGND VGND VPWR VPWR _32452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35240_ _35304_/CLK _35240_/D VGND VGND VPWR VPWR _35240_/Q sky130_fd_sc_hd__dfxtp_1
X_17386_ _35763_/Q _35123_/Q _34483_/Q _33843_/Q _17140_/X _17141_/X VGND VGND VPWR
+ VPWR _17386_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31403_ _31403_/A VGND VGND VPWR VPWR _35914_/D sky130_fd_sc_hd__clkbuf_1
X_19125_ _19121_/X _19124_/X _19083_/X _19084_/X VGND VGND VPWR VPWR _19140_/B sky130_fd_sc_hd__o211a_1
X_16337_ _35029_/Q _34965_/Q _34901_/Q _34837_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _16337_/X sky130_fd_sc_hd__mux4_1
X_35171_ _35299_/CLK _35171_/D VGND VGND VPWR VPWR _35171_/Q sky130_fd_sc_hd__dfxtp_1
X_32383_ _36031_/CLK _32383_/D VGND VGND VPWR VPWR _32383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34122_ _35273_/CLK _34122_/D VGND VGND VPWR VPWR _34122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19056_ _18946_/X _19054_/X _19055_/X _18949_/X VGND VGND VPWR VPWR _19056_/X sky130_fd_sc_hd__a22o_1
X_31334_ _31334_/A VGND VGND VPWR VPWR _35881_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16268_ _16087_/X _16266_/X _16267_/X _16097_/X VGND VGND VPWR VPWR _16268_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18007_ _17901_/X _18005_/X _18006_/X _17906_/X VGND VGND VPWR VPWR _18007_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34053_ _34053_/CLK _34053_/D VGND VGND VPWR VPWR _34053_/Q sky130_fd_sc_hd__dfxtp_1
X_31265_ _35849_/Q input55/X _31265_/S VGND VGND VPWR VPWR _31266_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16199_ _16074_/X _16197_/X _16198_/X _16084_/X VGND VGND VPWR VPWR _16199_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_60_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _33702_/CLK sky130_fd_sc_hd__clkbuf_16
X_33004_ _33007_/CLK _33004_/D VGND VGND VPWR VPWR _33004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30216_ _30327_/S VGND VGND VPWR VPWR _30235_/S sky130_fd_sc_hd__buf_4
XFILLER_153_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31196_ _35816_/Q input19/X _31202_/S VGND VGND VPWR VPWR _31197_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30147_ _35319_/Q _29179_/X _30163_/S VGND VGND VPWR VPWR _30148_/A sky130_fd_sc_hd__mux2_1
X_19958_ _19954_/X _19957_/X _19781_/X VGND VGND VPWR VPWR _19982_/A sky130_fd_sc_hd__o21ba_1
XFILLER_113_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18909_ _35805_/Q _32180_/Q _35677_/Q _35613_/Q _18907_/X _18908_/X VGND VGND VPWR
+ VPWR _18909_/X sky130_fd_sc_hd__mux4_1
X_34955_ _35788_/CLK _34955_/D VGND VGND VPWR VPWR _34955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30078_ _30078_/A VGND VGND VPWR VPWR _35286_/D sky130_fd_sc_hd__clkbuf_1
X_19889_ _33529_/Q _33465_/Q _33401_/Q _33337_/Q _19776_/X _19777_/X VGND VGND VPWR
+ VPWR _19889_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1070 _17128_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1081 _17194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1092 _17264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21920_ _21599_/X _21918_/X _21919_/X _21602_/X VGND VGND VPWR VPWR _21920_/X sky130_fd_sc_hd__a22o_1
X_33906_ _34286_/CLK _33906_/D VGND VGND VPWR VPWR _33906_/Q sky130_fd_sc_hd__dfxtp_1
X_34886_ _35078_/CLK _34886_/D VGND VGND VPWR VPWR _34886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33837_ _35564_/CLK _33837_/D VGND VGND VPWR VPWR _33837_/Q sky130_fd_sc_hd__dfxtp_1
X_21851_ _22557_/A VGND VGND VPWR VPWR _21851_/X sky130_fd_sc_hd__buf_4
XFILLER_55_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20802_ _20687_/X _20800_/X _20801_/X _20697_/X VGND VGND VPWR VPWR _20802_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24570_ _24570_/A VGND VGND VPWR VPWR _32777_/D sky130_fd_sc_hd__clkbuf_1
X_21782_ _35565_/Q _35501_/Q _35437_/Q _35373_/Q _21497_/X _21498_/X VGND VGND VPWR
+ VPWR _21782_/X sky130_fd_sc_hd__mux4_1
XFILLER_42_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33768_ _34281_/CLK _33768_/D VGND VGND VPWR VPWR _33768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23521_ _23521_/A VGND VGND VPWR VPWR _32314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35507_ _36019_/CLK _35507_/D VGND VGND VPWR VPWR _35507_/Q sky130_fd_sc_hd__dfxtp_1
X_20733_ _20729_/X _20732_/X _20700_/X VGND VGND VPWR VPWR _20734_/D sky130_fd_sc_hd__o21ba_1
XFILLER_180_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32719_ _36048_/CLK _32719_/D VGND VGND VPWR VPWR _32719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33699_ _34276_/CLK _33699_/D VGND VGND VPWR VPWR _33699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26240_ _25131_/X _33531_/Q _26248_/S VGND VGND VPWR VPWR _26241_/A sky130_fd_sc_hd__mux2_1
X_35438_ _35949_/CLK _35438_/D VGND VGND VPWR VPWR _35438_/Q sky130_fd_sc_hd__dfxtp_1
X_23452_ _23452_/A VGND VGND VPWR VPWR _32281_/D sky130_fd_sc_hd__clkbuf_1
X_20664_ _22362_/A VGND VGND VPWR VPWR _22532_/A sky130_fd_sc_hd__buf_12
XFILLER_211_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22403_ _32767_/Q _32703_/Q _32639_/Q _36095_/Q _22225_/X _22362_/X VGND VGND VPWR
+ VPWR _22403_/X sky130_fd_sc_hd__mux4_1
X_23383_ _23383_/A VGND VGND VPWR VPWR _32250_/D sky130_fd_sc_hd__clkbuf_1
X_26171_ _25029_/X _33498_/Q _26185_/S VGND VGND VPWR VPWR _26172_/A sky130_fd_sc_hd__mux2_1
X_20595_ _20595_/A VGND VGND VPWR VPWR _22369_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_167_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35369_ _35819_/CLK _35369_/D VGND VGND VPWR VPWR _35369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25122_ input37/X VGND VGND VPWR VPWR _25122_/X sky130_fd_sc_hd__buf_2
XFILLER_104_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22334_ _32509_/Q _32381_/Q _32061_/Q _36029_/Q _22229_/X _22017_/X VGND VGND VPWR
+ VPWR _22334_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29930_ _35216_/Q _29058_/X _29944_/S VGND VGND VPWR VPWR _29931_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22265_ _22261_/X _22264_/X _22089_/X _22090_/X VGND VGND VPWR VPWR _22282_/B sky130_fd_sc_hd__o211a_1
X_25053_ input13/X VGND VGND VPWR VPWR _25053_/X sky130_fd_sc_hd__buf_2
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_CLK clkbuf_leaf_57_CLK/A VGND VGND VPWR VPWR _34146_/CLK sky130_fd_sc_hd__clkbuf_16
X_24004_ _22923_/X _32540_/Q _24014_/S VGND VGND VPWR VPWR _24005_/A sky130_fd_sc_hd__mux2_1
X_21216_ _34781_/Q _34717_/Q _34653_/Q _34589_/Q _21182_/X _21183_/X VGND VGND VPWR
+ VPWR _21216_/X sky130_fd_sc_hd__mux4_1
X_29861_ _29861_/A VGND VGND VPWR VPWR _35183_/D sky130_fd_sc_hd__clkbuf_1
X_22196_ _32505_/Q _32377_/Q _32057_/Q _36025_/Q _21876_/X _22017_/X VGND VGND VPWR
+ VPWR _22196_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21147_ _33179_/Q _32539_/Q _35931_/Q _35867_/Q _20968_/X _20969_/X VGND VGND VPWR
+ VPWR _21147_/X sky130_fd_sc_hd__mux4_1
X_28812_ _28812_/A VGND VGND VPWR VPWR _34717_/D sky130_fd_sc_hd__clkbuf_1
X_29792_ _29792_/A VGND VGND VPWR VPWR _35150_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28743_ _26968_/X _34685_/Q _28747_/S VGND VGND VPWR VPWR _28744_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21078_ _20893_/X _21076_/X _21077_/X _20896_/X VGND VGND VPWR VPWR _21078_/X sky130_fd_sc_hd__a22o_1
X_25955_ _25109_/X _33396_/Q _25957_/S VGND VGND VPWR VPWR _25956_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20029_ _19855_/X _20025_/X _20028_/X _19858_/X VGND VGND VPWR VPWR _20029_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24906_ _22954_/X _32934_/Q _24916_/S VGND VGND VPWR VPWR _24907_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28674_ _26866_/X _34652_/Q _28684_/S VGND VGND VPWR VPWR _28675_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25886_ _25007_/X _33363_/Q _25894_/S VGND VGND VPWR VPWR _25887_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27625_ _34155_/Q _24335_/X _27625_/S VGND VGND VPWR VPWR _27626_/A sky130_fd_sc_hd__mux2_1
XFILLER_234_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24837_ _24837_/A VGND VGND VPWR VPWR _32901_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27556_ _27556_/A VGND VGND VPWR VPWR _34123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24768_ _24768_/A VGND VGND VPWR VPWR _32868_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26507_ _26507_/A VGND VGND VPWR VPWR _33657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23719_ _22904_/X _32406_/Q _23721_/S VGND VGND VPWR VPWR _23720_/A sky130_fd_sc_hd__mux2_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27487_ _27487_/A VGND VGND VPWR VPWR _34090_/D sky130_fd_sc_hd__clkbuf_1
X_24699_ _23050_/X _32837_/Q _24707_/S VGND VGND VPWR VPWR _24700_/A sky130_fd_sc_hd__mux2_1
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29226_ _34886_/Q _29225_/X _29235_/S VGND VGND VPWR VPWR _29227_/A sky130_fd_sc_hd__mux2_1
X_17240_ _32751_/Q _32687_/Q _32623_/Q _36079_/Q _16919_/X _17056_/X VGND VGND VPWR
+ VPWR _17240_/X sky130_fd_sc_hd__mux4_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26438_ _26438_/A VGND VGND VPWR VPWR _33624_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29157_ input28/X VGND VGND VPWR VPWR _29157_/X sky130_fd_sc_hd__clkbuf_4
X_17171_ _17167_/X _17170_/X _17128_/X VGND VGND VPWR VPWR _17193_/A sky130_fd_sc_hd__o21ba_1
X_26369_ _25122_/X _33592_/Q _26383_/S VGND VGND VPWR VPWR _26370_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16122_ _16044_/X _16120_/X _16121_/X _16054_/X VGND VGND VPWR VPWR _16122_/X sky130_fd_sc_hd__a22o_1
X_28108_ _28108_/A VGND VGND VPWR VPWR _34383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29088_ _29088_/A VGND VGND VPWR VPWR _34841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16053_ _17767_/A VGND VGND VPWR VPWR _17858_/A sky130_fd_sc_hd__buf_12
XFILLER_183_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28039_ _26925_/X _34351_/Q _28051_/S VGND VGND VPWR VPWR _28040_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_42_CLK clkbuf_6_6__f_CLK/X VGND VGND VPWR VPWR _34016_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_142_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1040 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_48__f_CLK clkbuf_5_24_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_48__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_237_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31050_ _31050_/A VGND VGND VPWR VPWR _35746_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30001_ _35250_/Q _29163_/X _30007_/S VGND VGND VPWR VPWR _30002_/A sky130_fd_sc_hd__mux2_1
X_19812_ _20165_/A VGND VGND VPWR VPWR _19812_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_233_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19743_ _20257_/A VGND VGND VPWR VPWR _19743_/X sky130_fd_sc_hd__buf_4
X_16955_ _16702_/X _16953_/X _16954_/X _16708_/X VGND VGND VPWR VPWR _16955_/X sky130_fd_sc_hd__a22o_1
XFILLER_238_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34740_ _35187_/CLK _34740_/D VGND VGND VPWR VPWR _34740_/Q sky130_fd_sc_hd__dfxtp_1
X_31952_ _34973_/CLK _31952_/D VGND VGND VPWR VPWR _31952_/Q sky130_fd_sc_hd__dfxtp_1
X_16886_ _16882_/X _16885_/X _16775_/X VGND VGND VPWR VPWR _16910_/A sky130_fd_sc_hd__o21ba_1
X_19674_ _20147_/A VGND VGND VPWR VPWR _19674_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18625_ _18621_/X _18624_/X _18340_/X _18342_/X VGND VGND VPWR VPWR _18640_/B sky130_fd_sc_hd__o211a_1
X_30903_ _35677_/Q _29098_/X _30911_/S VGND VGND VPWR VPWR _30904_/A sky130_fd_sc_hd__mux2_1
XTAP_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31883_ _31883_/A VGND VGND VPWR VPWR _36141_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34671_ _35242_/CLK _34671_/D VGND VGND VPWR VPWR _34671_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33622_ _34260_/CLK _33622_/D VGND VGND VPWR VPWR _33622_/Q sky130_fd_sc_hd__dfxtp_1
X_30834_ _30834_/A VGND VGND VPWR VPWR _35644_/D sky130_fd_sc_hd__clkbuf_1
X_18556_ _35795_/Q _32169_/Q _35667_/Q _35603_/Q _18554_/X _18555_/X VGND VGND VPWR
+ VPWR _18556_/X sky130_fd_sc_hd__mux4_1
XTAP_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17507_ _17860_/A VGND VGND VPWR VPWR _17507_/X sky130_fd_sc_hd__clkbuf_4
X_33553_ _34259_/CLK _33553_/D VGND VGND VPWR VPWR _33553_/Q sky130_fd_sc_hd__dfxtp_1
X_18487_ _18483_/X _18486_/X _18340_/X _18342_/X VGND VGND VPWR VPWR _18504_/B sky130_fd_sc_hd__o211a_1
X_30765_ _30765_/A VGND VGND VPWR VPWR _35611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_490 _31994_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32504_ _36025_/CLK _32504_/D VGND VGND VPWR VPWR _32504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17438_ _17434_/X _17437_/X _17161_/X VGND VGND VPWR VPWR _17439_/D sky130_fd_sc_hd__o21ba_1
XFILLER_178_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33484_ _33548_/CLK _33484_/D VGND VGND VPWR VPWR _33484_/Q sky130_fd_sc_hd__dfxtp_1
X_30696_ _35579_/Q _29191_/X _30704_/S VGND VGND VPWR VPWR _30697_/A sky130_fd_sc_hd__mux2_1
XANTENNA_15 _32115_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_26 _32116_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_37 _32117_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35223_ _36191_/CLK _35223_/D VGND VGND VPWR VPWR _35223_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_48 _32119_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32435_ _34805_/CLK _32435_/D VGND VGND VPWR VPWR _32435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17369_ _33779_/Q _33715_/Q _33651_/Q _33587_/Q _17196_/X _17197_/X VGND VGND VPWR
+ VPWR _17369_/X sky130_fd_sc_hd__mux4_1
XFILLER_242_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_59 _32126_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19108_ _20167_/A VGND VGND VPWR VPWR _19108_/X sky130_fd_sc_hd__clkbuf_4
X_20380_ _35783_/Q _35143_/Q _34503_/Q _33863_/Q _20146_/X _20147_/X VGND VGND VPWR
+ VPWR _20380_/X sky130_fd_sc_hd__mux4_1
X_35154_ _35282_/CLK _35154_/D VGND VGND VPWR VPWR _35154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32366_ _36015_/CLK _32366_/D VGND VGND VPWR VPWR _32366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34105_ _36152_/CLK _34105_/D VGND VGND VPWR VPWR _34105_/Q sky130_fd_sc_hd__dfxtp_1
X_19039_ _18789_/X _19035_/X _19038_/X _18794_/X VGND VGND VPWR VPWR _19039_/X sky130_fd_sc_hd__a22o_1
X_31317_ _31317_/A VGND VGND VPWR VPWR _35873_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35085_ _35789_/CLK _35085_/D VGND VGND VPWR VPWR _35085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput100 _31969_/Q VGND VGND VPWR VPWR D1[19] sky130_fd_sc_hd__buf_2
X_32297_ _35179_/CLK _32297_/D VGND VGND VPWR VPWR _32297_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput111 _31979_/Q VGND VGND VPWR VPWR D1[29] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_33_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _33692_/CLK sky130_fd_sc_hd__clkbuf_16
Xoutput122 _31989_/Q VGND VGND VPWR VPWR D1[39] sky130_fd_sc_hd__buf_2
X_22050_ _32757_/Q _32693_/Q _32629_/Q _36085_/Q _21872_/X _22009_/X VGND VGND VPWR
+ VPWR _22050_/X sky130_fd_sc_hd__mux4_1
Xoutput133 _31999_/Q VGND VGND VPWR VPWR D1[49] sky130_fd_sc_hd__buf_2
X_31248_ _31248_/A VGND VGND VPWR VPWR _35840_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_1230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34036_ _34228_/CLK _34036_/D VGND VGND VPWR VPWR _34036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput144 _32009_/Q VGND VGND VPWR VPWR D1[59] sky130_fd_sc_hd__buf_2
Xoutput155 _36184_/Q VGND VGND VPWR VPWR D2[10] sky130_fd_sc_hd__buf_2
XFILLER_173_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput166 _36194_/Q VGND VGND VPWR VPWR D2[20] sky130_fd_sc_hd__buf_2
X_21001_ _35543_/Q _35479_/Q _35415_/Q _35351_/Q _20791_/X _20792_/X VGND VGND VPWR
+ VPWR _21001_/X sky130_fd_sc_hd__mux4_1
Xoutput177 _36204_/Q VGND VGND VPWR VPWR D2[30] sky130_fd_sc_hd__buf_2
XFILLER_82_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput188 _36214_/Q VGND VGND VPWR VPWR D2[40] sky130_fd_sc_hd__buf_2
XFILLER_88_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31179_ _35808_/Q input10/X _31181_/S VGND VGND VPWR VPWR _31180_/A sky130_fd_sc_hd__mux2_1
Xoutput199 _36224_/Q VGND VGND VPWR VPWR D2[50] sky130_fd_sc_hd__buf_2
XFILLER_82_1059 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35987_ _35989_/CLK _35987_/D VGND VGND VPWR VPWR _35987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25740_ _25872_/S VGND VGND VPWR VPWR _25759_/S sky130_fd_sc_hd__buf_4
XFILLER_112_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34938_ _35002_/CLK _34938_/D VGND VGND VPWR VPWR _34938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22952_ _22951_/X _32037_/Q _22970_/S VGND VGND VPWR VPWR _22953_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21903_ _34033_/Q _33969_/Q _33905_/Q _32241_/Q _21620_/X _21621_/X VGND VGND VPWR
+ VPWR _21903_/X sky130_fd_sc_hd__mux4_1
X_25671_ _33262_/Q _24345_/X _25685_/S VGND VGND VPWR VPWR _25672_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22883_ input12/X VGND VGND VPWR VPWR _22883_/X sky130_fd_sc_hd__buf_4
XFILLER_56_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34869_ _35061_/CLK _34869_/D VGND VGND VPWR VPWR _34869_/Q sky130_fd_sc_hd__dfxtp_1
X_27410_ _34054_/Q _24419_/X _27416_/S VGND VGND VPWR VPWR _27411_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24622_ _24622_/A VGND VGND VPWR VPWR _32800_/D sky130_fd_sc_hd__clkbuf_1
X_28390_ _28390_/A VGND VGND VPWR VPWR _34517_/D sky130_fd_sc_hd__clkbuf_1
X_21834_ _34287_/Q _34223_/Q _34159_/Q _34095_/Q _21689_/X _21690_/X VGND VGND VPWR
+ VPWR _21834_/X sky130_fd_sc_hd__mux4_1
XFILLER_102_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27341_ _34021_/Q _24317_/X _27353_/S VGND VGND VPWR VPWR _27342_/A sky130_fd_sc_hd__mux2_1
X_24553_ _23038_/X _32769_/Q _24569_/S VGND VGND VPWR VPWR _24554_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21765_ _33773_/Q _33709_/Q _33645_/Q _33581_/Q _21443_/X _21444_/X VGND VGND VPWR
+ VPWR _21765_/X sky130_fd_sc_hd__mux4_1
XFILLER_246_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23504_ _23504_/A VGND VGND VPWR VPWR _32306_/D sky130_fd_sc_hd__clkbuf_1
X_27272_ _27272_/A VGND VGND VPWR VPWR _33988_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20716_ _32463_/Q _32335_/Q _32015_/Q _35983_/Q _20628_/X _22463_/A VGND VGND VPWR
+ VPWR _20716_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24484_ _24484_/A VGND VGND VPWR VPWR _32736_/D sky130_fd_sc_hd__clkbuf_1
X_21696_ _21692_/X _21695_/X _21375_/X VGND VGND VPWR VPWR _21718_/A sky130_fd_sc_hd__o21ba_1
XFILLER_225_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29011_ _34812_/Q _24388_/X _29017_/S VGND VGND VPWR VPWR _29012_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26223_ _25106_/X _33523_/Q _26227_/S VGND VGND VPWR VPWR _26224_/A sky130_fd_sc_hd__mux2_1
X_23435_ _23435_/A VGND VGND VPWR VPWR _32273_/D sky130_fd_sc_hd__clkbuf_1
X_20647_ _35790_/Q _32164_/Q _35662_/Q _35598_/Q _20645_/X _20646_/X VGND VGND VPWR
+ VPWR _20647_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26154_ _25004_/X _33490_/Q _26164_/S VGND VGND VPWR VPWR _26155_/A sky130_fd_sc_hd__mux2_1
X_20578_ input71/X VGND VGND VPWR VPWR _20657_/A sky130_fd_sc_hd__buf_8
XFILLER_221_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23366_ _23366_/A VGND VGND VPWR VPWR _32242_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_2_3_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_25105_ _25105_/A VGND VGND VPWR VPWR _33010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22317_ _35068_/Q _35004_/Q _34940_/Q _34876_/Q _22109_/X _22110_/X VGND VGND VPWR
+ VPWR _22317_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26085_ _26085_/A VGND VGND VPWR VPWR _33457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1076 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23297_ input43/X VGND VGND VPWR VPWR _23297_/X sky130_fd_sc_hd__buf_4
XFILLER_118_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _34205_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_3_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29913_ _29913_/A VGND VGND VPWR VPWR _35208_/D sky130_fd_sc_hd__clkbuf_1
X_25036_ _25035_/X _32988_/Q _25051_/S VGND VGND VPWR VPWR _25037_/A sky130_fd_sc_hd__mux2_1
X_22248_ _22107_/X _22246_/X _22247_/X _22112_/X VGND VGND VPWR VPWR _22248_/X sky130_fd_sc_hd__a22o_1
XFILLER_191_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22179_ _22532_/A VGND VGND VPWR VPWR _22179_/X sky130_fd_sc_hd__buf_4
X_29844_ _29844_/A VGND VGND VPWR VPWR _35175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29775_ _35143_/Q _29228_/X _29779_/S VGND VGND VPWR VPWR _29776_/A sky130_fd_sc_hd__mux2_1
X_26987_ input49/X VGND VGND VPWR VPWR _26987_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_59_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16740_ _33505_/Q _33441_/Q _33377_/Q _33313_/Q _16417_/X _16418_/X VGND VGND VPWR
+ VPWR _16740_/X sky130_fd_sc_hd__mux4_1
XFILLER_87_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28726_ _26943_/X _34677_/Q _28726_/S VGND VGND VPWR VPWR _28727_/A sky130_fd_sc_hd__mux2_1
X_25938_ _26007_/S VGND VGND VPWR VPWR _25957_/S sky130_fd_sc_hd__buf_4
XFILLER_4_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28657_ _26841_/X _34644_/Q _28663_/S VGND VGND VPWR VPWR _28658_/A sky130_fd_sc_hd__mux2_1
X_16671_ _16665_/X _16670_/X _16422_/X VGND VGND VPWR VPWR _16693_/A sky130_fd_sc_hd__o21ba_1
X_25869_ _25869_/A VGND VGND VPWR VPWR _33355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18410_ _33999_/Q _33935_/Q _33871_/Q _32143_/Q _18408_/X _18409_/X VGND VGND VPWR
+ VPWR _18410_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19390_ _20257_/A VGND VGND VPWR VPWR _19390_/X sky130_fd_sc_hd__buf_4
XFILLER_98_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27608_ _27608_/A VGND VGND VPWR VPWR _34146_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28588_ _28588_/A VGND VGND VPWR VPWR _34611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ input82/X VGND VGND VPWR VPWR _20143_/A sky130_fd_sc_hd__buf_12
XFILLER_167_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27539_ _26987_/X _34115_/Q _27551_/S VGND VGND VPWR VPWR _27540_/A sky130_fd_sc_hd__mux2_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18272_ _18268_/X _18271_/X _17867_/A VGND VGND VPWR VPWR _18273_/D sky130_fd_sc_hd__o21ba_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30550_ _30598_/S VGND VGND VPWR VPWR _30569_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_202_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17223_ _35310_/Q _35246_/Q _35182_/Q _32302_/Q _17006_/X _17007_/X VGND VGND VPWR
+ VPWR _17223_/X sky130_fd_sc_hd__mux4_1
X_29209_ _29209_/A VGND VGND VPWR VPWR _34880_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30481_ _23108_/X _35477_/Q _30485_/S VGND VGND VPWR VPWR _30482_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput13 DW[20] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_8
X_32220_ _35843_/CLK _32220_/D VGND VGND VPWR VPWR _32220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput24 DW[30] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__buf_4
X_17154_ _17154_/A VGND VGND VPWR VPWR _17154_/X sky130_fd_sc_hd__clkbuf_4
Xinput35 DW[40] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__buf_4
Xinput46 DW[50] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__buf_6
Xinput57 DW[60] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_16
Xinput68 R1[3] VGND VGND VPWR VPWR input68/X sky130_fd_sc_hd__buf_6
X_16105_ _34255_/Q _34191_/Q _34127_/Q _34063_/Q _16005_/X _16007_/X VGND VGND VPWR
+ VPWR _16105_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32151_ _36220_/CLK _32151_/D VGND VGND VPWR VPWR _32151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput79 R3[2] VGND VGND VPWR VPWR input79/X sky130_fd_sc_hd__clkbuf_4
X_17085_ _17081_/X _17084_/X _16808_/X VGND VGND VPWR VPWR _17086_/D sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_15_CLK clkbuf_6_6__f_CLK/X VGND VGND VPWR VPWR _36063_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31102_ _31102_/A VGND VGND VPWR VPWR _35771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16036_ _32974_/Q _32910_/Q _32846_/Q _32782_/Q _16033_/X _16035_/X VGND VGND VPWR
+ VPWR _16036_/X sky130_fd_sc_hd__mux4_1
X_32082_ _35038_/CLK _32082_/D VGND VGND VPWR VPWR _32082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35910_ _36168_/CLK _35910_/D VGND VGND VPWR VPWR _35910_/Q sky130_fd_sc_hd__dfxtp_1
X_31033_ _31033_/A VGND VGND VPWR VPWR _35738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35841_ _36034_/CLK _35841_/D VGND VGND VPWR VPWR _35841_/Q sky130_fd_sc_hd__dfxtp_1
X_17987_ _35844_/Q _32223_/Q _35716_/Q _35652_/Q _17666_/X _17667_/X VGND VGND VPWR
+ VPWR _17987_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19726_ _35572_/Q _35508_/Q _35444_/Q _35380_/Q _19550_/X _19551_/X VGND VGND VPWR
+ VPWR _19726_/X sky130_fd_sc_hd__mux4_1
X_35772_ _35772_/CLK _35772_/D VGND VGND VPWR VPWR _35772_/Q sky130_fd_sc_hd__dfxtp_1
X_16938_ _35302_/Q _35238_/Q _35174_/Q _32294_/Q _16653_/X _16654_/X VGND VGND VPWR
+ VPWR _16938_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32984_ _36121_/CLK _32984_/D VGND VGND VPWR VPWR _32984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34723_ _35298_/CLK _34723_/D VGND VGND VPWR VPWR _34723_/Q sky130_fd_sc_hd__dfxtp_1
X_31935_ _31935_/A VGND VGND VPWR VPWR _36166_/D sky130_fd_sc_hd__clkbuf_1
X_19657_ _19651_/X _19656_/X _19447_/X VGND VGND VPWR VPWR _19667_/C sky130_fd_sc_hd__o21ba_1
X_16869_ _34788_/Q _34724_/Q _34660_/Q _34596_/Q _16582_/X _16583_/X VGND VGND VPWR
+ VPWR _16869_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18608_ _18608_/A _18608_/B _18608_/C _18608_/D VGND VGND VPWR VPWR _18609_/A sky130_fd_sc_hd__or4_4
XFILLER_203_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34654_ _34781_/CLK _34654_/D VGND VGND VPWR VPWR _34654_/Q sky130_fd_sc_hd__dfxtp_1
X_31866_ _31866_/A VGND VGND VPWR VPWR _36133_/D sky130_fd_sc_hd__clkbuf_1
X_19588_ _20294_/A VGND VGND VPWR VPWR _19588_/X sky130_fd_sc_hd__buf_6
XFILLER_241_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33605_ _34308_/CLK _33605_/D VGND VGND VPWR VPWR _33605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18539_ _18539_/A VGND VGND VPWR VPWR _32082_/D sky130_fd_sc_hd__clkbuf_1
X_30817_ _30817_/A VGND VGND VPWR VPWR _35636_/D sky130_fd_sc_hd__clkbuf_1
X_31797_ _36101_/Q input51/X _31805_/S VGND VGND VPWR VPWR _31798_/A sky130_fd_sc_hd__mux2_1
X_34585_ _36201_/CLK _34585_/D VGND VGND VPWR VPWR _34585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33536_ _34305_/CLK _33536_/D VGND VGND VPWR VPWR _33536_/Q sky130_fd_sc_hd__dfxtp_1
X_21550_ _34023_/Q _33959_/Q _33895_/Q _32204_/Q _21267_/X _21268_/X VGND VGND VPWR
+ VPWR _21550_/X sky130_fd_sc_hd__mux4_1
X_30748_ _30748_/A VGND VGND VPWR VPWR _35603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20501_ _18277_/X _20499_/X _20500_/X _18287_/X VGND VGND VPWR VPWR _20501_/X sky130_fd_sc_hd__a22o_1
XFILLER_194_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21481_ _34277_/Q _34213_/Q _34149_/Q _34085_/Q _21336_/X _21337_/X VGND VGND VPWR
+ VPWR _21481_/X sky130_fd_sc_hd__mux4_1
X_33467_ _33787_/CLK _33467_/D VGND VGND VPWR VPWR _33467_/Q sky130_fd_sc_hd__dfxtp_1
X_30679_ _35571_/Q _29166_/X _30683_/S VGND VGND VPWR VPWR _30680_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35206_ _35339_/CLK _35206_/D VGND VGND VPWR VPWR _35206_/Q sky130_fd_sc_hd__dfxtp_1
X_20432_ _32777_/Q _32713_/Q _32649_/Q _36105_/Q _20278_/X _19173_/A VGND VGND VPWR
+ VPWR _20432_/X sky130_fd_sc_hd__mux4_1
X_23220_ input18/X VGND VGND VPWR VPWR _23220_/X sky130_fd_sc_hd__clkbuf_4
X_32418_ _35298_/CLK _32418_/D VGND VGND VPWR VPWR _32418_/Q sky130_fd_sc_hd__dfxtp_1
X_36186_ _36189_/CLK _36186_/D VGND VGND VPWR VPWR _36186_/Q sky130_fd_sc_hd__dfxtp_1
X_33398_ _34039_/CLK _33398_/D VGND VGND VPWR VPWR _33398_/Q sky130_fd_sc_hd__dfxtp_1
X_35137_ _35843_/CLK _35137_/D VGND VGND VPWR VPWR _35137_/Q sky130_fd_sc_hd__dfxtp_1
X_20363_ _20363_/A _20363_/B _20363_/C _20363_/D VGND VGND VPWR VPWR _20364_/A sky130_fd_sc_hd__or4_1
XFILLER_179_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23151_ _23151_/A VGND VGND VPWR VPWR _32162_/D sky130_fd_sc_hd__clkbuf_1
X_32349_ _36129_/CLK _32349_/D VGND VGND VPWR VPWR _32349_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_7008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22102_ _22455_/A VGND VGND VPWR VPWR _22102_/X sky130_fd_sc_hd__clkbuf_4
XTAP_7019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23082_ _23082_/A VGND VGND VPWR VPWR _27833_/A sky130_fd_sc_hd__buf_8
X_20294_ _20294_/A VGND VGND VPWR VPWR _20294_/X sky130_fd_sc_hd__buf_6
X_35068_ _35517_/CLK _35068_/D VGND VGND VPWR VPWR _35068_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_31__f_CLK clkbuf_5_15_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_31__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XTAP_6318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26910_ _26909_/X _33834_/Q _26913_/S VGND VGND VPWR VPWR _26911_/A sky130_fd_sc_hd__mux2_1
X_22033_ _35316_/Q _35252_/Q _35188_/Q _32308_/Q _21959_/X _21960_/X VGND VGND VPWR
+ VPWR _22033_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34019_ _34149_/CLK _34019_/D VGND VGND VPWR VPWR _34019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_923 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27890_ _27890_/A VGND VGND VPWR VPWR _34280_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26841_ input61/X VGND VGND VPWR VPWR _26841_/X sky130_fd_sc_hd__buf_4
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29560_ _35041_/Q _29110_/X _29560_/S VGND VGND VPWR VPWR _29561_/A sky130_fd_sc_hd__mux2_1
XTAP_4938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26772_ _33782_/Q _24369_/X _26790_/S VGND VGND VPWR VPWR _26773_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23984_ _23984_/A VGND VGND VPWR VPWR _32530_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28511_ _28511_/A VGND VGND VPWR VPWR _34574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25723_ _33287_/Q _24422_/X _25727_/S VGND VGND VPWR VPWR _25724_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29491_ _23303_/X _35008_/Q _29509_/S VGND VGND VPWR VPWR _29492_/A sky130_fd_sc_hd__mux2_1
X_22935_ input10/X VGND VGND VPWR VPWR _22935_/X sky130_fd_sc_hd__buf_4
XFILLER_17_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28442_ _26922_/X _34542_/Q _28456_/S VGND VGND VPWR VPWR _28443_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25654_ _33254_/Q _24320_/X _25664_/S VGND VGND VPWR VPWR _25655_/A sky130_fd_sc_hd__mux2_1
X_22866_ _34829_/Q _34765_/Q _34701_/Q _34637_/Q _22594_/X _22595_/X VGND VGND VPWR
+ VPWR _22866_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24605_ _22910_/X _32792_/Q _24623_/S VGND VGND VPWR VPWR _24606_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28373_ _28778_/B _28373_/B VGND VGND VPWR VPWR _28506_/S sky130_fd_sc_hd__nand2_8
X_21817_ _21594_/X _21815_/X _21816_/X _21597_/X VGND VGND VPWR VPWR _21817_/X sky130_fd_sc_hd__a22o_1
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25585_ _33223_/Q _24422_/X _25589_/S VGND VGND VPWR VPWR _25586_/A sky130_fd_sc_hd__mux2_1
X_22797_ _21754_/A _22795_/X _22796_/X _21759_/A VGND VGND VPWR VPWR _22797_/X sky130_fd_sc_hd__a22o_1
XFILLER_71_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27324_ _34013_/Q _24292_/X _27332_/S VGND VGND VPWR VPWR _27325_/A sky130_fd_sc_hd__mux2_1
XPHY_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24536_ _23013_/X _32761_/Q _24548_/S VGND VGND VPWR VPWR _24537_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21748_ _21743_/X _21746_/X _21747_/X VGND VGND VPWR VPWR _21763_/C sky130_fd_sc_hd__o21ba_1
XPHY_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27255_ _27255_/A VGND VGND VPWR VPWR _33980_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24467_ _22910_/X _32728_/Q _24485_/S VGND VGND VPWR VPWR _24468_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21679_ _34794_/Q _34730_/Q _34666_/Q _34602_/Q _21535_/X _21536_/X VGND VGND VPWR
+ VPWR _21679_/X sky130_fd_sc_hd__mux4_1
X_26206_ _25081_/X _33515_/Q _26206_/S VGND VGND VPWR VPWR _26207_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23418_ _23418_/A VGND VGND VPWR VPWR _32267_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27186_ _27186_/A VGND VGND VPWR VPWR _33947_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24398_ _32703_/Q _24397_/X _24398_/S VGND VGND VPWR VPWR _24399_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26137_ _26137_/A VGND VGND VPWR VPWR _33482_/D sky130_fd_sc_hd__clkbuf_1
X_23349_ _23349_/A VGND VGND VPWR VPWR _32234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26068_ _26068_/A VGND VGND VPWR VPWR _33449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17910_ _34050_/Q _33986_/Q _33922_/Q _32258_/Q _17726_/X _17727_/X VGND VGND VPWR
+ VPWR _17910_/X sky130_fd_sc_hd__mux4_1
X_25019_ input64/X VGND VGND VPWR VPWR _25019_/X sky130_fd_sc_hd__buf_4
XFILLER_238_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18890_ _18886_/X _18889_/X _18755_/X VGND VGND VPWR VPWR _18891_/D sky130_fd_sc_hd__o21ba_1
XTAP_6830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17841_ _17769_/X _17839_/X _17840_/X _17773_/X VGND VGND VPWR VPWR _17841_/X sky130_fd_sc_hd__a22o_1
X_29827_ _29827_/A VGND VGND VPWR VPWR _35167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17772_ _33022_/Q _32958_/Q _32894_/Q _32830_/Q _17695_/X _17696_/X VGND VGND VPWR
+ VPWR _17772_/X sky130_fd_sc_hd__mux4_1
X_29758_ _35135_/Q _29203_/X _29758_/S VGND VGND VPWR VPWR _29759_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19511_ _32494_/Q _32366_/Q _32046_/Q _36014_/Q _19223_/X _19364_/X VGND VGND VPWR
+ VPWR _19511_/X sky130_fd_sc_hd__mux4_1
X_16723_ _33184_/Q _32544_/Q _35936_/Q _35872_/Q _16721_/X _16722_/X VGND VGND VPWR
+ VPWR _16723_/X sky130_fd_sc_hd__mux4_1
X_28709_ _28709_/A VGND VGND VPWR VPWR _34668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29689_ _35102_/Q _29101_/X _29695_/S VGND VGND VPWR VPWR _29690_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19442_ _35756_/Q _35116_/Q _34476_/Q _33836_/Q _19440_/X _19441_/X VGND VGND VPWR
+ VPWR _19442_/X sky130_fd_sc_hd__mux4_1
X_16654_ _17007_/A VGND VGND VPWR VPWR _16654_/X sky130_fd_sc_hd__buf_4
X_31720_ _31720_/A VGND VGND VPWR VPWR _36064_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _34781_/CLK sky130_fd_sc_hd__clkbuf_16
X_31651_ _31678_/S VGND VGND VPWR VPWR _31670_/S sky130_fd_sc_hd__buf_6
X_19373_ _35562_/Q _35498_/Q _35434_/Q _35370_/Q _19197_/X _19198_/X VGND VGND VPWR
+ VPWR _19373_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16585_ _35292_/Q _35228_/Q _35164_/Q _32284_/Q _16300_/X _16301_/X VGND VGND VPWR
+ VPWR _16585_/X sky130_fd_sc_hd__mux4_1
XFILLER_15_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30602_ _35534_/Q _29048_/X _30620_/S VGND VGND VPWR VPWR _30603_/A sky130_fd_sc_hd__mux2_1
X_18324_ _18314_/X _18319_/X _18322_/X _18323_/X VGND VGND VPWR VPWR _18324_/X sky130_fd_sc_hd__a22o_1
X_34370_ _34562_/CLK _34370_/D VGND VGND VPWR VPWR _34370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31582_ _35999_/Q input9/X _31586_/S VGND VGND VPWR VPWR _31583_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18255_ _32525_/Q _32397_/Q _32077_/Q _36045_/Q _17982_/X _17007_/A VGND VGND VPWR
+ VPWR _18255_/X sky130_fd_sc_hd__mux4_1
X_33321_ _35002_/CLK _33321_/D VGND VGND VPWR VPWR _33321_/Q sky130_fd_sc_hd__dfxtp_1
X_30533_ _30533_/A VGND VGND VPWR VPWR _35501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17206_ _17202_/X _17203_/X _17204_/X _17205_/X VGND VGND VPWR VPWR _17206_/X sky130_fd_sc_hd__a22o_1
X_36040_ _36171_/CLK _36040_/D VGND VGND VPWR VPWR _36040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18186_ _34315_/Q _34251_/Q _34187_/Q _34123_/Q _16045_/X _16046_/X VGND VGND VPWR
+ VPWR _18186_/X sky130_fd_sc_hd__mux4_1
X_30464_ _30464_/A VGND VGND VPWR VPWR _35469_/D sky130_fd_sc_hd__clkbuf_1
X_33252_ _36134_/CLK _33252_/D VGND VGND VPWR VPWR _33252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32203_ _36018_/CLK _32203_/D VGND VGND VPWR VPWR _32203_/Q sky130_fd_sc_hd__dfxtp_1
X_17137_ _17843_/A VGND VGND VPWR VPWR _17137_/X sky130_fd_sc_hd__clkbuf_4
X_33183_ _35935_/CLK _33183_/D VGND VGND VPWR VPWR _33183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30395_ _23237_/X _35436_/Q _30413_/S VGND VGND VPWR VPWR _30396_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32134_ _35750_/CLK _32134_/D VGND VGND VPWR VPWR _32134_/Q sky130_fd_sc_hd__dfxtp_1
X_17068_ _17063_/X _17065_/X _17066_/X _17067_/X VGND VGND VPWR VPWR _17068_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16019_ _32718_/Q _32654_/Q _32590_/Q _36046_/Q _17862_/A _17713_/A VGND VGND VPWR
+ VPWR _16019_/X sky130_fd_sc_hd__mux4_1
X_32065_ _36032_/CLK _32065_/D VGND VGND VPWR VPWR _32065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31016_ _31016_/A VGND VGND VPWR VPWR _35730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35824_ _35951_/CLK _35824_/D VGND VGND VPWR VPWR _35824_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19709_ _20062_/A VGND VGND VPWR VPWR _19709_/X sky130_fd_sc_hd__clkbuf_4
X_35755_ _35945_/CLK _35755_/D VGND VGND VPWR VPWR _35755_/Q sky130_fd_sc_hd__dfxtp_1
X_32967_ _32967_/CLK _32967_/D VGND VGND VPWR VPWR _32967_/Q sky130_fd_sc_hd__dfxtp_1
X_20981_ _20981_/A VGND VGND VPWR VPWR _36182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22720_ _35080_/Q _35016_/Q _34952_/Q _34888_/Q _22462_/X _22463_/X VGND VGND VPWR
+ VPWR _22720_/X sky130_fd_sc_hd__mux4_1
X_34706_ _34706_/CLK _34706_/D VGND VGND VPWR VPWR _34706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31918_ _31918_/A VGND VGND VPWR VPWR _36158_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35686_ _35750_/CLK _35686_/D VGND VGND VPWR VPWR _35686_/Q sky130_fd_sc_hd__dfxtp_1
X_32898_ _32965_/CLK _32898_/D VGND VGND VPWR VPWR _32898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34637_ _35341_/CLK _34637_/D VGND VGND VPWR VPWR _34637_/Q sky130_fd_sc_hd__dfxtp_1
X_22651_ _20577_/X _22649_/X _22650_/X _20587_/X VGND VGND VPWR VPWR _22651_/X sky130_fd_sc_hd__a22o_1
XFILLER_213_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31849_ _31849_/A VGND VGND VPWR VPWR _36125_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21602_ _22465_/A VGND VGND VPWR VPWR _21602_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_34_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25370_ _25370_/A VGND VGND VPWR VPWR _33122_/D sky130_fd_sc_hd__clkbuf_1
X_34568_ _35080_/CLK _34568_/D VGND VGND VPWR VPWR _34568_/Q sky130_fd_sc_hd__dfxtp_1
X_22582_ _22582_/A VGND VGND VPWR VPWR _22582_/X sky130_fd_sc_hd__buf_6
XFILLER_146_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24321_ _32678_/Q _24320_/X _24336_/S VGND VGND VPWR VPWR _24322_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21533_ _21246_/X _21531_/X _21532_/X _21249_/X VGND VGND VPWR VPWR _21533_/X sky130_fd_sc_hd__a22o_1
X_33519_ _33520_/CLK _33519_/D VGND VGND VPWR VPWR _33519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34499_ _35778_/CLK _34499_/D VGND VGND VPWR VPWR _34499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27040_ _27040_/A VGND VGND VPWR VPWR _33878_/D sky130_fd_sc_hd__clkbuf_1
X_24252_ input23/X VGND VGND VPWR VPWR _24252_/X sky130_fd_sc_hd__buf_6
X_21464_ _21241_/X _21462_/X _21463_/X _21244_/X VGND VGND VPWR VPWR _21464_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23203_ _23203_/A VGND VGND VPWR VPWR _32183_/D sky130_fd_sc_hd__clkbuf_1
X_20415_ _20411_/X _20414_/X _20153_/X VGND VGND VPWR VPWR _20423_/C sky130_fd_sc_hd__o21ba_1
XFILLER_175_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36169_ _36169_/CLK _36169_/D VGND VGND VPWR VPWR _36169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21395_ _21390_/X _21393_/X _21394_/X VGND VGND VPWR VPWR _21410_/C sky130_fd_sc_hd__o21ba_1
X_24183_ _24183_/A VGND VGND VPWR VPWR _32624_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23134_ _32157_/Q _23133_/X _23146_/S VGND VGND VPWR VPWR _23135_/A sky130_fd_sc_hd__mux2_1
X_20346_ _33030_/Q _32966_/Q _32902_/Q _32838_/Q _18280_/X _18283_/X VGND VGND VPWR
+ VPWR _20346_/X sky130_fd_sc_hd__mux4_1
X_28991_ _28991_/A VGND VGND VPWR VPWR _34802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23065_ input57/X VGND VGND VPWR VPWR _23065_/X sky130_fd_sc_hd__buf_2
X_20277_ _20273_/X _20276_/X _20134_/X VGND VGND VPWR VPWR _20303_/A sky130_fd_sc_hd__o21ba_1
XTAP_6115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27942_ _34305_/Q _24404_/X _27958_/S VGND VGND VPWR VPWR _27943_/A sky130_fd_sc_hd__mux2_1
XTAP_6126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22016_ _22508_/A VGND VGND VPWR VPWR _22016_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27873_ _27873_/A VGND VGND VPWR VPWR _34272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29612_ _29612_/A VGND VGND VPWR VPWR _35065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26824_ _26821_/X _33806_/Q _26851_/S VGND VGND VPWR VPWR _26825_/A sky130_fd_sc_hd__mux2_1
XTAP_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29543_ _29543_/A VGND VGND VPWR VPWR _35032_/D sky130_fd_sc_hd__clkbuf_1
X_26755_ _33774_/Q _24345_/X _26769_/S VGND VGND VPWR VPWR _26756_/A sky130_fd_sc_hd__mux2_1
X_23967_ _23967_/A VGND VGND VPWR VPWR _32523_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25706_ _33279_/Q _24397_/X _25706_/S VGND VGND VPWR VPWR _25707_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22918_ _22917_/X _32026_/Q _22939_/S VGND VGND VPWR VPWR _22919_/A sky130_fd_sc_hd__mux2_1
X_26686_ _26686_/A VGND VGND VPWR VPWR _26819_/S sky130_fd_sc_hd__buf_12
X_29474_ _23277_/X _35000_/Q _29488_/S VGND VGND VPWR VPWR _29475_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23898_ _23898_/A VGND VGND VPWR VPWR _32490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28425_ _26897_/X _34534_/Q _28435_/S VGND VGND VPWR VPWR _28426_/A sky130_fd_sc_hd__mux2_1
X_25637_ _33246_/Q _24295_/X _25643_/S VGND VGND VPWR VPWR _25638_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22849_ _34061_/Q _33997_/Q _33933_/Q _32269_/Q _20658_/X _20660_/X VGND VGND VPWR
+ VPWR _22849_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28356_ _28356_/A VGND VGND VPWR VPWR _34501_/D sky130_fd_sc_hd__clkbuf_1
X_16370_ _33174_/Q _32534_/Q _35926_/Q _35862_/Q _16368_/X _16369_/X VGND VGND VPWR
+ VPWR _16370_/X sky130_fd_sc_hd__mux4_1
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25568_ _33215_/Q _24397_/X _25568_/S VGND VGND VPWR VPWR _25569_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27307_ _34005_/Q _24267_/X _27311_/S VGND VGND VPWR VPWR _27308_/A sky130_fd_sc_hd__mux2_1
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24519_ _22988_/X _32753_/Q _24527_/S VGND VGND VPWR VPWR _24520_/A sky130_fd_sc_hd__mux2_1
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28287_ _28287_/A VGND VGND VPWR VPWR _34468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25499_ _33182_/Q _24295_/X _25505_/S VGND VGND VPWR VPWR _25500_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18040_ _17908_/X _18038_/X _18039_/X _17911_/X VGND VGND VPWR VPWR _18040_/X sky130_fd_sc_hd__a22o_1
X_27238_ _27238_/A VGND VGND VPWR VPWR _33972_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27169_ _27169_/A VGND VGND VPWR VPWR _33939_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30180_ _35335_/Q _29228_/X _30184_/S VGND VGND VPWR VPWR _30181_/A sky130_fd_sc_hd__mux2_1
X_19991_ _32764_/Q _32700_/Q _32636_/Q _36092_/Q _19925_/X _19709_/X VGND VGND VPWR
+ VPWR _19991_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18942_ _35806_/Q _32181_/Q _35678_/Q _35614_/Q _18907_/X _18908_/X VGND VGND VPWR
+ VPWR _18942_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18873_ _18657_/X _18871_/X _18872_/X _18661_/X VGND VGND VPWR VPWR _18873_/X sky130_fd_sc_hd__a22o_1
XTAP_6660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17824_ _17824_/A _17824_/B _17824_/C _17824_/D VGND VGND VPWR VPWR _17825_/A sky130_fd_sc_hd__or4_4
X_33870_ _34262_/CLK _33870_/D VGND VGND VPWR VPWR _33870_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32821_ _36021_/CLK _32821_/D VGND VGND VPWR VPWR _32821_/Q sky130_fd_sc_hd__dfxtp_1
X_17755_ _34302_/Q _34238_/Q _34174_/Q _34110_/Q _17442_/X _17443_/X VGND VGND VPWR
+ VPWR _17755_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35540_ _35797_/CLK _35540_/D VGND VGND VPWR VPWR _35540_/Q sky130_fd_sc_hd__dfxtp_1
X_16706_ _17903_/A VGND VGND VPWR VPWR _16706_/X sky130_fd_sc_hd__clkbuf_4
X_32752_ _33009_/CLK _32752_/D VGND VGND VPWR VPWR _32752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17686_ _17548_/X _17684_/X _17685_/X _17553_/X VGND VGND VPWR VPWR _17686_/X sky130_fd_sc_hd__a22o_1
XFILLER_223_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31703_ _36056_/Q input2/X _31721_/S VGND VGND VPWR VPWR _31704_/A sky130_fd_sc_hd__mux2_1
X_19425_ _33516_/Q _33452_/Q _33388_/Q _33324_/Q _19423_/X _19424_/X VGND VGND VPWR
+ VPWR _19425_/X sky130_fd_sc_hd__mux4_2
XFILLER_90_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35471_ _35791_/CLK _35471_/D VGND VGND VPWR VPWR _35471_/Q sky130_fd_sc_hd__dfxtp_1
X_16637_ _17830_/A VGND VGND VPWR VPWR _16637_/X sky130_fd_sc_hd__clkbuf_4
X_32683_ _36137_/CLK _32683_/D VGND VGND VPWR VPWR _32683_/Q sky130_fd_sc_hd__dfxtp_1
X_34422_ _35319_/CLK _34422_/D VGND VGND VPWR VPWR _34422_/Q sky130_fd_sc_hd__dfxtp_1
X_19356_ _20062_/A VGND VGND VPWR VPWR _19356_/X sky130_fd_sc_hd__buf_6
X_31634_ _31634_/A VGND VGND VPWR VPWR _36023_/D sky130_fd_sc_hd__clkbuf_1
X_16568_ _33244_/Q _36124_/Q _33116_/Q _33052_/Q _16352_/X _16353_/X VGND VGND VPWR
+ VPWR _16568_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18307_ _20257_/A VGND VGND VPWR VPWR _18307_/X sky130_fd_sc_hd__buf_4
XFILLER_52_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34353_ _34866_/CLK _34353_/D VGND VGND VPWR VPWR _34353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31565_ _35991_/Q input64/X _31565_/S VGND VGND VPWR VPWR _31566_/A sky130_fd_sc_hd__mux2_1
X_16499_ _17865_/A VGND VGND VPWR VPWR _16499_/X sky130_fd_sc_hd__buf_4
X_19287_ _19002_/X _19285_/X _19286_/X _19008_/X VGND VGND VPWR VPWR _19287_/X sky130_fd_sc_hd__a22o_1
XFILLER_206_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33304_ _36194_/CLK _33304_/D VGND VGND VPWR VPWR _33304_/Q sky130_fd_sc_hd__dfxtp_1
X_18238_ _16044_/X _18236_/X _18237_/X _16054_/X VGND VGND VPWR VPWR _18238_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30516_ _30516_/A VGND VGND VPWR VPWR _35493_/D sky130_fd_sc_hd__clkbuf_1
X_34284_ _35252_/CLK _34284_/D VGND VGND VPWR VPWR _34284_/Q sky130_fd_sc_hd__dfxtp_1
X_31496_ _23270_/X _35958_/Q _31514_/S VGND VGND VPWR VPWR _31497_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36023_ _36023_/CLK _36023_/D VGND VGND VPWR VPWR _36023_/Q sky130_fd_sc_hd__dfxtp_1
X_30447_ _23319_/X _35461_/Q _30455_/S VGND VGND VPWR VPWR _30448_/A sky130_fd_sc_hd__mux2_1
X_33235_ _36115_/CLK _33235_/D VGND VGND VPWR VPWR _33235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18169_ _35850_/Q _32230_/Q _35722_/Q _35658_/Q _15989_/X _15991_/X VGND VGND VPWR
+ VPWR _18169_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20200_ _20200_/A VGND VGND VPWR VPWR _32129_/D sky130_fd_sc_hd__buf_4
XFILLER_116_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21180_ _20893_/X _21178_/X _21179_/X _20896_/X VGND VGND VPWR VPWR _21180_/X sky130_fd_sc_hd__a22o_1
XFILLER_239_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33166_ _35919_/CLK _33166_/D VGND VGND VPWR VPWR _33166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30378_ _23175_/X _35428_/Q _30392_/S VGND VGND VPWR VPWR _30379_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_1298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20131_ _33536_/Q _33472_/Q _33408_/Q _33344_/Q _20129_/X _20130_/X VGND VGND VPWR
+ VPWR _20131_/X sky130_fd_sc_hd__mux4_1
X_32117_ _35811_/CLK _32117_/D VGND VGND VPWR VPWR _32117_/Q sky130_fd_sc_hd__dfxtp_1
X_33097_ _36169_/CLK _33097_/D VGND VGND VPWR VPWR _33097_/Q sky130_fd_sc_hd__dfxtp_1
X_20062_ _20062_/A VGND VGND VPWR VPWR _20062_/X sky130_fd_sc_hd__clkbuf_4
X_32048_ _36077_/CLK _32048_/D VGND VGND VPWR VPWR _32048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24870_ _22901_/X _32917_/Q _24874_/S VGND VGND VPWR VPWR _24871_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1096 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23821_ _23821_/A VGND VGND VPWR VPWR _32454_/D sky130_fd_sc_hd__clkbuf_1
X_35807_ _35807_/CLK _35807_/D VGND VGND VPWR VPWR _35807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33999_ _34262_/CLK _33999_/D VGND VGND VPWR VPWR _33999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26540_ _26540_/A VGND VGND VPWR VPWR _33673_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_308 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23752_ _23752_/A VGND VGND VPWR VPWR _32421_/D sky130_fd_sc_hd__clkbuf_1
X_35738_ _35738_/CLK _35738_/D VGND VGND VPWR VPWR _35738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20964_ _35798_/Q _32173_/Q _35670_/Q _35606_/Q _20854_/X _20855_/X VGND VGND VPWR
+ VPWR _20964_/X sky130_fd_sc_hd__mux4_1
XANTENNA_319 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22703_ _33288_/Q _36168_/Q _33160_/Q _33096_/Q _20628_/X _21757_/A VGND VGND VPWR
+ VPWR _22703_/X sky130_fd_sc_hd__mux4_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26471_ _26471_/A VGND VGND VPWR VPWR _33640_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23683_ _23683_/A VGND VGND VPWR VPWR _32390_/D sky130_fd_sc_hd__clkbuf_1
X_35669_ _35669_/CLK _35669_/D VGND VGND VPWR VPWR _35669_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20895_ _33172_/Q _32532_/Q _35924_/Q _35860_/Q _20663_/X _20665_/X VGND VGND VPWR
+ VPWR _20895_/X sky130_fd_sc_hd__mux4_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28210_ _26977_/X _34432_/Q _28228_/S VGND VGND VPWR VPWR _28211_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25422_ _25422_/A VGND VGND VPWR VPWR _33147_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22634_ _22634_/A VGND VGND VPWR VPWR _36229_/D sky130_fd_sc_hd__clkbuf_1
X_29190_ _29190_/A VGND VGND VPWR VPWR _34874_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28141_ _28141_/A VGND VGND VPWR VPWR _34399_/D sky130_fd_sc_hd__clkbuf_1
X_25353_ _25353_/A VGND VGND VPWR VPWR _33114_/D sky130_fd_sc_hd__clkbuf_1
X_22565_ _34563_/Q _32451_/Q _34435_/Q _34371_/Q _22531_/X _22532_/X VGND VGND VPWR
+ VPWR _22565_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1086 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_946 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24304_ input11/X VGND VGND VPWR VPWR _24304_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_70_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28072_ _26974_/X _34367_/Q _28072_/S VGND VGND VPWR VPWR _28073_/A sky130_fd_sc_hd__mux2_1
X_21516_ _34022_/Q _33958_/Q _33894_/Q _32193_/Q _21267_/X _21268_/X VGND VGND VPWR
+ VPWR _21516_/X sky130_fd_sc_hd__mux4_1
X_25284_ _25284_/A VGND VGND VPWR VPWR _33082_/D sky130_fd_sc_hd__clkbuf_1
X_22496_ _35073_/Q _35009_/Q _34945_/Q _34881_/Q _22462_/X _22463_/X VGND VGND VPWR
+ VPWR _22496_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27023_ _26821_/X _33870_/Q _27041_/S VGND VGND VPWR VPWR _27024_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24235_ _24235_/A VGND VGND VPWR VPWR _32649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21447_ _22506_/A VGND VGND VPWR VPWR _21447_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_120_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24166_ _24166_/A VGND VGND VPWR VPWR _32616_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21378_ _33250_/Q _36130_/Q _33122_/Q _33058_/Q _21305_/X _21306_/X VGND VGND VPWR
+ VPWR _21378_/X sky130_fd_sc_hd__mux4_1
XFILLER_218_1127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23117_ input2/X VGND VGND VPWR VPWR _23117_/X sky130_fd_sc_hd__clkbuf_8
X_20329_ _34565_/Q _32453_/Q _34437_/Q _34373_/Q _20231_/X _20232_/X VGND VGND VPWR
+ VPWR _20329_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24097_ _24097_/A VGND VGND VPWR VPWR _32584_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28974_ _28974_/A VGND VGND VPWR VPWR _34794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23048_ _23047_/X _32068_/Q _23063_/S VGND VGND VPWR VPWR _23049_/A sky130_fd_sc_hd__mux2_1
XTAP_5200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27925_ _34297_/Q _24379_/X _27937_/S VGND VGND VPWR VPWR _27926_/A sky130_fd_sc_hd__mux2_1
XTAP_5211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27856_ _34264_/Q _24276_/X _27874_/S VGND VGND VPWR VPWR _27857_/A sky130_fd_sc_hd__mux2_1
XTAP_5266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26807_ _33799_/Q _24422_/X _26811_/S VGND VGND VPWR VPWR _26808_/A sky130_fd_sc_hd__mux2_1
XTAP_5299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24999_ _24998_/X _32976_/Q _25020_/S VGND VGND VPWR VPWR _25000_/A sky130_fd_sc_hd__mux2_1
XTAP_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27787_ _27787_/A VGND VGND VPWR VPWR _34231_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29526_ _29526_/A VGND VGND VPWR VPWR _35024_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17540_ _35319_/Q _35255_/Q _35191_/Q _32311_/Q _17359_/X _17360_/X VGND VGND VPWR
+ VPWR _17540_/X sky130_fd_sc_hd__mux4_1
XTAP_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26738_ _33766_/Q _24320_/X _26748_/S VGND VGND VPWR VPWR _26739_/A sky130_fd_sc_hd__mux2_1
XTAP_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_820 _23003_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_831 _23133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_842 _23330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17471_ _17471_/A _17471_/B _17471_/C _17471_/D VGND VGND VPWR VPWR _17472_/A sky130_fd_sc_hd__or4_1
X_26669_ _25165_/X _33734_/Q _26675_/S VGND VGND VPWR VPWR _26670_/A sky130_fd_sc_hd__mux2_1
X_29457_ _23250_/X _34992_/Q _29467_/S VGND VGND VPWR VPWR _29458_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_853 _24264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_864 _24413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_875 _24979_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19210_ _19210_/A _19210_/B _19210_/C _19210_/D VGND VGND VPWR VPWR _19211_/A sky130_fd_sc_hd__or4_4
XFILLER_220_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_886 _25171_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16422_ _17834_/A VGND VGND VPWR VPWR _16422_/X sky130_fd_sc_hd__clkbuf_4
X_28408_ _26872_/X _34526_/Q _28414_/S VGND VGND VPWR VPWR _28409_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29388_ _23090_/X _34959_/Q _29404_/S VGND VGND VPWR VPWR _29389_/A sky130_fd_sc_hd__mux2_1
XANTENNA_897 _26007_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16353_ _17903_/A VGND VGND VPWR VPWR _16353_/X sky130_fd_sc_hd__clkbuf_4
X_19141_ _19141_/A VGND VGND VPWR VPWR _32099_/D sky130_fd_sc_hd__clkbuf_1
X_28339_ _28339_/A VGND VGND VPWR VPWR _34493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19072_ _33506_/Q _33442_/Q _33378_/Q _33314_/Q _19070_/X _19071_/X VGND VGND VPWR
+ VPWR _19072_/X sky130_fd_sc_hd__mux4_1
X_31350_ _35889_/Q input29/X _31358_/S VGND VGND VPWR VPWR _31351_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16284_ _17830_/A VGND VGND VPWR VPWR _16284_/X sky130_fd_sc_hd__buf_4
XFILLER_125_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30301_ _35392_/Q _29206_/X _30319_/S VGND VGND VPWR VPWR _30302_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18023_ _33221_/Q _32581_/Q _35973_/Q _35909_/Q _17780_/X _17781_/X VGND VGND VPWR
+ VPWR _18023_/X sky130_fd_sc_hd__mux4_1
X_31281_ _35856_/Q input23/X _31295_/S VGND VGND VPWR VPWR _31282_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33020_ _36095_/CLK _33020_/D VGND VGND VPWR VPWR _33020_/Q sky130_fd_sc_hd__dfxtp_1
X_30232_ _30232_/A VGND VGND VPWR VPWR _35359_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30163_ _35327_/Q _29203_/X _30163_/S VGND VGND VPWR VPWR _30164_/A sky130_fd_sc_hd__mux2_1
X_19974_ _19970_/X _19973_/X _19800_/X VGND VGND VPWR VPWR _19982_/C sky130_fd_sc_hd__o21ba_1
XFILLER_113_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18925_ _33758_/Q _33694_/Q _33630_/Q _33566_/Q _18790_/X _18791_/X VGND VGND VPWR
+ VPWR _18925_/X sky130_fd_sc_hd__mux4_1
X_30094_ _35294_/Q _29101_/X _30100_/S VGND VGND VPWR VPWR _30095_/A sky130_fd_sc_hd__mux2_1
X_34971_ _35166_/CLK _34971_/D VGND VGND VPWR VPWR _34971_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1230 _24416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1241 _25872_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_295_CLK clkbuf_6_51__f_CLK/X VGND VGND VPWR VPWR _35837_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_1252 _26853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33922_ _33922_/CLK _33922_/D VGND VGND VPWR VPWR _33922_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1263 _29098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18856_ _18852_/X _18855_/X _18755_/X VGND VGND VPWR VPWR _18857_/D sky130_fd_sc_hd__o21ba_1
XFILLER_67_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1274 _31543_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1285 _17843_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1296 _17154_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17807_ _33023_/Q _32959_/Q _32895_/Q _32831_/Q _17695_/X _17696_/X VGND VGND VPWR
+ VPWR _17807_/X sky130_fd_sc_hd__mux4_1
X_33853_ _35711_/CLK _33853_/D VGND VGND VPWR VPWR _33853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18787_ _18787_/A _18787_/B _18787_/C _18787_/D VGND VGND VPWR VPWR _18788_/A sky130_fd_sc_hd__or4_2
X_15999_ _17796_/A VGND VGND VPWR VPWR _15999_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_94_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32804_ _36067_/CLK _32804_/D VGND VGND VPWR VPWR _32804_/Q sky130_fd_sc_hd__dfxtp_1
X_17738_ _35837_/Q _32216_/Q _35709_/Q _35645_/Q _17666_/X _17667_/X VGND VGND VPWR
+ VPWR _17738_/X sky130_fd_sc_hd__mux4_1
X_33784_ _34296_/CLK _33784_/D VGND VGND VPWR VPWR _33784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30996_ _30996_/A VGND VGND VPWR VPWR _35721_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35523_ _35909_/CLK _35523_/D VGND VGND VPWR VPWR _35523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32735_ _35801_/CLK _32735_/D VGND VGND VPWR VPWR _32735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17669_ _35771_/Q _35131_/Q _34491_/Q _33851_/Q _17493_/X _17494_/X VGND VGND VPWR
+ VPWR _17669_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19408_ _33195_/Q _32555_/Q _35947_/Q _35883_/Q _19374_/X _19375_/X VGND VGND VPWR
+ VPWR _19408_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35454_ _35966_/CLK _35454_/D VGND VGND VPWR VPWR _35454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20680_ _22362_/A VGND VGND VPWR VPWR _21607_/A sky130_fd_sc_hd__buf_12
X_32666_ _32666_/CLK _32666_/D VGND VGND VPWR VPWR _32666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34405_ _35942_/CLK _34405_/D VGND VGND VPWR VPWR _34405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31617_ _31617_/A VGND VGND VPWR VPWR _36015_/D sky130_fd_sc_hd__clkbuf_1
X_19339_ _34793_/Q _34729_/Q _34665_/Q _34601_/Q _19235_/X _19236_/X VGND VGND VPWR
+ VPWR _19339_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35385_ _35577_/CLK _35385_/D VGND VGND VPWR VPWR _35385_/Q sky130_fd_sc_hd__dfxtp_1
X_32597_ _36116_/CLK _32597_/D VGND VGND VPWR VPWR _32597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22350_ _22107_/X _22348_/X _22349_/X _22112_/X VGND VGND VPWR VPWR _22350_/X sky130_fd_sc_hd__a22o_1
X_34336_ _35039_/CLK _34336_/D VGND VGND VPWR VPWR _34336_/Q sky130_fd_sc_hd__dfxtp_1
X_31548_ _31548_/A VGND VGND VPWR VPWR _35982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21301_ _21297_/X _21300_/X _21022_/X VGND VGND VPWR VPWR _21333_/A sky130_fd_sc_hd__o21ba_1
XFILLER_163_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22281_ _22277_/X _22280_/X _22114_/X VGND VGND VPWR VPWR _22282_/D sky130_fd_sc_hd__o21ba_1
X_34267_ _34267_/CLK _34267_/D VGND VGND VPWR VPWR _34267_/Q sky130_fd_sc_hd__dfxtp_1
X_31479_ _23244_/X _35950_/Q _31493_/S VGND VGND VPWR VPWR _31480_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24020_ _24020_/A VGND VGND VPWR VPWR _32547_/D sky130_fd_sc_hd__clkbuf_1
X_36006_ _36007_/CLK _36006_/D VGND VGND VPWR VPWR _36006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33218_ _35906_/CLK _33218_/D VGND VGND VPWR VPWR _33218_/Q sky130_fd_sc_hd__dfxtp_1
X_21232_ _32734_/Q _32670_/Q _32606_/Q _36062_/Q _21166_/X _20950_/X VGND VGND VPWR
+ VPWR _21232_/X sky130_fd_sc_hd__mux4_1
X_34198_ _35664_/CLK _34198_/D VGND VGND VPWR VPWR _34198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33149_ _36095_/CLK _33149_/D VGND VGND VPWR VPWR _33149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21163_ _34012_/Q _33948_/Q _33884_/Q _32156_/Q _20914_/X _20915_/X VGND VGND VPWR
+ VPWR _21163_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20114_ _33215_/Q _32575_/Q _35967_/Q _35903_/Q _20080_/X _20081_/X VGND VGND VPWR
+ VPWR _20114_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25971_ _25971_/A VGND VGND VPWR VPWR _33403_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21094_ _22458_/A VGND VGND VPWR VPWR _21094_/X sky130_fd_sc_hd__buf_4
XFILLER_58_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_286_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _36028_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27710_ _34195_/Q _24261_/X _27718_/S VGND VGND VPWR VPWR _27711_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_1193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20045_ _34813_/Q _34749_/Q _34685_/Q _34621_/Q _19941_/X _19942_/X VGND VGND VPWR
+ VPWR _20045_/X sky130_fd_sc_hd__mux4_1
XFILLER_24_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24922_ _24922_/A VGND VGND VPWR VPWR _32941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28690_ _28690_/A VGND VGND VPWR VPWR _34659_/D sky130_fd_sc_hd__clkbuf_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24853_ _24853_/A VGND VGND VPWR VPWR _32909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27641_ _27641_/A VGND VGND VPWR VPWR _34162_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23804_ _23804_/A VGND VGND VPWR VPWR _32446_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27572_ _27572_/A VGND VGND VPWR VPWR _34129_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 _32128_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24784_ _22972_/X _32876_/Q _24802_/S VGND VGND VPWR VPWR _24785_/A sky130_fd_sc_hd__mux2_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _32130_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21996_ _35059_/Q _34995_/Q _34931_/Q _34867_/Q _21756_/X _21757_/X VGND VGND VPWR
+ VPWR _21996_/X sky130_fd_sc_hd__mux4_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26523_ _25150_/X _33665_/Q _26539_/S VGND VGND VPWR VPWR _26524_/A sky130_fd_sc_hd__mux2_1
XANTENNA_127 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29311_ _23234_/X _34923_/Q _29311_/S VGND VGND VPWR VPWR _29312_/A sky130_fd_sc_hd__mux2_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23735_ _23735_/A VGND VGND VPWR VPWR _32413_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20947_ _20743_/X _20945_/X _20946_/X _20746_/X VGND VGND VPWR VPWR _20947_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_149 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29242_ _29242_/A VGND VGND VPWR VPWR _34891_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26454_ _26454_/A VGND VGND VPWR VPWR _33632_/D sky130_fd_sc_hd__clkbuf_1
X_23666_ _23666_/A VGND VGND VPWR VPWR _32382_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20878_ _20874_/X _20877_/X _20611_/X VGND VGND VPWR VPWR _20908_/A sky130_fd_sc_hd__o21ba_2
XFILLER_230_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25405_ _25405_/A VGND VGND VPWR VPWR _33139_/D sky130_fd_sc_hd__clkbuf_1
X_22617_ _22369_/X _22615_/X _22616_/X _22373_/X VGND VGND VPWR VPWR _22617_/X sky130_fd_sc_hd__a22o_1
XFILLER_197_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29173_ _34869_/Q _29172_/X _29173_/S VGND VGND VPWR VPWR _29174_/A sky130_fd_sc_hd__mux2_1
X_26385_ _26412_/S VGND VGND VPWR VPWR _26404_/S sky130_fd_sc_hd__buf_6
X_23597_ _23597_/A VGND VGND VPWR VPWR _32349_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_210_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _35845_/CLK sky130_fd_sc_hd__clkbuf_16
X_28124_ _28124_/A VGND VGND VPWR VPWR _34391_/D sky130_fd_sc_hd__clkbuf_1
X_25336_ _25336_/A VGND VGND VPWR VPWR _33106_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22548_ _22361_/X _22546_/X _22547_/X _22367_/X VGND VGND VPWR VPWR _22548_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_5_9_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_9_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_28055_ _28055_/A VGND VGND VPWR VPWR _34358_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25267_ _25267_/A VGND VGND VPWR VPWR _33074_/D sky130_fd_sc_hd__clkbuf_1
X_22479_ _33281_/Q _36161_/Q _33153_/Q _33089_/Q _22364_/X _22365_/X VGND VGND VPWR
+ VPWR _22479_/X sky130_fd_sc_hd__mux4_1
X_27006_ _27005_/X _33865_/Q _27006_/S VGND VGND VPWR VPWR _27007_/A sky130_fd_sc_hd__mux2_1
X_24218_ _23038_/X _32641_/Q _24234_/S VGND VGND VPWR VPWR _24219_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25198_ _25198_/A VGND VGND VPWR VPWR _33041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24149_ _24149_/A VGND VGND VPWR VPWR _32608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28957_ _34786_/Q _24307_/X _28975_/S VGND VGND VPWR VPWR _28958_/A sky130_fd_sc_hd__mux2_1
X_16971_ _16796_/X _16969_/X _16970_/X _16799_/X VGND VGND VPWR VPWR _16971_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_277_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _34298_/CLK sky130_fd_sc_hd__clkbuf_16
X_18710_ _18387_/X _18708_/X _18709_/X _18397_/X VGND VGND VPWR VPWR _18710_/X sky130_fd_sc_hd__a22o_1
XTAP_5030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27908_ _34289_/Q _24354_/X _27916_/S VGND VGND VPWR VPWR _27909_/A sky130_fd_sc_hd__mux2_1
XTAP_5041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19690_ _19652_/X _19688_/X _19689_/X _19655_/X VGND VGND VPWR VPWR _19690_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28888_ _28888_/A VGND VGND VPWR VPWR _34753_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18641_ _18641_/A VGND VGND VPWR VPWR _32085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27839_ _34256_/Q _24252_/X _27853_/S VGND VGND VPWR VPWR _27840_/A sky130_fd_sc_hd__mux2_1
XTAP_5085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18572_ _33748_/Q _33684_/Q _33620_/Q _33556_/Q _18437_/X _18438_/X VGND VGND VPWR
+ VPWR _18572_/X sky130_fd_sc_hd__mux4_1
X_30850_ _23316_/X _35652_/Q _30860_/S VGND VGND VPWR VPWR _30851_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29509_ _23333_/X _35017_/Q _29509_/S VGND VGND VPWR VPWR _29510_/A sky130_fd_sc_hd__mux2_1
XTAP_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17523_ _17202_/X _17521_/X _17522_/X _17205_/X VGND VGND VPWR VPWR _17523_/X sky130_fd_sc_hd__a22o_1
XTAP_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30781_ _23152_/X _35619_/Q _30797_/S VGND VGND VPWR VPWR _30782_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_650 _20206_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_661 _20423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32520_ _35975_/CLK _32520_/D VGND VGND VPWR VPWR _32520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_672 _22460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17454_ _33013_/Q _32949_/Q _32885_/Q _32821_/Q _17342_/X _17343_/X VGND VGND VPWR
+ VPWR _17454_/X sky130_fd_sc_hd__mux4_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1097 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_683 _22434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_694 _22595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16405_ _34775_/Q _34711_/Q _34647_/Q _34583_/Q _16229_/X _16230_/X VGND VGND VPWR
+ VPWR _16405_/X sky130_fd_sc_hd__mux4_1
X_32451_ _34562_/CLK _32451_/D VGND VGND VPWR VPWR _32451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17385_ _35827_/Q _32205_/Q _35699_/Q _35635_/Q _17313_/X _17314_/X VGND VGND VPWR
+ VPWR _17385_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_201_CLK clkbuf_6_54__f_CLK/X VGND VGND VPWR VPWR _36034_/CLK sky130_fd_sc_hd__clkbuf_16
X_31402_ _35914_/Q input57/X _31408_/S VGND VGND VPWR VPWR _31403_/A sky130_fd_sc_hd__mux2_1
X_19124_ _19010_/X _19122_/X _19123_/X _19014_/X VGND VGND VPWR VPWR _19124_/X sky130_fd_sc_hd__a22o_1
XFILLER_201_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16336_ _34517_/Q _32405_/Q _34389_/Q _34325_/Q _16166_/X _16167_/X VGND VGND VPWR
+ VPWR _16336_/X sky130_fd_sc_hd__mux4_1
X_35170_ _35298_/CLK _35170_/D VGND VGND VPWR VPWR _35170_/Q sky130_fd_sc_hd__dfxtp_1
X_32382_ _36033_/CLK _32382_/D VGND VGND VPWR VPWR _32382_/Q sky130_fd_sc_hd__dfxtp_1
X_34121_ _34816_/CLK _34121_/D VGND VGND VPWR VPWR _34121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16267_ _35027_/Q _34963_/Q _34899_/Q _34835_/Q _16092_/X _16094_/X VGND VGND VPWR
+ VPWR _16267_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19055_ _33185_/Q _32545_/Q _35937_/Q _35873_/Q _19021_/X _19022_/X VGND VGND VPWR
+ VPWR _19055_/X sky130_fd_sc_hd__mux4_1
X_31333_ _35881_/Q input20/X _31337_/S VGND VGND VPWR VPWR _31334_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18006_ _34309_/Q _34245_/Q _34181_/Q _34117_/Q _17795_/X _17796_/X VGND VGND VPWR
+ VPWR _18006_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34052_ _34306_/CLK _34052_/D VGND VGND VPWR VPWR _34052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31264_ _31264_/A VGND VGND VPWR VPWR _35848_/D sky130_fd_sc_hd__clkbuf_1
X_16198_ _35281_/Q _35217_/Q _35153_/Q _32273_/Q _16079_/X _16081_/X VGND VGND VPWR
+ VPWR _16198_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33003_ _36137_/CLK _33003_/D VGND VGND VPWR VPWR _33003_/Q sky130_fd_sc_hd__dfxtp_1
X_30215_ _30215_/A VGND VGND VPWR VPWR _35351_/D sky130_fd_sc_hd__clkbuf_1
X_31195_ _31195_/A VGND VGND VPWR VPWR _35815_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30146_ _30146_/A VGND VGND VPWR VPWR _35318_/D sky130_fd_sc_hd__clkbuf_1
X_19957_ _19855_/X _19955_/X _19956_/X _19858_/X VGND VGND VPWR VPWR _19957_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_268_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _33793_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18908_ _20096_/A VGND VGND VPWR VPWR _18908_/X sky130_fd_sc_hd__clkbuf_4
X_34954_ _35788_/CLK _34954_/D VGND VGND VPWR VPWR _34954_/Q sky130_fd_sc_hd__dfxtp_1
X_30077_ _35286_/Q _29076_/X _30079_/S VGND VGND VPWR VPWR _30078_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19888_ _19848_/X _19886_/X _19887_/X _19853_/X VGND VGND VPWR VPWR _19888_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1060 _16623_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1071 _17128_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1082 _17194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33905_ _34286_/CLK _33905_/D VGND VGND VPWR VPWR _33905_/Q sky130_fd_sc_hd__dfxtp_1
X_18839_ _18657_/X _18837_/X _18838_/X _18661_/X VGND VGND VPWR VPWR _18839_/X sky130_fd_sc_hd__a22o_1
XANTENNA_1093 _17264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34885_ _35781_/CLK _34885_/D VGND VGND VPWR VPWR _34885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33836_ _35054_/CLK _33836_/D VGND VGND VPWR VPWR _33836_/Q sky130_fd_sc_hd__dfxtp_1
X_21850_ _22556_/A VGND VGND VPWR VPWR _21850_/X sky130_fd_sc_hd__buf_6
XFILLER_208_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20801_ _35025_/Q _34961_/Q _34897_/Q _34833_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _20801_/X sky130_fd_sc_hd__mux4_1
XFILLER_24_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33767_ _34279_/CLK _33767_/D VGND VGND VPWR VPWR _33767_/Q sky130_fd_sc_hd__dfxtp_1
X_21781_ _21594_/X _21779_/X _21780_/X _21597_/X VGND VGND VPWR VPWR _21781_/X sky130_fd_sc_hd__a22o_1
XFILLER_58_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30979_ _35713_/Q _29210_/X _30995_/S VGND VGND VPWR VPWR _30980_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23520_ _23016_/X _32314_/Q _23530_/S VGND VGND VPWR VPWR _23521_/A sky130_fd_sc_hd__mux2_1
X_35506_ _36018_/CLK _35506_/D VGND VGND VPWR VPWR _35506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_440_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _33255_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_224_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20732_ _20687_/X _20730_/X _20731_/X _20697_/X VGND VGND VPWR VPWR _20732_/X sky130_fd_sc_hd__a22o_1
XFILLER_169_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32718_ _36049_/CLK _32718_/D VGND VGND VPWR VPWR _32718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33698_ _34276_/CLK _33698_/D VGND VGND VPWR VPWR _33698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35437_ _35562_/CLK _35437_/D VGND VGND VPWR VPWR _35437_/Q sky130_fd_sc_hd__dfxtp_1
X_23451_ _22914_/X _32281_/Q _23467_/S VGND VGND VPWR VPWR _23452_/A sky130_fd_sc_hd__mux2_1
X_20663_ _22531_/A VGND VGND VPWR VPWR _20663_/X sky130_fd_sc_hd__buf_6
X_32649_ _36105_/CLK _32649_/D VGND VGND VPWR VPWR _32649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22402_ _22398_/X _22401_/X _22081_/X VGND VGND VPWR VPWR _22424_/A sky130_fd_sc_hd__o21ba_1
XFILLER_195_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26170_ _26170_/A VGND VGND VPWR VPWR _33497_/D sky130_fd_sc_hd__clkbuf_1
X_23382_ _32250_/Q _23283_/X _23392_/S VGND VGND VPWR VPWR _23383_/A sky130_fd_sc_hd__mux2_1
X_35368_ _35945_/CLK _35368_/D VGND VGND VPWR VPWR _35368_/Q sky130_fd_sc_hd__dfxtp_1
X_20594_ input73/X input74/X VGND VGND VPWR VPWR _20595_/A sky130_fd_sc_hd__and2_1
XFILLER_164_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25121_ _25121_/A VGND VGND VPWR VPWR _33015_/D sky130_fd_sc_hd__clkbuf_1
X_34319_ _34638_/CLK _34319_/D VGND VGND VPWR VPWR _34319_/Q sky130_fd_sc_hd__dfxtp_1
X_22333_ _22008_/X _22331_/X _22332_/X _22014_/X VGND VGND VPWR VPWR _22333_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35299_ _35299_/CLK _35299_/D VGND VGND VPWR VPWR _35299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25052_ _25052_/A VGND VGND VPWR VPWR _32993_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22264_ _22016_/X _22262_/X _22263_/X _22020_/X VGND VGND VPWR VPWR _22264_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24003_ _24003_/A VGND VGND VPWR VPWR _32539_/D sky130_fd_sc_hd__clkbuf_1
X_21215_ _21211_/X _21214_/X _21041_/X VGND VGND VPWR VPWR _21223_/C sky130_fd_sc_hd__o21ba_1
XFILLER_191_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29860_ _35183_/Q _29154_/X _29872_/S VGND VGND VPWR VPWR _29861_/A sky130_fd_sc_hd__mux2_1
X_22195_ _22008_/X _22193_/X _22194_/X _22014_/X VGND VGND VPWR VPWR _22195_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28811_ _26869_/X _34717_/Q _28819_/S VGND VGND VPWR VPWR _28812_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21146_ _35547_/Q _35483_/Q _35419_/Q _35355_/Q _21144_/X _21145_/X VGND VGND VPWR
+ VPWR _21146_/X sky130_fd_sc_hd__mux4_1
X_29791_ _35150_/Q _29048_/X _29809_/S VGND VGND VPWR VPWR _29792_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_259_CLK clkbuf_6_60__f_CLK/X VGND VGND VPWR VPWR _33026_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28742_ _28742_/A VGND VGND VPWR VPWR _34684_/D sky130_fd_sc_hd__clkbuf_1
X_21077_ _33177_/Q _32537_/Q _35929_/Q _35865_/Q _20968_/X _20969_/X VGND VGND VPWR
+ VPWR _21077_/X sky130_fd_sc_hd__mux4_1
X_25954_ _25954_/A VGND VGND VPWR VPWR _33395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20028_ _34045_/Q _33981_/Q _33917_/Q _32253_/Q _20026_/X _20027_/X VGND VGND VPWR
+ VPWR _20028_/X sky130_fd_sc_hd__mux4_1
X_24905_ _24905_/A VGND VGND VPWR VPWR _32933_/D sky130_fd_sc_hd__clkbuf_1
X_25885_ _25885_/A VGND VGND VPWR VPWR _33362_/D sky130_fd_sc_hd__clkbuf_1
X_28673_ _28673_/A VGND VGND VPWR VPWR _34651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27624_ _27624_/A VGND VGND VPWR VPWR _34154_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24836_ _23050_/X _32901_/Q _24844_/S VGND VGND VPWR VPWR _24837_/A sky130_fd_sc_hd__mux2_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27555_ _27011_/X _34123_/Q _27559_/S VGND VGND VPWR VPWR _27556_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24767_ _22948_/X _32868_/Q _24781_/S VGND VGND VPWR VPWR _24768_/A sky130_fd_sc_hd__mux2_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21979_ _33267_/Q _36147_/Q _33139_/Q _33075_/Q _21658_/X _21659_/X VGND VGND VPWR
+ VPWR _21979_/X sky130_fd_sc_hd__mux4_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_431_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _34282_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_226_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23718_ _23718_/A VGND VGND VPWR VPWR _32405_/D sky130_fd_sc_hd__clkbuf_1
X_26506_ _25125_/X _33657_/Q _26518_/S VGND VGND VPWR VPWR _26507_/A sky130_fd_sc_hd__mux2_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27486_ _26909_/X _34090_/Q _27488_/S VGND VGND VPWR VPWR _27487_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24698_ _24698_/A VGND VGND VPWR VPWR _32836_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29225_ input52/X VGND VGND VPWR VPWR _29225_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26437_ _25022_/X _33624_/Q _26455_/S VGND VGND VPWR VPWR _26438_/A sky130_fd_sc_hd__mux2_1
X_23649_ _32374_/Q _23270_/X _23667_/S VGND VGND VPWR VPWR _23650_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17170_ _16849_/X _17168_/X _17169_/X _16852_/X VGND VGND VPWR VPWR _17170_/X sky130_fd_sc_hd__a22o_1
X_29156_ _29156_/A VGND VGND VPWR VPWR _34863_/D sky130_fd_sc_hd__clkbuf_1
X_26368_ _26368_/A VGND VGND VPWR VPWR _33591_/D sky130_fd_sc_hd__clkbuf_1
X_16121_ _35727_/Q _35087_/Q _34447_/Q _33807_/Q _16049_/X _16051_/X VGND VGND VPWR
+ VPWR _16121_/X sky130_fd_sc_hd__mux4_1
X_28107_ _26826_/X _34383_/Q _28123_/S VGND VGND VPWR VPWR _28108_/A sky130_fd_sc_hd__mux2_1
X_25319_ _25319_/A VGND VGND VPWR VPWR _33099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26299_ _25019_/X _33559_/Q _26299_/S VGND VGND VPWR VPWR _26300_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29087_ _34841_/Q _29086_/X _29111_/S VGND VGND VPWR VPWR _29088_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16052_ _35726_/Q _35086_/Q _34446_/Q _33806_/Q _16049_/X _16051_/X VGND VGND VPWR
+ VPWR _16052_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28038_ _28038_/A VGND VGND VPWR VPWR _34350_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1052 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_CLK CLK VGND VGND VPWR VPWR clkbuf_0_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_123_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30000_ _30000_/A VGND VGND VPWR VPWR _35249_/D sky130_fd_sc_hd__clkbuf_1
X_19811_ _35062_/Q _34998_/Q _34934_/Q _34870_/Q _19809_/X _19810_/X VGND VGND VPWR
+ VPWR _19811_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29989_ _35244_/Q _29144_/X _30007_/S VGND VGND VPWR VPWR _29990_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19742_ _20256_/A VGND VGND VPWR VPWR _19742_/X sky130_fd_sc_hd__buf_4
X_16954_ _33255_/Q _36135_/Q _33127_/Q _33063_/Q _16705_/X _16706_/X VGND VGND VPWR
+ VPWR _16954_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31951_ _34973_/CLK _31951_/D VGND VGND VPWR VPWR _31951_/Q sky130_fd_sc_hd__dfxtp_1
X_19673_ _20146_/A VGND VGND VPWR VPWR _19673_/X sky130_fd_sc_hd__buf_4
XFILLER_49_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16885_ _16849_/X _16883_/X _16884_/X _16852_/X VGND VGND VPWR VPWR _16885_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18624_ _18326_/X _18622_/X _18623_/X _18337_/X VGND VGND VPWR VPWR _18624_/X sky130_fd_sc_hd__a22o_1
XFILLER_49_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30902_ _30902_/A VGND VGND VPWR VPWR _35676_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34670_ _35304_/CLK _34670_/D VGND VGND VPWR VPWR _34670_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31882_ _23241_/X _36141_/Q _31898_/S VGND VGND VPWR VPWR _31883_/A sky130_fd_sc_hd__mux2_1
XTAP_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33621_ _33685_/CLK _33621_/D VGND VGND VPWR VPWR _33621_/Q sky130_fd_sc_hd__dfxtp_1
X_30833_ _23289_/X _35644_/Q _30839_/S VGND VGND VPWR VPWR _30834_/A sky130_fd_sc_hd__mux2_1
X_18555_ _20096_/A VGND VGND VPWR VPWR _18555_/X sky130_fd_sc_hd__buf_4
XFILLER_240_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_422_CLK clkbuf_6_36__f_CLK/X VGND VGND VPWR VPWR _36074_/CLK sky130_fd_sc_hd__clkbuf_16
X_17506_ _17502_/X _17503_/X _17504_/X _17505_/X VGND VGND VPWR VPWR _17506_/X sky130_fd_sc_hd__a22o_1
X_33552_ _34194_/CLK _33552_/D VGND VGND VPWR VPWR _33552_/Q sky130_fd_sc_hd__dfxtp_1
X_18486_ _18326_/X _18484_/X _18485_/X _18337_/X VGND VGND VPWR VPWR _18486_/X sky130_fd_sc_hd__a22o_1
X_30764_ _23127_/X _35611_/Q _30776_/S VGND VGND VPWR VPWR _30765_/A sky130_fd_sc_hd__mux2_1
XANTENNA_480 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_491 _31994_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32503_ _36022_/CLK _32503_/D VGND VGND VPWR VPWR _32503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17437_ _17154_/X _17435_/X _17436_/X _17159_/X VGND VGND VPWR VPWR _17437_/X sky130_fd_sc_hd__a22o_1
X_33483_ _36107_/CLK _33483_/D VGND VGND VPWR VPWR _33483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30695_ _30695_/A VGND VGND VPWR VPWR _35578_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_16 _32115_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35222_ _35286_/CLK _35222_/D VGND VGND VPWR VPWR _35222_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_27 _32116_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_38 _32117_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32434_ _34866_/CLK _32434_/D VGND VGND VPWR VPWR _32434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_49 _32119_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17368_ _17368_/A VGND VGND VPWR VPWR _31986_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_1433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19107_ _19101_/X _19102_/X _19105_/X _19106_/X VGND VGND VPWR VPWR _19107_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35153_ _36216_/CLK _35153_/D VGND VGND VPWR VPWR _35153_/Q sky130_fd_sc_hd__dfxtp_1
X_16319_ _32725_/Q _32661_/Q _32597_/Q _36053_/Q _16213_/X _17713_/A VGND VGND VPWR
+ VPWR _16319_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32365_ _36013_/CLK _32365_/D VGND VGND VPWR VPWR _32365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17299_ _33777_/Q _33713_/Q _33649_/Q _33585_/Q _17196_/X _17197_/X VGND VGND VPWR
+ VPWR _17299_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34104_ _36152_/CLK _34104_/D VGND VGND VPWR VPWR _34104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19038_ _34273_/Q _34209_/Q _34145_/Q _34081_/Q _19036_/X _19037_/X VGND VGND VPWR
+ VPWR _19038_/X sky130_fd_sc_hd__mux4_1
X_31316_ _35873_/Q input11/X _31316_/S VGND VGND VPWR VPWR _31317_/A sky130_fd_sc_hd__mux2_1
X_35084_ _35340_/CLK _35084_/D VGND VGND VPWR VPWR _35084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput101 _31951_/Q VGND VGND VPWR VPWR D1[1] sky130_fd_sc_hd__buf_2
X_32296_ _35179_/CLK _32296_/D VGND VGND VPWR VPWR _32296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput112 _31952_/Q VGND VGND VPWR VPWR D1[2] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_489_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _35809_/CLK sky130_fd_sc_hd__clkbuf_16
Xoutput123 _31953_/Q VGND VGND VPWR VPWR D1[3] sky130_fd_sc_hd__buf_2
X_34035_ _34227_/CLK _34035_/D VGND VGND VPWR VPWR _34035_/Q sky130_fd_sc_hd__dfxtp_1
X_31247_ _35840_/Q input46/X _31265_/S VGND VGND VPWR VPWR _31248_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput134 _31954_/Q VGND VGND VPWR VPWR D1[4] sky130_fd_sc_hd__buf_2
Xoutput145 _31955_/Q VGND VGND VPWR VPWR D1[5] sky130_fd_sc_hd__buf_2
Xoutput156 _36185_/Q VGND VGND VPWR VPWR D2[11] sky130_fd_sc_hd__buf_2
XFILLER_138_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21000_ _20888_/X _20998_/X _20999_/X _20891_/X VGND VGND VPWR VPWR _21000_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput167 _36195_/Q VGND VGND VPWR VPWR D2[21] sky130_fd_sc_hd__buf_2
XFILLER_86_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput178 _36205_/Q VGND VGND VPWR VPWR D2[31] sky130_fd_sc_hd__buf_2
XFILLER_47_1158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput189 _36215_/Q VGND VGND VPWR VPWR D2[41] sky130_fd_sc_hd__buf_2
XFILLER_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31178_ _31178_/A VGND VGND VPWR VPWR _35807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30129_ _30129_/A VGND VGND VPWR VPWR _35310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35986_ _35986_/CLK _35986_/D VGND VGND VPWR VPWR _35986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34937_ _35386_/CLK _34937_/D VGND VGND VPWR VPWR _34937_/Q sky130_fd_sc_hd__dfxtp_1
X_22951_ input16/X VGND VGND VPWR VPWR _22951_/X sky130_fd_sc_hd__buf_2
XFILLER_68_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21902_ _33521_/Q _33457_/Q _33393_/Q _33329_/Q _21723_/X _21724_/X VGND VGND VPWR
+ VPWR _21902_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25670_ _25670_/A VGND VGND VPWR VPWR _33261_/D sky130_fd_sc_hd__clkbuf_1
X_22882_ _22882_/A VGND VGND VPWR VPWR _32014_/D sky130_fd_sc_hd__clkbuf_1
X_34868_ _34932_/CLK _34868_/D VGND VGND VPWR VPWR _34868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24621_ _22935_/X _32800_/Q _24623_/S VGND VGND VPWR VPWR _24622_/A sky130_fd_sc_hd__mux2_1
X_33819_ _35098_/CLK _33819_/D VGND VGND VPWR VPWR _33819_/Q sky130_fd_sc_hd__dfxtp_1
X_21833_ _33775_/Q _33711_/Q _33647_/Q _33583_/Q _21796_/X _21797_/X VGND VGND VPWR
+ VPWR _21833_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34799_ _34866_/CLK _34799_/D VGND VGND VPWR VPWR _34799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_413_CLK clkbuf_6_33__f_CLK/X VGND VGND VPWR VPWR _35242_/CLK sky130_fd_sc_hd__clkbuf_16
X_27340_ _27340_/A VGND VGND VPWR VPWR _34020_/D sky130_fd_sc_hd__clkbuf_1
X_24552_ _24552_/A VGND VGND VPWR VPWR _32768_/D sky130_fd_sc_hd__clkbuf_1
X_21764_ _21764_/A VGND VGND VPWR VPWR _36204_/D sky130_fd_sc_hd__buf_6
XFILLER_19_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23503_ _22991_/X _32306_/Q _23509_/S VGND VGND VPWR VPWR _23504_/A sky130_fd_sc_hd__mux2_1
X_27271_ _26990_/X _33988_/Q _27281_/S VGND VGND VPWR VPWR _27272_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_6_54__f_CLK clkbuf_5_27_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_54__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20715_ _20614_/X _20713_/X _20714_/X _20623_/X VGND VGND VPWR VPWR _20715_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24483_ _22935_/X _32736_/Q _24485_/S VGND VGND VPWR VPWR _24484_/A sky130_fd_sc_hd__mux2_1
X_21695_ _21449_/X _21693_/X _21694_/X _21452_/X VGND VGND VPWR VPWR _21695_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29010_ _29010_/A VGND VGND VPWR VPWR _34811_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26222_ _26222_/A VGND VGND VPWR VPWR _33522_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23434_ _22889_/X _32273_/Q _23446_/S VGND VGND VPWR VPWR _23435_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20646_ _22396_/A VGND VGND VPWR VPWR _20646_/X sky130_fd_sc_hd__buf_6
XFILLER_165_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26153_ _26153_/A VGND VGND VPWR VPWR _33489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23365_ _32242_/Q _23256_/X _23371_/S VGND VGND VPWR VPWR _23366_/A sky130_fd_sc_hd__mux2_1
X_20577_ _22455_/A VGND VGND VPWR VPWR _20577_/X sky130_fd_sc_hd__buf_4
XFILLER_20_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25104_ _25103_/X _33010_/Q _25113_/S VGND VGND VPWR VPWR _25105_/A sky130_fd_sc_hd__mux2_1
X_22316_ _34556_/Q _32444_/Q _34428_/Q _34364_/Q _22178_/X _22179_/X VGND VGND VPWR
+ VPWR _22316_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26084_ _25100_/X _33457_/Q _26092_/S VGND VGND VPWR VPWR _26085_/A sky130_fd_sc_hd__mux2_1
X_23296_ _23296_/A VGND VGND VPWR VPWR _32216_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29912_ _35208_/Q _29231_/X _29914_/S VGND VGND VPWR VPWR _29913_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25035_ input6/X VGND VGND VPWR VPWR _25035_/X sky130_fd_sc_hd__buf_2
X_22247_ _35066_/Q _35002_/Q _34938_/Q _34874_/Q _22109_/X _22110_/X VGND VGND VPWR
+ VPWR _22247_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29843_ _35175_/Q _29129_/X _29851_/S VGND VGND VPWR VPWR _29844_/A sky130_fd_sc_hd__mux2_1
X_22178_ _22531_/A VGND VGND VPWR VPWR _22178_/X sky130_fd_sc_hd__buf_6
XFILLER_78_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21129_ _21089_/X _21127_/X _21128_/X _21094_/X VGND VGND VPWR VPWR _21129_/X sky130_fd_sc_hd__a22o_1
X_29774_ _29774_/A VGND VGND VPWR VPWR _35142_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26986_ _26986_/A VGND VGND VPWR VPWR _33858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28725_ _28725_/A VGND VGND VPWR VPWR _34676_/D sky130_fd_sc_hd__clkbuf_1
X_25937_ _25937_/A VGND VGND VPWR VPWR _33387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28656_ _28656_/A VGND VGND VPWR VPWR _34643_/D sky130_fd_sc_hd__clkbuf_1
X_16670_ _16496_/X _16666_/X _16669_/X _16499_/X VGND VGND VPWR VPWR _16670_/X sky130_fd_sc_hd__a22o_1
X_25868_ _25180_/X _33355_/Q _25872_/S VGND VGND VPWR VPWR _25869_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27607_ _34146_/Q _24307_/X _27625_/S VGND VGND VPWR VPWR _27608_/A sky130_fd_sc_hd__mux2_1
XFILLER_234_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24819_ _23025_/X _32893_/Q _24823_/S VGND VGND VPWR VPWR _24820_/A sky130_fd_sc_hd__mux2_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28587_ _26937_/X _34611_/Q _28591_/S VGND VGND VPWR VPWR _28588_/A sky130_fd_sc_hd__mux2_1
X_25799_ _25078_/X _33322_/Q _25801_/S VGND VGND VPWR VPWR _25800_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_404_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _35945_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _20142_/A VGND VGND VPWR VPWR _18340_/X sky130_fd_sc_hd__buf_2
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27538_ _27538_/A VGND VGND VPWR VPWR _34114_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18271_ _16056_/X _18269_/X _18270_/X _16068_/X VGND VGND VPWR VPWR _18271_/X sky130_fd_sc_hd__a22o_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27469_ _27559_/S VGND VGND VPWR VPWR _27488_/S sky130_fd_sc_hd__buf_4
XFILLER_204_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29208_ _34880_/Q _29206_/X _29235_/S VGND VGND VPWR VPWR _29209_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17222_ _34798_/Q _34734_/Q _34670_/Q _34606_/Q _16935_/X _16936_/X VGND VGND VPWR
+ VPWR _17222_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30480_ _30480_/A VGND VGND VPWR VPWR _35476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput14 DW[21] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_8
Xinput25 DW[31] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_4
X_17153_ _17149_/X _17150_/X _17151_/X _17152_/X VGND VGND VPWR VPWR _17153_/X sky130_fd_sc_hd__a22o_1
X_29139_ _34858_/Q _29138_/X _29142_/S VGND VGND VPWR VPWR _29140_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput36 DW[41] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__buf_4
XFILLER_167_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput47 DW[51] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__buf_8
X_16104_ _33743_/Q _33679_/Q _33615_/Q _33551_/Q _15980_/X _15983_/X VGND VGND VPWR
+ VPWR _16104_/X sky130_fd_sc_hd__mux4_1
Xinput58 DW[61] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__buf_8
Xinput69 R1[4] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__buf_2
X_32150_ _34006_/CLK _32150_/D VGND VGND VPWR VPWR _32150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17084_ _16801_/X _17082_/X _17083_/X _16806_/X VGND VGND VPWR VPWR _17084_/X sky130_fd_sc_hd__a22o_1
XFILLER_156_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31101_ _35771_/Q _29191_/X _31109_/S VGND VGND VPWR VPWR _31102_/A sky130_fd_sc_hd__mux2_1
X_16035_ _17830_/A VGND VGND VPWR VPWR _16035_/X sky130_fd_sc_hd__clkbuf_4
X_32081_ _34973_/CLK _32081_/D VGND VGND VPWR VPWR _32081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31032_ _35738_/Q _29089_/X _31046_/S VGND VGND VPWR VPWR _31033_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35840_ _35971_/CLK _35840_/D VGND VGND VPWR VPWR _35840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17986_ _17981_/X _17985_/X _17842_/X _17843_/X VGND VGND VPWR VPWR _18003_/B sky130_fd_sc_hd__o211a_1
XFILLER_112_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19725_ _19647_/X _19723_/X _19724_/X _19650_/X VGND VGND VPWR VPWR _19725_/X sky130_fd_sc_hd__a22o_1
XFILLER_84_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35771_ _35771_/CLK _35771_/D VGND VGND VPWR VPWR _35771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16937_ _34790_/Q _34726_/Q _34662_/Q _34598_/Q _16935_/X _16936_/X VGND VGND VPWR
+ VPWR _16937_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32983_ _32983_/CLK _32983_/D VGND VGND VPWR VPWR _32983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34722_ _35928_/CLK _34722_/D VGND VGND VPWR VPWR _34722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31934_ _23322_/X _36166_/Q _31940_/S VGND VGND VPWR VPWR _31935_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19656_ _19652_/X _19653_/X _19654_/X _19655_/X VGND VGND VPWR VPWR _19656_/X sky130_fd_sc_hd__a22o_1
X_16868_ _16864_/X _16867_/X _16794_/X VGND VGND VPWR VPWR _16878_/C sky130_fd_sc_hd__o21ba_1
XFILLER_42_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18607_ _18603_/X _18606_/X _18400_/X VGND VGND VPWR VPWR _18608_/D sky130_fd_sc_hd__o21ba_1
X_34653_ _35164_/CLK _34653_/D VGND VGND VPWR VPWR _34653_/Q sky130_fd_sc_hd__dfxtp_1
X_19587_ _19583_/X _19586_/X _19447_/X VGND VGND VPWR VPWR _19597_/C sky130_fd_sc_hd__o21ba_1
X_31865_ _23199_/X _36133_/Q _31877_/S VGND VGND VPWR VPWR _31866_/A sky130_fd_sc_hd__mux2_1
X_16799_ _17152_/A VGND VGND VPWR VPWR _16799_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_206_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33604_ _33795_/CLK _33604_/D VGND VGND VPWR VPWR _33604_/Q sky130_fd_sc_hd__dfxtp_1
X_18538_ _18538_/A _18538_/B _18538_/C _18538_/D VGND VGND VPWR VPWR _18539_/A sky130_fd_sc_hd__or4_4
XFILLER_34_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30816_ _23264_/X _35636_/Q _30818_/S VGND VGND VPWR VPWR _30817_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34584_ _34777_/CLK _34584_/D VGND VGND VPWR VPWR _34584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31796_ _31796_/A VGND VGND VPWR VPWR _36100_/D sky130_fd_sc_hd__clkbuf_1
X_33535_ _34303_/CLK _33535_/D VGND VGND VPWR VPWR _33535_/Q sky130_fd_sc_hd__dfxtp_1
X_18469_ _35024_/Q _34960_/Q _34896_/Q _34832_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _18469_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30747_ _23102_/X _35603_/Q _30755_/S VGND VGND VPWR VPWR _30748_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20500_ _35787_/Q _35147_/Q _34507_/Q _33867_/Q _18408_/X _18409_/X VGND VGND VPWR
+ VPWR _20500_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33466_ _33787_/CLK _33466_/D VGND VGND VPWR VPWR _33466_/Q sky130_fd_sc_hd__dfxtp_1
X_21480_ _33765_/Q _33701_/Q _33637_/Q _33573_/Q _21443_/X _21444_/X VGND VGND VPWR
+ VPWR _21480_/X sky130_fd_sc_hd__mux4_1
XFILLER_193_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30678_ _30678_/A VGND VGND VPWR VPWR _35570_/D sky130_fd_sc_hd__clkbuf_1
X_35205_ _35333_/CLK _35205_/D VGND VGND VPWR VPWR _35205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20431_ _20427_/X _20430_/X _20134_/X VGND VGND VPWR VPWR _20453_/A sky130_fd_sc_hd__o21ba_2
X_32417_ _35296_/CLK _32417_/D VGND VGND VPWR VPWR _32417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36185_ _36185_/CLK _36185_/D VGND VGND VPWR VPWR _36185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33397_ _34292_/CLK _33397_/D VGND VGND VPWR VPWR _33397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35136_ _35843_/CLK _35136_/D VGND VGND VPWR VPWR _35136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23150_ _32162_/Q _23148_/X _23350_/S VGND VGND VPWR VPWR _23151_/A sky130_fd_sc_hd__mux2_1
X_20362_ _20358_/X _20361_/X _20167_/X VGND VGND VPWR VPWR _20363_/D sky130_fd_sc_hd__o21ba_1
XFILLER_173_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32348_ _33244_/CLK _32348_/D VGND VGND VPWR VPWR _32348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22101_ _22096_/X _22099_/X _22100_/X VGND VGND VPWR VPWR _22116_/C sky130_fd_sc_hd__o21ba_1
XTAP_7009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23081_ _30329_/B _29049_/B _30329_/A VGND VGND VPWR VPWR _23082_/A sky130_fd_sc_hd__or3b_1
X_35067_ _35515_/CLK _35067_/D VGND VGND VPWR VPWR _35067_/Q sky130_fd_sc_hd__dfxtp_1
X_20293_ _20289_/X _20292_/X _20153_/X VGND VGND VPWR VPWR _20303_/C sky130_fd_sc_hd__o21ba_1
X_32279_ _36185_/CLK _32279_/D VGND VGND VPWR VPWR _32279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22032_ _34804_/Q _34740_/Q _34676_/Q _34612_/Q _21888_/X _21889_/X VGND VGND VPWR
+ VPWR _22032_/X sky130_fd_sc_hd__mux4_1
X_34018_ _34149_/CLK _34018_/D VGND VGND VPWR VPWR _34018_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26840_ _26840_/A VGND VGND VPWR VPWR _33811_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23983_ _22892_/X _32530_/Q _23993_/S VGND VGND VPWR VPWR _23984_/A sky130_fd_sc_hd__mux2_1
X_26771_ _26819_/S VGND VGND VPWR VPWR _26790_/S sky130_fd_sc_hd__buf_4
X_35969_ _35970_/CLK _35969_/D VGND VGND VPWR VPWR _35969_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28510_ _26821_/X _34574_/Q _28528_/S VGND VGND VPWR VPWR _28511_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25722_ _25722_/A VGND VGND VPWR VPWR _33286_/D sky130_fd_sc_hd__clkbuf_1
X_22934_ _22934_/A VGND VGND VPWR VPWR _32031_/D sky130_fd_sc_hd__clkbuf_1
X_29490_ _29517_/S VGND VGND VPWR VPWR _29509_/S sky130_fd_sc_hd__buf_4
XFILLER_228_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28441_ _28441_/A VGND VGND VPWR VPWR _34541_/D sky130_fd_sc_hd__clkbuf_1
X_22865_ _22861_/X _22864_/X _22453_/A VGND VGND VPWR VPWR _22873_/C sky130_fd_sc_hd__o21ba_1
XFILLER_16_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25653_ _25653_/A VGND VGND VPWR VPWR _33253_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21816_ _35758_/Q _35118_/Q _34478_/Q _33838_/Q _21740_/X _21741_/X VGND VGND VPWR
+ VPWR _21816_/X sky130_fd_sc_hd__mux4_1
X_24604_ _24715_/S VGND VGND VPWR VPWR _24623_/S sky130_fd_sc_hd__buf_4
X_28372_ _28372_/A VGND VGND VPWR VPWR _34509_/D sky130_fd_sc_hd__clkbuf_1
X_25584_ _25584_/A VGND VGND VPWR VPWR _33222_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22796_ _33035_/Q _32971_/Q _32907_/Q _32843_/Q _20580_/X _20583_/X VGND VGND VPWR
+ VPWR _22796_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24535_ _24535_/A VGND VGND VPWR VPWR _32760_/D sky130_fd_sc_hd__clkbuf_1
X_27323_ _27323_/A VGND VGND VPWR VPWR _34012_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21747_ _22453_/A VGND VGND VPWR VPWR _21747_/X sky130_fd_sc_hd__buf_4
XPHY_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27254_ _26965_/X _33980_/Q _27260_/S VGND VGND VPWR VPWR _27255_/A sky130_fd_sc_hd__mux2_1
X_24466_ _24577_/S VGND VGND VPWR VPWR _24485_/S sky130_fd_sc_hd__buf_6
XFILLER_185_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21678_ _21672_/X _21677_/X _21394_/X VGND VGND VPWR VPWR _21686_/C sky130_fd_sc_hd__o21ba_1
XFILLER_32_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23417_ _32267_/Q _23339_/X _23421_/S VGND VGND VPWR VPWR _23418_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26205_ _26205_/A VGND VGND VPWR VPWR _33514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20629_ _20659_/A VGND VGND VPWR VPWR _22370_/A sky130_fd_sc_hd__buf_12
X_27185_ _26863_/X _33947_/Q _27197_/S VGND VGND VPWR VPWR _27186_/A sky130_fd_sc_hd__mux2_1
X_24397_ input44/X VGND VGND VPWR VPWR _24397_/X sky130_fd_sc_hd__clkbuf_4
X_26136_ _25177_/X _33482_/Q _26142_/S VGND VGND VPWR VPWR _26137_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23348_ _32234_/Q _23231_/X _23350_/S VGND VGND VPWR VPWR _23349_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26067_ _25075_/X _33449_/Q _26071_/S VGND VGND VPWR VPWR _26068_/A sky130_fd_sc_hd__mux2_1
X_23279_ _23279_/A VGND VGND VPWR VPWR _32210_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25018_ _25018_/A VGND VGND VPWR VPWR _32982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17840_ _33024_/Q _32960_/Q _32896_/Q _32832_/Q _17695_/X _17696_/X VGND VGND VPWR
+ VPWR _17840_/X sky130_fd_sc_hd__mux4_1
X_29826_ _35167_/Q _29104_/X _29830_/S VGND VGND VPWR VPWR _29827_/A sky130_fd_sc_hd__mux2_1
XTAP_6853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17771_ _32510_/Q _32382_/Q _32062_/Q _36030_/Q _17629_/X _17770_/X VGND VGND VPWR
+ VPWR _17771_/X sky130_fd_sc_hd__mux4_1
X_29757_ _29757_/A VGND VGND VPWR VPWR _35134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26969_ _26968_/X _33853_/Q _26975_/S VGND VGND VPWR VPWR _26970_/A sky130_fd_sc_hd__mux2_1
X_19510_ _19355_/X _19508_/X _19509_/X _19361_/X VGND VGND VPWR VPWR _19510_/X sky130_fd_sc_hd__a22o_1
X_16722_ _17932_/A VGND VGND VPWR VPWR _16722_/X sky130_fd_sc_hd__buf_4
XFILLER_47_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28708_ _26915_/X _34668_/Q _28726_/S VGND VGND VPWR VPWR _28709_/A sky130_fd_sc_hd__mux2_1
X_29688_ _29688_/A VGND VGND VPWR VPWR _35101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19441_ _20295_/A VGND VGND VPWR VPWR _19441_/X sky130_fd_sc_hd__buf_4
X_28639_ _27014_/X _34636_/Q _28641_/S VGND VGND VPWR VPWR _28640_/A sky130_fd_sc_hd__mux2_1
X_16653_ _17712_/A VGND VGND VPWR VPWR _16653_/X sky130_fd_sc_hd__buf_6
XFILLER_165_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31650_ _31650_/A VGND VGND VPWR VPWR _36031_/D sky130_fd_sc_hd__clkbuf_1
X_19372_ _19294_/X _19370_/X _19371_/X _19297_/X VGND VGND VPWR VPWR _19372_/X sky130_fd_sc_hd__a22o_1
X_16584_ _34780_/Q _34716_/Q _34652_/Q _34588_/Q _16582_/X _16583_/X VGND VGND VPWR
+ VPWR _16584_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30601_ _30733_/S VGND VGND VPWR VPWR _30620_/S sky130_fd_sc_hd__buf_4
X_18323_ _20206_/A VGND VGND VPWR VPWR _18323_/X sky130_fd_sc_hd__buf_2
XFILLER_128_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31581_ _31581_/A VGND VGND VPWR VPWR _35998_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33320_ _34278_/CLK _33320_/D VGND VGND VPWR VPWR _33320_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ _17149_/A _18252_/X _18253_/X _17152_/A VGND VGND VPWR VPWR _18254_/X sky130_fd_sc_hd__a22o_1
X_30532_ _23241_/X _35501_/Q _30548_/S VGND VGND VPWR VPWR _30533_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17205_ _17911_/A VGND VGND VPWR VPWR _17205_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_141_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33251_ _36132_/CLK _33251_/D VGND VGND VPWR VPWR _33251_/Q sky130_fd_sc_hd__dfxtp_1
X_18185_ _33803_/Q _33739_/Q _33675_/Q _33611_/Q _17902_/X _17903_/X VGND VGND VPWR
+ VPWR _18185_/X sky130_fd_sc_hd__mux4_1
X_30463_ _23345_/X _35469_/Q _30463_/S VGND VGND VPWR VPWR _30464_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32202_ _35955_/CLK _32202_/D VGND VGND VPWR VPWR _32202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17136_ _17842_/A VGND VGND VPWR VPWR _17136_/X sky130_fd_sc_hd__clkbuf_4
X_33182_ _35935_/CLK _33182_/D VGND VGND VPWR VPWR _33182_/Q sky130_fd_sc_hd__dfxtp_1
X_30394_ _30463_/S VGND VGND VPWR VPWR _30413_/S sky130_fd_sc_hd__buf_6
XFILLER_195_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32133_ _35750_/CLK _32133_/D VGND VGND VPWR VPWR _32133_/Q sky130_fd_sc_hd__dfxtp_1
X_17067_ _17911_/A VGND VGND VPWR VPWR _17067_/X sky130_fd_sc_hd__buf_4
XFILLER_98_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16018_ _17762_/A VGND VGND VPWR VPWR _17713_/A sky130_fd_sc_hd__buf_4
X_32064_ _36032_/CLK _32064_/D VGND VGND VPWR VPWR _32064_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31015_ _35730_/Q _29064_/X _31025_/S VGND VGND VPWR VPWR _31016_/A sky130_fd_sc_hd__mux2_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35823_ _35951_/CLK _35823_/D VGND VGND VPWR VPWR _35823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17969_ _17969_/A _17969_/B _17969_/C _17969_/D VGND VGND VPWR VPWR _17970_/A sky130_fd_sc_hd__or4_4
XFILLER_22_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19708_ _20201_/A VGND VGND VPWR VPWR _19708_/X sky130_fd_sc_hd__clkbuf_4
X_35754_ _35945_/CLK _35754_/D VGND VGND VPWR VPWR _35754_/Q sky130_fd_sc_hd__dfxtp_1
X_32966_ _32967_/CLK _32966_/D VGND VGND VPWR VPWR _32966_/Q sky130_fd_sc_hd__dfxtp_1
X_20980_ _20980_/A _20980_/B _20980_/C _20980_/D VGND VGND VPWR VPWR _20981_/A sky130_fd_sc_hd__or4_1
XFILLER_38_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34705_ _36220_/CLK _34705_/D VGND VGND VPWR VPWR _34705_/Q sky130_fd_sc_hd__dfxtp_1
X_31917_ _23297_/X _36158_/Q _31919_/S VGND VGND VPWR VPWR _31918_/A sky130_fd_sc_hd__mux2_1
X_19639_ _33266_/Q _36146_/Q _33138_/Q _33074_/Q _19358_/X _19359_/X VGND VGND VPWR
+ VPWR _19639_/X sky130_fd_sc_hd__mux4_1
X_35685_ _35748_/CLK _35685_/D VGND VGND VPWR VPWR _35685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_2_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_2_2_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_32897_ _36033_/CLK _32897_/D VGND VGND VPWR VPWR _32897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34636_ _35341_/CLK _34636_/D VGND VGND VPWR VPWR _34636_/Q sky130_fd_sc_hd__dfxtp_1
X_22650_ _35782_/Q _35142_/Q _34502_/Q _33862_/Q _22446_/X _22447_/X VGND VGND VPWR
+ VPWR _22650_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31848_ _23133_/X _36125_/Q _31856_/S VGND VGND VPWR VPWR _31849_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21601_ _33192_/Q _32552_/Q _35944_/Q _35880_/Q _21321_/X _21322_/X VGND VGND VPWR
+ VPWR _21601_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34567_ _35079_/CLK _34567_/D VGND VGND VPWR VPWR _34567_/Q sky130_fd_sc_hd__dfxtp_1
X_22581_ _22361_/X _22579_/X _22580_/X _22367_/X VGND VGND VPWR VPWR _22581_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31779_ _31779_/A VGND VGND VPWR VPWR _36092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24320_ input17/X VGND VGND VPWR VPWR _24320_/X sky130_fd_sc_hd__buf_4
XFILLER_107_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21532_ _33190_/Q _32550_/Q _35942_/Q _35878_/Q _21321_/X _21322_/X VGND VGND VPWR
+ VPWR _21532_/X sky130_fd_sc_hd__mux4_1
X_33518_ _33520_/CLK _33518_/D VGND VGND VPWR VPWR _33518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34498_ _35779_/CLK _34498_/D VGND VGND VPWR VPWR _34498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36237_ _36237_/CLK _36237_/D VGND VGND VPWR VPWR _36237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24251_ _24251_/A VGND VGND VPWR VPWR _32655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33449_ _35386_/CLK _33449_/D VGND VGND VPWR VPWR _33449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21463_ _35748_/Q _35108_/Q _34468_/Q _33828_/Q _21387_/X _21388_/X VGND VGND VPWR
+ VPWR _21463_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23202_ _32183_/Q _23139_/X _23206_/S VGND VGND VPWR VPWR _23203_/A sky130_fd_sc_hd__mux2_1
X_20414_ _18297_/X _20412_/X _20413_/X _18303_/X VGND VGND VPWR VPWR _20414_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36168_ _36168_/CLK _36168_/D VGND VGND VPWR VPWR _36168_/Q sky130_fd_sc_hd__dfxtp_1
X_24182_ _22985_/X _32624_/Q _24192_/S VGND VGND VPWR VPWR _24183_/A sky130_fd_sc_hd__mux2_1
X_21394_ _22453_/A VGND VGND VPWR VPWR _21394_/X sky130_fd_sc_hd__buf_2
XFILLER_88_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35119_ _35822_/CLK _35119_/D VGND VGND VPWR VPWR _35119_/Q sky130_fd_sc_hd__dfxtp_1
X_23133_ input7/X VGND VGND VPWR VPWR _23133_/X sky130_fd_sc_hd__buf_6
X_20345_ _32518_/Q _32390_/Q _32070_/Q _36038_/Q _20282_/X _20070_/X VGND VGND VPWR
+ VPWR _20345_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36099_ _36100_/CLK _36099_/D VGND VGND VPWR VPWR _36099_/Q sky130_fd_sc_hd__dfxtp_1
X_28990_ _34802_/Q _24357_/X _28996_/S VGND VGND VPWR VPWR _28991_/A sky130_fd_sc_hd__mux2_1
XTAP_6105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27941_ _27941_/A VGND VGND VPWR VPWR _34304_/D sky130_fd_sc_hd__clkbuf_1
X_23064_ _23064_/A VGND VGND VPWR VPWR _32073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20276_ _20208_/X _20274_/X _20275_/X _20211_/X VGND VGND VPWR VPWR _20276_/X sky130_fd_sc_hd__a22o_1
XTAP_6116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22015_ _22008_/X _22010_/X _22013_/X _22014_/X VGND VGND VPWR VPWR _22015_/X sky130_fd_sc_hd__a22o_1
XTAP_6149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27872_ _34272_/Q _24301_/X _27874_/S VGND VGND VPWR VPWR _27873_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29611_ _35065_/Q _29185_/X _29623_/S VGND VGND VPWR VPWR _29612_/A sky130_fd_sc_hd__mux2_1
XTAP_5448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26823_ _27018_/S VGND VGND VPWR VPWR _26851_/S sky130_fd_sc_hd__buf_4
XTAP_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29542_ _35032_/Q _29082_/X _29560_/S VGND VGND VPWR VPWR _29543_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26754_ _26754_/A VGND VGND VPWR VPWR _33773_/D sky130_fd_sc_hd__clkbuf_1
X_23966_ _23068_/X _32523_/Q _23970_/S VGND VGND VPWR VPWR _23967_/A sky130_fd_sc_hd__mux2_1
XTAP_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25705_ _25705_/A VGND VGND VPWR VPWR _33278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29473_ _29473_/A VGND VGND VPWR VPWR _34999_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22917_ input4/X VGND VGND VPWR VPWR _22917_/X sky130_fd_sc_hd__buf_4
X_26685_ _31140_/B _26685_/B VGND VGND VPWR VPWR _26686_/A sky130_fd_sc_hd__and2b_1
X_23897_ _22966_/X _32490_/Q _23899_/S VGND VGND VPWR VPWR _23898_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28424_ _28424_/A VGND VGND VPWR VPWR _34533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22848_ _33549_/Q _33485_/Q _33421_/Q _33357_/Q _20633_/X _20635_/X VGND VGND VPWR
+ VPWR _22848_/X sky130_fd_sc_hd__mux4_1
X_25636_ _25636_/A VGND VGND VPWR VPWR _33245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28355_ _34501_/Q _24416_/X _28363_/S VGND VGND VPWR VPWR _28356_/A sky130_fd_sc_hd__mux2_1
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22779_ _34570_/Q _32458_/Q _34442_/Q _34378_/Q _22531_/X _22532_/X VGND VGND VPWR
+ VPWR _22779_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25567_ _25567_/A VGND VGND VPWR VPWR _33214_/D sky130_fd_sc_hd__clkbuf_1
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27306_ _27306_/A VGND VGND VPWR VPWR _34004_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24518_ _24518_/A VGND VGND VPWR VPWR _32752_/D sky130_fd_sc_hd__clkbuf_1
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28286_ _34468_/Q _24314_/X _28300_/S VGND VGND VPWR VPWR _28287_/A sky130_fd_sc_hd__mux2_1
X_25498_ _25498_/A VGND VGND VPWR VPWR _33181_/D sky130_fd_sc_hd__clkbuf_1
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27237_ _26940_/X _33972_/Q _27239_/S VGND VGND VPWR VPWR _27238_/A sky130_fd_sc_hd__mux2_1
X_24449_ _24449_/A VGND VGND VPWR VPWR _32719_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27168_ _26838_/X _33939_/Q _27176_/S VGND VGND VPWR VPWR _27169_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26119_ _26119_/A VGND VGND VPWR VPWR _33473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19990_ _19986_/X _19989_/X _19781_/X VGND VGND VPWR VPWR _20020_/A sky130_fd_sc_hd__o21ba_1
X_27099_ _27099_/A VGND VGND VPWR VPWR _33906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18941_ _20155_/A VGND VGND VPWR VPWR _18941_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18872_ _32988_/Q _32924_/Q _32860_/Q _32796_/Q _18583_/X _18584_/X VGND VGND VPWR
+ VPWR _18872_/X sky130_fd_sc_hd__mux4_1
XTAP_6650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17823_ _17819_/X _17822_/X _17514_/X VGND VGND VPWR VPWR _17824_/D sky130_fd_sc_hd__o21ba_1
X_29809_ _35159_/Q _29079_/X _29809_/S VGND VGND VPWR VPWR _29810_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32820_ _33013_/CLK _32820_/D VGND VGND VPWR VPWR _32820_/Q sky130_fd_sc_hd__dfxtp_1
X_17754_ _33790_/Q _33726_/Q _33662_/Q _33598_/Q _17549_/X _17550_/X VGND VGND VPWR
+ VPWR _17754_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16705_ _17902_/A VGND VGND VPWR VPWR _16705_/X sky130_fd_sc_hd__buf_4
X_32751_ _36078_/CLK _32751_/D VGND VGND VPWR VPWR _32751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17685_ _34300_/Q _34236_/Q _34172_/Q _34108_/Q _17442_/X _17443_/X VGND VGND VPWR
+ VPWR _17685_/X sky130_fd_sc_hd__mux4_1
X_31702_ _31813_/S VGND VGND VPWR VPWR _31721_/S sky130_fd_sc_hd__buf_6
XFILLER_63_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19424_ _20130_/A VGND VGND VPWR VPWR _19424_/X sky130_fd_sc_hd__buf_4
X_35470_ _35919_/CLK _35470_/D VGND VGND VPWR VPWR _35470_/Q sky130_fd_sc_hd__dfxtp_1
X_16636_ _17829_/A VGND VGND VPWR VPWR _16636_/X sky130_fd_sc_hd__buf_4
XFILLER_223_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32682_ _36139_/CLK _32682_/D VGND VGND VPWR VPWR _32682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34421_ _34805_/CLK _34421_/D VGND VGND VPWR VPWR _34421_/Q sky130_fd_sc_hd__dfxtp_1
X_19355_ _20201_/A VGND VGND VPWR VPWR _19355_/X sky130_fd_sc_hd__buf_4
X_31633_ _36023_/Q input36/X _31649_/S VGND VGND VPWR VPWR _31634_/A sky130_fd_sc_hd__mux2_1
X_16567_ _32732_/Q _32668_/Q _32604_/Q _36060_/Q _16566_/X _16350_/X VGND VGND VPWR
+ VPWR _16567_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18306_ _18359_/A VGND VGND VPWR VPWR _20257_/A sky130_fd_sc_hd__buf_12
XFILLER_200_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34352_ _34866_/CLK _34352_/D VGND VGND VPWR VPWR _34352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31564_ _31564_/A VGND VGND VPWR VPWR _35990_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19286_ _33256_/Q _36136_/Q _33128_/Q _33064_/Q _19005_/X _19006_/X VGND VGND VPWR
+ VPWR _19286_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16498_ _34010_/Q _33946_/Q _33882_/Q _32154_/Q _16314_/X _16315_/X VGND VGND VPWR
+ VPWR _16498_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33303_ _36228_/CLK _33303_/D VGND VGND VPWR VPWR _33303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18237_ _35340_/Q _35276_/Q _35212_/Q _32332_/Q _16088_/X _16090_/X VGND VGND VPWR
+ VPWR _18237_/X sky130_fd_sc_hd__mux4_1
X_30515_ _23199_/X _35493_/Q _30527_/S VGND VGND VPWR VPWR _30516_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34283_ _34283_/CLK _34283_/D VGND VGND VPWR VPWR _34283_/Q sky130_fd_sc_hd__dfxtp_1
X_31495_ _31543_/S VGND VGND VPWR VPWR _31514_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_102_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36022_ _36022_/CLK _36022_/D VGND VGND VPWR VPWR _36022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33234_ _33234_/CLK _33234_/D VGND VGND VPWR VPWR _33234_/Q sky130_fd_sc_hd__dfxtp_1
X_30446_ _30446_/A VGND VGND VPWR VPWR _35460_/D sky130_fd_sc_hd__clkbuf_1
X_18168_ _18164_/X _18167_/X _17842_/A _17843_/A VGND VGND VPWR VPWR _18183_/B sky130_fd_sc_hd__o211a_1
XFILLER_15_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17119_ _17119_/A VGND VGND VPWR VPWR _31979_/D sky130_fd_sc_hd__clkbuf_1
X_33165_ _34316_/CLK _33165_/D VGND VGND VPWR VPWR _33165_/Q sky130_fd_sc_hd__dfxtp_1
X_18099_ _34056_/Q _33992_/Q _33928_/Q _32264_/Q _16058_/X _16060_/X VGND VGND VPWR
+ VPWR _18099_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30377_ _30377_/A VGND VGND VPWR VPWR _35427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20130_ _20130_/A VGND VGND VPWR VPWR _20130_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_132_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32116_ _35555_/CLK _32116_/D VGND VGND VPWR VPWR _32116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33096_ _35909_/CLK _33096_/D VGND VGND VPWR VPWR _33096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20061_ _20061_/A VGND VGND VPWR VPWR _20061_/X sky130_fd_sc_hd__clkbuf_4
X_32047_ _36013_/CLK _32047_/D VGND VGND VPWR VPWR _32047_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23820_ _23053_/X _32454_/Q _23826_/S VGND VGND VPWR VPWR _23821_/A sky130_fd_sc_hd__mux2_1
X_35806_ _35809_/CLK _35806_/D VGND VGND VPWR VPWR _35806_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33998_ _35792_/CLK _33998_/D VGND VGND VPWR VPWR _33998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23751_ _22951_/X _32421_/Q _23763_/S VGND VGND VPWR VPWR _23752_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_309 _32140_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20963_ _20956_/X _20962_/X _20640_/X _20642_/X VGND VGND VPWR VPWR _20980_/B sky130_fd_sc_hd__o211a_1
X_35737_ _35929_/CLK _35737_/D VGND VGND VPWR VPWR _35737_/Q sky130_fd_sc_hd__dfxtp_1
X_32949_ _35829_/CLK _32949_/D VGND VGND VPWR VPWR _32949_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22702_ _32776_/Q _32712_/Q _32648_/Q _36104_/Q _22578_/X _21473_/A VGND VGND VPWR
+ VPWR _22702_/X sky130_fd_sc_hd__mux4_1
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23682_ _32390_/Q _23322_/X _23688_/S VGND VGND VPWR VPWR _23683_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26470_ _25072_/X _33640_/Q _26476_/S VGND VGND VPWR VPWR _26471_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20894_ _35540_/Q _35476_/Q _35412_/Q _35348_/Q _20791_/X _20792_/X VGND VGND VPWR
+ VPWR _20894_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35668_ _35669_/CLK _35668_/D VGND VGND VPWR VPWR _35668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22633_ _22633_/A _22633_/B _22633_/C _22633_/D VGND VGND VPWR VPWR _22634_/A sky130_fd_sc_hd__or4_4
X_25421_ _25131_/X _33147_/Q _25429_/S VGND VGND VPWR VPWR _25422_/A sky130_fd_sc_hd__mux2_1
X_34619_ _35707_/CLK _34619_/D VGND VGND VPWR VPWR _34619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_1070 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35599_ _35792_/CLK _35599_/D VGND VGND VPWR VPWR _35599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28140_ _26875_/X _34399_/Q _28144_/S VGND VGND VPWR VPWR _28141_/A sky130_fd_sc_hd__mux2_1
X_25352_ _25029_/X _33114_/Q _25366_/S VGND VGND VPWR VPWR _25353_/A sky130_fd_sc_hd__mux2_1
X_22564_ _22455_/X _22562_/X _22563_/X _22458_/X VGND VGND VPWR VPWR _22564_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21515_ _33510_/Q _33446_/Q _33382_/Q _33318_/Q _21370_/X _21371_/X VGND VGND VPWR
+ VPWR _21515_/X sky130_fd_sc_hd__mux4_1
X_24303_ _24303_/A VGND VGND VPWR VPWR _32672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28071_ _28071_/A VGND VGND VPWR VPWR _34366_/D sky130_fd_sc_hd__clkbuf_1
X_25283_ _25128_/X _33082_/Q _25293_/S VGND VGND VPWR VPWR _25284_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22495_ _34561_/Q _32449_/Q _34433_/Q _34369_/Q _22178_/X _22179_/X VGND VGND VPWR
+ VPWR _22495_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27022_ _27154_/S VGND VGND VPWR VPWR _27041_/S sky130_fd_sc_hd__buf_4
X_24234_ _23062_/X _32649_/Q _24234_/S VGND VGND VPWR VPWR _24235_/A sky130_fd_sc_hd__mux2_1
X_21446_ _34276_/Q _34212_/Q _34148_/Q _34084_/Q _21336_/X _21337_/X VGND VGND VPWR
+ VPWR _21446_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24165_ _22960_/X _32616_/Q _24171_/S VGND VGND VPWR VPWR _24166_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21377_ _32738_/Q _32674_/Q _32610_/Q _36066_/Q _21166_/X _21303_/X VGND VGND VPWR
+ VPWR _21377_/X sky130_fd_sc_hd__mux4_1
X_23116_ _23116_/A VGND VGND VPWR VPWR _32151_/D sky130_fd_sc_hd__clkbuf_1
X_20328_ _20155_/X _20326_/X _20327_/X _20158_/X VGND VGND VPWR VPWR _20328_/X sky130_fd_sc_hd__a22o_1
XFILLER_218_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24096_ _23059_/X _32584_/Q _24098_/S VGND VGND VPWR VPWR _24097_/A sky130_fd_sc_hd__mux2_1
X_28973_ _34794_/Q _24332_/X _28975_/S VGND VGND VPWR VPWR _28974_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23047_ input50/X VGND VGND VPWR VPWR _23047_/X sky130_fd_sc_hd__buf_4
XFILLER_122_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27924_ _27924_/A VGND VGND VPWR VPWR _34296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20259_ _33219_/Q _32579_/Q _35971_/Q _35907_/Q _20080_/X _20081_/X VGND VGND VPWR
+ VPWR _20259_/X sky130_fd_sc_hd__mux4_1
XTAP_5201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27855_ _27966_/S VGND VGND VPWR VPWR _27874_/S sky130_fd_sc_hd__buf_4
XTAP_5256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_1__f_CLK clkbuf_5_0_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_9_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_95_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26806_ _26806_/A VGND VGND VPWR VPWR _33798_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27786_ _34231_/Q _24373_/X _27802_/S VGND VGND VPWR VPWR _27787_/A sky130_fd_sc_hd__mux2_1
X_24998_ input23/X VGND VGND VPWR VPWR _24998_/X sky130_fd_sc_hd__buf_4
XTAP_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29525_ _35024_/Q _29058_/X _29539_/S VGND VGND VPWR VPWR _29526_/A sky130_fd_sc_hd__mux2_1
XTAP_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26737_ _26737_/A VGND VGND VPWR VPWR _33765_/D sky130_fd_sc_hd__clkbuf_1
X_23949_ _23949_/A VGND VGND VPWR VPWR _32514_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_923 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_810 _22907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_821 _23421_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29456_ _29456_/A VGND VGND VPWR VPWR _34991_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17470_ _17466_/X _17469_/X _17161_/X VGND VGND VPWR VPWR _17471_/D sky130_fd_sc_hd__o21ba_1
XANTENNA_832 _23133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26668_ _26668_/A VGND VGND VPWR VPWR _33733_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_843 _23333_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_854 _24301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_865 _24425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16421_ _16143_/X _16419_/X _16420_/X _16146_/X VGND VGND VPWR VPWR _16421_/X sky130_fd_sc_hd__a22o_1
X_28407_ _28407_/A VGND VGND VPWR VPWR _34525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25619_ _25619_/A VGND VGND VPWR VPWR _33237_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_876 _25187_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29387_ _29387_/A VGND VGND VPWR VPWR _34958_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_887 _25322_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_898 _26007_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26599_ _26599_/A VGND VGND VPWR VPWR _33700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19140_ _19140_/A _19140_/B _19140_/C _19140_/D VGND VGND VPWR VPWR _19141_/A sky130_fd_sc_hd__or4_2
X_28338_ _34493_/Q _24391_/X _28342_/S VGND VGND VPWR VPWR _28339_/A sky130_fd_sc_hd__mux2_1
X_16352_ _17902_/A VGND VGND VPWR VPWR _16352_/X sky130_fd_sc_hd__buf_4
XFILLER_73_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19071_ _20130_/A VGND VGND VPWR VPWR _19071_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_40_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16283_ _17829_/A VGND VGND VPWR VPWR _16283_/X sky130_fd_sc_hd__buf_4
X_28269_ _34460_/Q _24289_/X _28279_/S VGND VGND VPWR VPWR _28270_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30300_ _30327_/S VGND VGND VPWR VPWR _30319_/S sky130_fd_sc_hd__buf_4
X_18022_ _35589_/Q _35525_/Q _35461_/Q _35397_/Q _17956_/X _17957_/X VGND VGND VPWR
+ VPWR _18022_/X sky130_fd_sc_hd__mux4_1
X_31280_ _31280_/A VGND VGND VPWR VPWR _35855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30231_ _35359_/Q _29104_/X _30235_/S VGND VGND VPWR VPWR _30232_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30162_ _30162_/A VGND VGND VPWR VPWR _35326_/D sky130_fd_sc_hd__clkbuf_1
X_19973_ _19652_/X _19971_/X _19972_/X _19655_/X VGND VGND VPWR VPWR _19973_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18924_ _18924_/A VGND VGND VPWR VPWR _32093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1220 _24273_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_34970_ _34970_/CLK _34970_/D VGND VGND VPWR VPWR _34970_/Q sky130_fd_sc_hd__dfxtp_1
X_30093_ _30093_/A VGND VGND VPWR VPWR _35293_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1231 _24416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1242 _25872_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33921_ _36165_/CLK _33921_/D VGND VGND VPWR VPWR _33921_/Q sky130_fd_sc_hd__dfxtp_1
X_18855_ _18748_/X _18853_/X _18854_/X _18753_/X VGND VGND VPWR VPWR _18855_/X sky130_fd_sc_hd__a22o_1
XANTENNA_1253 _26863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1264 _29213_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1275 _31813_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17806_ _32511_/Q _32383_/Q _32063_/Q _36031_/Q _17629_/X _17770_/X VGND VGND VPWR
+ VPWR _17806_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1286 _17858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33852_ _35772_/CLK _33852_/D VGND VGND VPWR VPWR _33852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1297 _17157_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18786_ _18782_/X _18785_/X _18755_/X VGND VGND VPWR VPWR _18787_/D sky130_fd_sc_hd__o21ba_1
X_15998_ _17795_/A VGND VGND VPWR VPWR _15998_/X sky130_fd_sc_hd__buf_4
XFILLER_212_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32803_ _32994_/CLK _32803_/D VGND VGND VPWR VPWR _32803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17737_ _17733_/X _17736_/X _17489_/X _17490_/X VGND VGND VPWR VPWR _17752_/B sky130_fd_sc_hd__o211a_1
XFILLER_208_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33783_ _34039_/CLK _33783_/D VGND VGND VPWR VPWR _33783_/Q sky130_fd_sc_hd__dfxtp_1
X_30995_ _35721_/Q _29234_/X _30995_/S VGND VGND VPWR VPWR _30996_/A sky130_fd_sc_hd__mux2_1
X_35522_ _35585_/CLK _35522_/D VGND VGND VPWR VPWR _35522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32734_ _36062_/CLK _32734_/D VGND VGND VPWR VPWR _32734_/Q sky130_fd_sc_hd__dfxtp_1
X_17668_ _35835_/Q _32213_/Q _35707_/Q _35643_/Q _17666_/X _17667_/X VGND VGND VPWR
+ VPWR _17668_/X sky130_fd_sc_hd__mux4_1
XFILLER_247_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19407_ _35563_/Q _35499_/Q _35435_/Q _35371_/Q _19197_/X _19198_/X VGND VGND VPWR
+ VPWR _19407_/X sky130_fd_sc_hd__mux4_1
X_35453_ _35517_/CLK _35453_/D VGND VGND VPWR VPWR _35453_/Q sky130_fd_sc_hd__dfxtp_1
X_16619_ _34525_/Q _32413_/Q _34397_/Q _34333_/Q _16519_/X _16520_/X VGND VGND VPWR
+ VPWR _16619_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32665_ _35799_/CLK _32665_/D VGND VGND VPWR VPWR _32665_/Q sky130_fd_sc_hd__dfxtp_1
X_17599_ _17595_/X _17598_/X _17489_/X _17490_/X VGND VGND VPWR VPWR _17616_/B sky130_fd_sc_hd__o211a_1
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34404_ _35042_/CLK _34404_/D VGND VGND VPWR VPWR _34404_/Q sky130_fd_sc_hd__dfxtp_1
X_19338_ _19334_/X _19337_/X _19094_/X VGND VGND VPWR VPWR _19346_/C sky130_fd_sc_hd__o21ba_1
X_31616_ _36015_/Q input27/X _31628_/S VGND VGND VPWR VPWR _31617_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35384_ _35638_/CLK _35384_/D VGND VGND VPWR VPWR _35384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32596_ _36116_/CLK _32596_/D VGND VGND VPWR VPWR _32596_/Q sky130_fd_sc_hd__dfxtp_1
X_34335_ _35039_/CLK _34335_/D VGND VGND VPWR VPWR _34335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31547_ _35982_/Q input1/X _31565_/S VGND VGND VPWR VPWR _31548_/A sky130_fd_sc_hd__mux2_1
X_19269_ _34791_/Q _34727_/Q _34663_/Q _34599_/Q _19235_/X _19236_/X VGND VGND VPWR
+ VPWR _19269_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21300_ _21096_/X _21298_/X _21299_/X _21099_/X VGND VGND VPWR VPWR _21300_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22280_ _22107_/X _22278_/X _22279_/X _22112_/X VGND VGND VPWR VPWR _22280_/X sky130_fd_sc_hd__a22o_1
XFILLER_129_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34266_ _34266_/CLK _34266_/D VGND VGND VPWR VPWR _34266_/Q sky130_fd_sc_hd__dfxtp_1
X_31478_ _31478_/A VGND VGND VPWR VPWR _35949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36005_ _36005_/CLK _36005_/D VGND VGND VPWR VPWR _36005_/Q sky130_fd_sc_hd__dfxtp_1
X_33217_ _35906_/CLK _33217_/D VGND VGND VPWR VPWR _33217_/Q sky130_fd_sc_hd__dfxtp_1
X_21231_ _21227_/X _21230_/X _21022_/X VGND VGND VPWR VPWR _21261_/A sky130_fd_sc_hd__o21ba_1
X_30429_ _30429_/A VGND VGND VPWR VPWR _35452_/D sky130_fd_sc_hd__clkbuf_1
X_34197_ _34197_/CLK _34197_/D VGND VGND VPWR VPWR _34197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33148_ _36095_/CLK _33148_/D VGND VGND VPWR VPWR _33148_/Q sky130_fd_sc_hd__dfxtp_1
X_21162_ _33500_/Q _33436_/Q _33372_/Q _33308_/Q _21017_/X _21018_/X VGND VGND VPWR
+ VPWR _21162_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20113_ _35583_/Q _35519_/Q _35455_/Q _35391_/Q _19903_/X _19904_/X VGND VGND VPWR
+ VPWR _20113_/X sky130_fd_sc_hd__mux4_1
XFILLER_160_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25970_ _25131_/X _33403_/Q _25978_/S VGND VGND VPWR VPWR _25971_/A sky130_fd_sc_hd__mux2_1
X_33079_ _36088_/CLK _33079_/D VGND VGND VPWR VPWR _33079_/Q sky130_fd_sc_hd__dfxtp_1
X_21093_ _34266_/Q _34202_/Q _34138_/Q _34074_/Q _20983_/X _20984_/X VGND VGND VPWR
+ VPWR _21093_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_860 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20044_ _20040_/X _20043_/X _19800_/X VGND VGND VPWR VPWR _20052_/C sky130_fd_sc_hd__o21ba_1
X_24921_ _22976_/X _32941_/Q _24937_/S VGND VGND VPWR VPWR _24922_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27640_ _34162_/Q _24357_/X _27646_/S VGND VGND VPWR VPWR _27641_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24852_ _23074_/X _32909_/Q _24852_/S VGND VGND VPWR VPWR _24853_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_1479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_928 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23803_ _23028_/X _32446_/Q _23805_/S VGND VGND VPWR VPWR _23804_/A sky130_fd_sc_hd__mux2_1
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27571_ _34129_/Q _24255_/X _27583_/S VGND VGND VPWR VPWR _27572_/A sky130_fd_sc_hd__mux2_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ _34547_/Q _32435_/Q _34419_/Q _34355_/Q _21825_/X _21826_/X VGND VGND VPWR
+ VPWR _21995_/X sky130_fd_sc_hd__mux4_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24783_ _24852_/S VGND VGND VPWR VPWR _24802_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_227_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_106 _32129_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_117 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29310_ _29310_/A VGND VGND VPWR VPWR _34922_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26522_ _26522_/A VGND VGND VPWR VPWR _33664_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_128 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20946_ _34006_/Q _33942_/Q _33878_/Q _32150_/Q _20914_/X _20915_/X VGND VGND VPWR
+ VPWR _20946_/X sky130_fd_sc_hd__mux4_1
XANTENNA_139 _32132_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23734_ _22926_/X _32413_/Q _23742_/S VGND VGND VPWR VPWR _23735_/A sky130_fd_sc_hd__mux2_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29241_ _34891_/Q _29240_/X _29247_/S VGND VGND VPWR VPWR _29242_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26453_ _25047_/X _33632_/Q _26455_/S VGND VGND VPWR VPWR _26454_/A sky130_fd_sc_hd__mux2_1
X_20877_ _20743_/X _20875_/X _20876_/X _20746_/X VGND VGND VPWR VPWR _20877_/X sky130_fd_sc_hd__a22o_1
XFILLER_214_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23665_ _32382_/Q _23297_/X _23667_/S VGND VGND VPWR VPWR _23666_/A sky130_fd_sc_hd__mux2_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25404_ _25106_/X _33139_/Q _25408_/S VGND VGND VPWR VPWR _25405_/A sky130_fd_sc_hd__mux2_1
X_22616_ _33029_/Q _32965_/Q _32901_/Q _32837_/Q _22295_/X _22296_/X VGND VGND VPWR
+ VPWR _22616_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29172_ input33/X VGND VGND VPWR VPWR _29172_/X sky130_fd_sc_hd__clkbuf_4
X_26384_ _26384_/A VGND VGND VPWR VPWR _33599_/D sky130_fd_sc_hd__clkbuf_1
X_23596_ _32349_/Q _23133_/X _23604_/S VGND VGND VPWR VPWR _23597_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28123_ _26850_/X _34391_/Q _28123_/S VGND VGND VPWR VPWR _28124_/A sky130_fd_sc_hd__mux2_1
X_22547_ _33283_/Q _36163_/Q _33155_/Q _33091_/Q _22364_/X _22365_/X VGND VGND VPWR
+ VPWR _22547_/X sky130_fd_sc_hd__mux4_1
X_25335_ _25004_/X _33106_/Q _25345_/S VGND VGND VPWR VPWR _25336_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28054_ _26946_/X _34358_/Q _28072_/S VGND VGND VPWR VPWR _28055_/A sky130_fd_sc_hd__mux2_1
X_22478_ _32769_/Q _32705_/Q _32641_/Q _36097_/Q _22225_/X _22362_/X VGND VGND VPWR
+ VPWR _22478_/X sky130_fd_sc_hd__mux4_1
X_25266_ _25103_/X _33074_/Q _25272_/S VGND VGND VPWR VPWR _25267_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27005_ input55/X VGND VGND VPWR VPWR _27005_/X sky130_fd_sc_hd__buf_4
XFILLER_202_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24217_ _24217_/A VGND VGND VPWR VPWR _32640_/D sky130_fd_sc_hd__clkbuf_1
X_21429_ _35555_/Q _35491_/Q _35427_/Q _35363_/Q _21144_/X _21145_/X VGND VGND VPWR
+ VPWR _21429_/X sky130_fd_sc_hd__mux4_1
X_25197_ _25001_/X _33041_/Q _25209_/S VGND VGND VPWR VPWR _25198_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24148_ _22935_/X _32608_/Q _24150_/S VGND VGND VPWR VPWR _24149_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24079_ _24106_/S VGND VGND VPWR VPWR _24098_/S sky130_fd_sc_hd__buf_4
X_16970_ _35303_/Q _35239_/Q _35175_/Q _32295_/Q _16653_/X _16654_/X VGND VGND VPWR
+ VPWR _16970_/X sky130_fd_sc_hd__mux4_1
X_28956_ _28998_/A VGND VGND VPWR VPWR _28975_/S sky130_fd_sc_hd__buf_4
XFILLER_110_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27907_ _27907_/A VGND VGND VPWR VPWR _34288_/D sky130_fd_sc_hd__clkbuf_1
X_28887_ _26981_/X _34753_/Q _28903_/S VGND VGND VPWR VPWR _28888_/A sky130_fd_sc_hd__mux2_1
XTAP_5031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18640_ _18640_/A _18640_/B _18640_/C _18640_/D VGND VGND VPWR VPWR _18641_/A sky130_fd_sc_hd__or4_4
X_27838_ _27838_/A VGND VGND VPWR VPWR _34255_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ _18571_/A VGND VGND VPWR VPWR _32083_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27769_ _34223_/Q _24348_/X _27781_/S VGND VGND VPWR VPWR _27770_/A sky130_fd_sc_hd__mux2_1
XTAP_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29508_ _29508_/A VGND VGND VPWR VPWR _35016_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ _34039_/Q _33975_/Q _33911_/Q _32247_/Q _17373_/X _17374_/X VGND VGND VPWR
+ VPWR _17522_/X sky130_fd_sc_hd__mux4_1
XTAP_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30780_ _30780_/A VGND VGND VPWR VPWR _35618_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_640 _19347_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_651 _20208_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_662 _22455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29439_ _29439_/A VGND VGND VPWR VPWR _34983_/D sky130_fd_sc_hd__clkbuf_1
X_17453_ _32501_/Q _32373_/Q _32053_/Q _36021_/Q _17276_/X _17417_/X VGND VGND VPWR
+ VPWR _17453_/X sky130_fd_sc_hd__mux4_1
XANTENNA_673 _22460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_684 _22434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_695 _22595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16404_ _16400_/X _16403_/X _16071_/X VGND VGND VPWR VPWR _16412_/C sky130_fd_sc_hd__o21ba_1
X_32450_ _35330_/CLK _32450_/D VGND VGND VPWR VPWR _32450_/Q sky130_fd_sc_hd__dfxtp_1
X_17384_ _17380_/X _17383_/X _17136_/X _17137_/X VGND VGND VPWR VPWR _17399_/B sky130_fd_sc_hd__o211a_1
XFILLER_198_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31401_ _31401_/A VGND VGND VPWR VPWR _35913_/D sky130_fd_sc_hd__clkbuf_1
X_19123_ _32995_/Q _32931_/Q _32867_/Q _32803_/Q _18936_/X _18937_/X VGND VGND VPWR
+ VPWR _19123_/X sky130_fd_sc_hd__mux4_1
X_16335_ _16074_/X _16333_/X _16334_/X _16084_/X VGND VGND VPWR VPWR _16335_/X sky130_fd_sc_hd__a22o_1
X_32381_ _36029_/CLK _32381_/D VGND VGND VPWR VPWR _32381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34120_ _34819_/CLK _34120_/D VGND VGND VPWR VPWR _34120_/Q sky130_fd_sc_hd__dfxtp_1
X_19054_ _35553_/Q _35489_/Q _35425_/Q _35361_/Q _18844_/X _18845_/X VGND VGND VPWR
+ VPWR _19054_/X sky130_fd_sc_hd__mux4_1
X_31332_ _31332_/A VGND VGND VPWR VPWR _35880_/D sky130_fd_sc_hd__clkbuf_1
X_16266_ _34515_/Q _32403_/Q _34387_/Q _34323_/Q _16166_/X _16167_/X VGND VGND VPWR
+ VPWR _16266_/X sky130_fd_sc_hd__mux4_1
XFILLER_199_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_930 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18005_ _33797_/Q _33733_/Q _33669_/Q _33605_/Q _17902_/X _17903_/X VGND VGND VPWR
+ VPWR _18005_/X sky130_fd_sc_hd__mux4_1
X_34051_ _34053_/CLK _34051_/D VGND VGND VPWR VPWR _34051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31263_ _35848_/Q input54/X _31265_/S VGND VGND VPWR VPWR _31264_/A sky130_fd_sc_hd__mux2_1
X_16197_ _34769_/Q _34705_/Q _34641_/Q _34577_/Q _16075_/X _16076_/X VGND VGND VPWR
+ VPWR _16197_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33002_ _36137_/CLK _33002_/D VGND VGND VPWR VPWR _33002_/Q sky130_fd_sc_hd__dfxtp_1
X_30214_ _35351_/Q _29079_/X _30214_/S VGND VGND VPWR VPWR _30215_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31194_ _35815_/Q input18/X _31202_/S VGND VGND VPWR VPWR _31195_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30145_ _35318_/Q _29175_/X _30163_/S VGND VGND VPWR VPWR _30146_/A sky130_fd_sc_hd__mux2_1
X_19956_ _34043_/Q _33979_/Q _33915_/Q _32251_/Q _19673_/X _19674_/X VGND VGND VPWR
+ VPWR _19956_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18907_ _20095_/A VGND VGND VPWR VPWR _18907_/X sky130_fd_sc_hd__buf_4
XANTENNA_1050 _17867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_34953_ _35784_/CLK _34953_/D VGND VGND VPWR VPWR _34953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30076_ _30076_/A VGND VGND VPWR VPWR _35285_/D sky130_fd_sc_hd__clkbuf_1
X_19887_ _34297_/Q _34233_/Q _34169_/Q _34105_/Q _19742_/X _19743_/X VGND VGND VPWR
+ VPWR _19887_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1061 _16733_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1072 _17164_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1083 _17232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33904_ _34032_/CLK _33904_/D VGND VGND VPWR VPWR _33904_/Q sky130_fd_sc_hd__dfxtp_1
X_18838_ _32987_/Q _32923_/Q _32859_/Q _32795_/Q _18583_/X _18584_/X VGND VGND VPWR
+ VPWR _18838_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1094 _17264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_34884_ _35779_/CLK _34884_/D VGND VGND VPWR VPWR _34884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18769_ _32473_/Q _32345_/Q _32025_/Q _35993_/Q _18517_/X _18658_/X VGND VGND VPWR
+ VPWR _18769_/X sky130_fd_sc_hd__mux4_1
X_33835_ _35944_/CLK _33835_/D VGND VGND VPWR VPWR _33835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20800_ _34513_/Q _32401_/Q _34385_/Q _34321_/Q _20766_/X _20767_/X VGND VGND VPWR
+ VPWR _20800_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33766_ _34278_/CLK _33766_/D VGND VGND VPWR VPWR _33766_/Q sky130_fd_sc_hd__dfxtp_1
X_21780_ _35757_/Q _35117_/Q _34477_/Q _33837_/Q _21740_/X _21741_/X VGND VGND VPWR
+ VPWR _21780_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30978_ _30978_/A VGND VGND VPWR VPWR _35712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20731_ _35023_/Q _34959_/Q _34895_/Q _34831_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _20731_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35505_ _35889_/CLK _35505_/D VGND VGND VPWR VPWR _35505_/Q sky130_fd_sc_hd__dfxtp_1
X_32717_ _36173_/CLK _32717_/D VGND VGND VPWR VPWR _32717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33697_ _34145_/CLK _33697_/D VGND VGND VPWR VPWR _33697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23450_ _23450_/A VGND VGND VPWR VPWR _32280_/D sky130_fd_sc_hd__clkbuf_1
X_32648_ _36169_/CLK _32648_/D VGND VGND VPWR VPWR _32648_/Q sky130_fd_sc_hd__dfxtp_1
X_35436_ _35562_/CLK _35436_/D VGND VGND VPWR VPWR _35436_/Q sky130_fd_sc_hd__dfxtp_1
X_20662_ _22578_/A VGND VGND VPWR VPWR _22531_/A sky130_fd_sc_hd__buf_12
XFILLER_23_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22401_ _22155_/X _22399_/X _22400_/X _22158_/X VGND VGND VPWR VPWR _22401_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23381_ _23381_/A VGND VGND VPWR VPWR _32249_/D sky130_fd_sc_hd__clkbuf_1
X_20593_ _20577_/X _20584_/X _20587_/X _20592_/X VGND VGND VPWR VPWR _20593_/X sky130_fd_sc_hd__a22o_1
XFILLER_220_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32579_ _36037_/CLK _32579_/D VGND VGND VPWR VPWR _32579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35367_ _35750_/CLK _35367_/D VGND VGND VPWR VPWR _35367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22332_ _33277_/Q _36157_/Q _33149_/Q _33085_/Q _22011_/X _22012_/X VGND VGND VPWR
+ VPWR _22332_/X sky130_fd_sc_hd__mux4_1
X_25120_ _25119_/X _33015_/Q _25144_/S VGND VGND VPWR VPWR _25121_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34318_ _34638_/CLK _34318_/D VGND VGND VPWR VPWR _34318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35298_ _35298_/CLK _35298_/D VGND VGND VPWR VPWR _35298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25051_ _25050_/X _32993_/Q _25051_/S VGND VGND VPWR VPWR _25052_/A sky130_fd_sc_hd__mux2_1
X_34249_ _34816_/CLK _34249_/D VGND VGND VPWR VPWR _34249_/Q sky130_fd_sc_hd__dfxtp_1
X_22263_ _33019_/Q _32955_/Q _32891_/Q _32827_/Q _21942_/X _21943_/X VGND VGND VPWR
+ VPWR _22263_/X sky130_fd_sc_hd__mux4_1
X_24002_ _22920_/X _32539_/Q _24014_/S VGND VGND VPWR VPWR _24003_/A sky130_fd_sc_hd__mux2_1
X_21214_ _20893_/X _21212_/X _21213_/X _20896_/X VGND VGND VPWR VPWR _21214_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22194_ _33273_/Q _36153_/Q _33145_/Q _33081_/Q _22011_/X _22012_/X VGND VGND VPWR
+ VPWR _22194_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28810_ _28810_/A VGND VGND VPWR VPWR _34716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21145_ _22557_/A VGND VGND VPWR VPWR _21145_/X sky130_fd_sc_hd__clkbuf_4
X_29790_ _29922_/S VGND VGND VPWR VPWR _29809_/S sky130_fd_sc_hd__buf_6
XFILLER_116_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_14__f_CLK clkbuf_5_7_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_14__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_28741_ _26965_/X _34684_/Q _28747_/S VGND VGND VPWR VPWR _28742_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21076_ _35545_/Q _35481_/Q _35417_/Q _35353_/Q _20791_/X _20792_/X VGND VGND VPWR
+ VPWR _21076_/X sky130_fd_sc_hd__mux4_1
X_25953_ _25106_/X _33395_/Q _25957_/S VGND VGND VPWR VPWR _25954_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20027_ _20147_/A VGND VGND VPWR VPWR _20027_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_189_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24904_ _22951_/X _32933_/Q _24916_/S VGND VGND VPWR VPWR _24905_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28672_ _26863_/X _34651_/Q _28684_/S VGND VGND VPWR VPWR _28673_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25884_ _25004_/X _33362_/Q _25894_/S VGND VGND VPWR VPWR _25885_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27623_ _34154_/Q _24332_/X _27625_/S VGND VGND VPWR VPWR _27624_/A sky130_fd_sc_hd__mux2_1
X_24835_ _24835_/A VGND VGND VPWR VPWR _32900_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27554_ _27554_/A VGND VGND VPWR VPWR _34122_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24766_ _24766_/A VGND VGND VPWR VPWR _32867_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21978_ _32755_/Q _32691_/Q _32627_/Q _36083_/Q _21872_/X _21656_/X VGND VGND VPWR
+ VPWR _21978_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26505_ _26505_/A VGND VGND VPWR VPWR _33656_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23717_ _22901_/X _32405_/Q _23721_/S VGND VGND VPWR VPWR _23718_/A sky130_fd_sc_hd__mux2_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20929_ _35541_/Q _35477_/Q _35413_/Q _35349_/Q _20791_/X _20792_/X VGND VGND VPWR
+ VPWR _20929_/X sky130_fd_sc_hd__mux4_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27485_ _27485_/A VGND VGND VPWR VPWR _34089_/D sky130_fd_sc_hd__clkbuf_1
X_24697_ _23047_/X _32836_/Q _24707_/S VGND VGND VPWR VPWR _24698_/A sky130_fd_sc_hd__mux2_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29224_ _29224_/A VGND VGND VPWR VPWR _34885_/D sky130_fd_sc_hd__clkbuf_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26436_ _26547_/S VGND VGND VPWR VPWR _26455_/S sky130_fd_sc_hd__buf_4
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23648_ _23696_/S VGND VGND VPWR VPWR _23667_/S sky130_fd_sc_hd__buf_4
XFILLER_109_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29155_ _34863_/Q _29154_/X _29173_/S VGND VGND VPWR VPWR _29156_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_195_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _35585_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26367_ _25119_/X _33591_/Q _26383_/S VGND VGND VPWR VPWR _26368_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23579_ _32341_/Q _23108_/X _23583_/S VGND VGND VPWR VPWR _23580_/A sky130_fd_sc_hd__mux2_1
X_16120_ _35791_/Q _32165_/Q _35663_/Q _35599_/Q _16045_/X _16046_/X VGND VGND VPWR
+ VPWR _16120_/X sky130_fd_sc_hd__mux4_1
X_28106_ _28106_/A VGND VGND VPWR VPWR _34382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25318_ _25180_/X _33099_/Q _25322_/S VGND VGND VPWR VPWR _25319_/A sky130_fd_sc_hd__mux2_1
X_29086_ input3/X VGND VGND VPWR VPWR _29086_/X sky130_fd_sc_hd__clkbuf_4
X_26298_ _26298_/A VGND VGND VPWR VPWR _33558_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16051_ _17995_/A VGND VGND VPWR VPWR _16051_/X sky130_fd_sc_hd__clkbuf_4
X_28037_ _26922_/X _34350_/Q _28051_/S VGND VGND VPWR VPWR _28038_/A sky130_fd_sc_hd__mux2_1
X_25249_ _25078_/X _33066_/Q _25251_/S VGND VGND VPWR VPWR _25250_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19810_ _20163_/A VGND VGND VPWR VPWR _19810_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_124_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29988_ _30057_/S VGND VGND VPWR VPWR _30007_/S sky130_fd_sc_hd__buf_4
XFILLER_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16953_ _32743_/Q _32679_/Q _32615_/Q _36071_/Q _16919_/X _16703_/X VGND VGND VPWR
+ VPWR _16953_/X sky130_fd_sc_hd__mux4_1
X_19741_ _33781_/Q _33717_/Q _33653_/Q _33589_/Q _19496_/X _19497_/X VGND VGND VPWR
+ VPWR _19741_/X sky130_fd_sc_hd__mux4_1
X_28939_ _28939_/A VGND VGND VPWR VPWR _34777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31950_ _34973_/CLK _31950_/D VGND VGND VPWR VPWR _31950_/Q sky130_fd_sc_hd__dfxtp_1
X_19672_ _33523_/Q _33459_/Q _33395_/Q _33331_/Q _19423_/X _19424_/X VGND VGND VPWR
+ VPWR _19672_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16884_ _34021_/Q _33957_/Q _33893_/Q _32182_/Q _16667_/X _16668_/X VGND VGND VPWR
+ VPWR _16884_/X sky130_fd_sc_hd__mux4_1
X_18623_ _32981_/Q _32917_/Q _32853_/Q _32789_/Q _18583_/X _18584_/X VGND VGND VPWR
+ VPWR _18623_/X sky130_fd_sc_hd__mux4_1
X_30901_ _35676_/Q _29095_/X _30911_/S VGND VGND VPWR VPWR _30902_/A sky130_fd_sc_hd__mux2_1
XTAP_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31881_ _31881_/A VGND VGND VPWR VPWR _36140_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33620_ _33685_/CLK _33620_/D VGND VGND VPWR VPWR _33620_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30832_ _30832_/A VGND VGND VPWR VPWR _35643_/D sky130_fd_sc_hd__clkbuf_1
X_18554_ _20095_/A VGND VGND VPWR VPWR _18554_/X sky130_fd_sc_hd__buf_6
XFILLER_18_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17505_ _17858_/A VGND VGND VPWR VPWR _17505_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33551_ _35341_/CLK _33551_/D VGND VGND VPWR VPWR _33551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18485_ _32977_/Q _32913_/Q _32849_/Q _32785_/Q _18333_/X _18335_/X VGND VGND VPWR
+ VPWR _18485_/X sky130_fd_sc_hd__mux4_1
X_30763_ _30763_/A VGND VGND VPWR VPWR _35610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_470 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_481 _31993_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32502_ _36022_/CLK _32502_/D VGND VGND VPWR VPWR _32502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17436_ _35060_/Q _34996_/Q _34932_/Q _34868_/Q _17156_/X _17157_/X VGND VGND VPWR
+ VPWR _17436_/X sky130_fd_sc_hd__mux4_1
XANTENNA_492 _31994_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33482_ _36107_/CLK _33482_/D VGND VGND VPWR VPWR _33482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30694_ _35578_/Q _29188_/X _30704_/S VGND VGND VPWR VPWR _30695_/A sky130_fd_sc_hd__mux2_1
XANTENNA_17 _32115_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35221_ _36202_/CLK _35221_/D VGND VGND VPWR VPWR _35221_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_28 _32116_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32433_ _34866_/CLK _32433_/D VGND VGND VPWR VPWR _32433_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_186_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _35386_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_39 _32117_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17367_ _17367_/A _17367_/B _17367_/C _17367_/D VGND VGND VPWR VPWR _17368_/A sky130_fd_sc_hd__or4_4
XFILLER_53_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19106_ _19459_/A VGND VGND VPWR VPWR _19106_/X sky130_fd_sc_hd__buf_4
XFILLER_105_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16318_ _16312_/X _16317_/X _16011_/X VGND VGND VPWR VPWR _16340_/A sky130_fd_sc_hd__o21ba_1
X_35152_ _35280_/CLK _35152_/D VGND VGND VPWR VPWR _35152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32364_ _36013_/CLK _32364_/D VGND VGND VPWR VPWR _32364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17298_ _17298_/A VGND VGND VPWR VPWR _31984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34103_ _36150_/CLK _34103_/D VGND VGND VPWR VPWR _34103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31315_ _31315_/A VGND VGND VPWR VPWR _35872_/D sky130_fd_sc_hd__clkbuf_1
X_19037_ _20257_/A VGND VGND VPWR VPWR _19037_/X sky130_fd_sc_hd__buf_4
X_35083_ _35338_/CLK _35083_/D VGND VGND VPWR VPWR _35083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16249_ _16014_/X _16247_/X _16248_/X _16023_/X VGND VGND VPWR VPWR _16249_/X sky130_fd_sc_hd__a22o_1
X_32295_ _36005_/CLK _32295_/D VGND VGND VPWR VPWR _32295_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput102 _31970_/Q VGND VGND VPWR VPWR D1[20] sky130_fd_sc_hd__buf_2
X_34034_ _34288_/CLK _34034_/D VGND VGND VPWR VPWR _34034_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput113 _31980_/Q VGND VGND VPWR VPWR D1[30] sky130_fd_sc_hd__buf_2
X_31246_ _31273_/S VGND VGND VPWR VPWR _31265_/S sky130_fd_sc_hd__buf_4
Xoutput124 _31990_/Q VGND VGND VPWR VPWR D1[40] sky130_fd_sc_hd__buf_2
XFILLER_138_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput135 _32000_/Q VGND VGND VPWR VPWR D1[50] sky130_fd_sc_hd__buf_2
Xoutput146 _32010_/Q VGND VGND VPWR VPWR D1[60] sky130_fd_sc_hd__buf_2
Xoutput157 _36186_/Q VGND VGND VPWR VPWR D2[12] sky130_fd_sc_hd__buf_2
XFILLER_86_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput168 _36196_/Q VGND VGND VPWR VPWR D2[22] sky130_fd_sc_hd__buf_2
XFILLER_138_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput179 _36206_/Q VGND VGND VPWR VPWR D2[32] sky130_fd_sc_hd__buf_2
X_31177_ _35807_/Q input9/X _31181_/S VGND VGND VPWR VPWR _31178_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30128_ _35310_/Q _29151_/X _30142_/S VGND VGND VPWR VPWR _30129_/A sky130_fd_sc_hd__mux2_1
X_19939_ _19652_/X _19937_/X _19938_/X _19655_/X VGND VGND VPWR VPWR _19939_/X sky130_fd_sc_hd__a22o_1
X_35985_ _35985_/CLK _35985_/D VGND VGND VPWR VPWR _35985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_110_CLK clkbuf_6_20__f_CLK/X VGND VGND VPWR VPWR _35215_/CLK sky130_fd_sc_hd__clkbuf_16
X_30059_ _30059_/A _31140_/B VGND VGND VPWR VPWR _30192_/S sky130_fd_sc_hd__nor2_8
X_34936_ _35257_/CLK _34936_/D VGND VGND VPWR VPWR _34936_/Q sky130_fd_sc_hd__dfxtp_1
X_22950_ _22950_/A VGND VGND VPWR VPWR _32036_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21901_ _21795_/X _21899_/X _21900_/X _21800_/X VGND VGND VPWR VPWR _21901_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_5_8_0_CLK clkbuf_5_9_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_8_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22881_ _22875_/X _32014_/Q _22908_/S VGND VGND VPWR VPWR _22882_/A sky130_fd_sc_hd__mux2_1
X_34867_ _34997_/CLK _34867_/D VGND VGND VPWR VPWR _34867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24620_ _24620_/A VGND VGND VPWR VPWR _32799_/D sky130_fd_sc_hd__clkbuf_1
X_21832_ _21832_/A VGND VGND VPWR VPWR _36206_/D sky130_fd_sc_hd__buf_6
X_33818_ _35738_/CLK _33818_/D VGND VGND VPWR VPWR _33818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34798_ _35313_/CLK _34798_/D VGND VGND VPWR VPWR _34798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24551_ _23034_/X _32768_/Q _24569_/S VGND VGND VPWR VPWR _24552_/A sky130_fd_sc_hd__mux2_1
X_21763_ _21763_/A _21763_/B _21763_/C _21763_/D VGND VGND VPWR VPWR _21764_/A sky130_fd_sc_hd__or4_1
XFILLER_93_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33749_ _34260_/CLK _33749_/D VGND VGND VPWR VPWR _33749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20714_ _33231_/Q _36111_/Q _33103_/Q _33039_/Q _20620_/X _20621_/X VGND VGND VPWR
+ VPWR _20714_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23502_ _23502_/A VGND VGND VPWR VPWR _32305_/D sky130_fd_sc_hd__clkbuf_1
X_27270_ _27270_/A VGND VGND VPWR VPWR _33987_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24482_ _24482_/A VGND VGND VPWR VPWR _32735_/D sky130_fd_sc_hd__clkbuf_1
X_21694_ _34027_/Q _33963_/Q _33899_/Q _32235_/Q _21620_/X _21621_/X VGND VGND VPWR
+ VPWR _21694_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26221_ _25103_/X _33522_/Q _26227_/S VGND VGND VPWR VPWR _26222_/A sky130_fd_sc_hd__mux2_1
X_20645_ _22395_/A VGND VGND VPWR VPWR _20645_/X sky130_fd_sc_hd__buf_8
X_23433_ _23433_/A VGND VGND VPWR VPWR _32272_/D sky130_fd_sc_hd__clkbuf_1
X_35419_ _35869_/CLK _35419_/D VGND VGND VPWR VPWR _35419_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_177_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _33548_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26152_ _25001_/X _33489_/Q _26164_/S VGND VGND VPWR VPWR _26153_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23364_ _23364_/A VGND VGND VPWR VPWR _32241_/D sky130_fd_sc_hd__clkbuf_1
X_20576_ _22361_/A VGND VGND VPWR VPWR _22455_/A sky130_fd_sc_hd__buf_12
XFILLER_137_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25103_ input30/X VGND VGND VPWR VPWR _25103_/X sky130_fd_sc_hd__clkbuf_4
X_22315_ _22102_/X _22311_/X _22314_/X _22105_/X VGND VGND VPWR VPWR _22315_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23295_ _32216_/Q _23294_/X _23301_/S VGND VGND VPWR VPWR _23296_/A sky130_fd_sc_hd__mux2_1
X_26083_ _26083_/A VGND VGND VPWR VPWR _33456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29911_ _29911_/A VGND VGND VPWR VPWR _35207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22246_ _34554_/Q _32442_/Q _34426_/Q _34362_/Q _22178_/X _22179_/X VGND VGND VPWR
+ VPWR _22246_/X sky130_fd_sc_hd__mux4_1
X_25034_ _25034_/A VGND VGND VPWR VPWR _32987_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29842_ _29842_/A VGND VGND VPWR VPWR _35174_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22177_ _22102_/X _22175_/X _22176_/X _22105_/X VGND VGND VPWR VPWR _22177_/X sky130_fd_sc_hd__a22o_1
XFILLER_160_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21128_ _34267_/Q _34203_/Q _34139_/Q _34075_/Q _20983_/X _20984_/X VGND VGND VPWR
+ VPWR _21128_/X sky130_fd_sc_hd__mux4_1
XFILLER_87_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29773_ _35142_/Q _29225_/X _29779_/S VGND VGND VPWR VPWR _29774_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26985_ _26984_/X _33858_/Q _27006_/S VGND VGND VPWR VPWR _26986_/A sky130_fd_sc_hd__mux2_1
X_28724_ _26940_/X _34676_/Q _28726_/S VGND VGND VPWR VPWR _28725_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_101_CLK clkbuf_leaf_99_CLK/A VGND VGND VPWR VPWR _35026_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21059_ _33753_/Q _33689_/Q _33625_/Q _33561_/Q _20737_/X _20738_/X VGND VGND VPWR
+ VPWR _21059_/X sky130_fd_sc_hd__mux4_1
X_25936_ _25081_/X _33387_/Q _25936_/S VGND VGND VPWR VPWR _25937_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28655_ _26838_/X _34643_/Q _28663_/S VGND VGND VPWR VPWR _28656_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25867_ _25867_/A VGND VGND VPWR VPWR _33354_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27606_ _27696_/S VGND VGND VPWR VPWR _27625_/S sky130_fd_sc_hd__buf_4
X_24818_ _24818_/A VGND VGND VPWR VPWR _32892_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28586_ _28586_/A VGND VGND VPWR VPWR _34610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25798_ _25798_/A VGND VGND VPWR VPWR _33321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27537_ _26984_/X _34114_/Q _27551_/S VGND VGND VPWR VPWR _27538_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24749_ _24749_/A VGND VGND VPWR VPWR _32859_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _35085_/Q _35021_/Q _34957_/Q _34893_/Q _16079_/X _16081_/X VGND VGND VPWR
+ VPWR _18270_/X sky130_fd_sc_hd__mux4_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27468_ _27468_/A VGND VGND VPWR VPWR _34081_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29207_ _29247_/S VGND VGND VPWR VPWR _29235_/S sky130_fd_sc_hd__buf_4
X_17221_ _17217_/X _17220_/X _17147_/X VGND VGND VPWR VPWR _17231_/C sky130_fd_sc_hd__o21ba_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26419_ _26419_/A VGND VGND VPWR VPWR _33615_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_168_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _36173_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_230_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27399_ _27399_/A VGND VGND VPWR VPWR _34048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1011 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29138_ input21/X VGND VGND VPWR VPWR _29138_/X sky130_fd_sc_hd__clkbuf_4
X_17152_ _17152_/A VGND VGND VPWR VPWR _17152_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_204_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput15 DW[22] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_8
XFILLER_196_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput26 DW[32] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_4
Xinput37 DW[42] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__buf_4
Xinput48 DW[52] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__buf_8
X_16103_ _16103_/A VGND VGND VPWR VPWR _31950_/D sky130_fd_sc_hd__clkbuf_1
Xinput59 DW[62] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__clkbuf_16
X_29069_ _29069_/A VGND VGND VPWR VPWR _34835_/D sky130_fd_sc_hd__clkbuf_1
X_17083_ _35050_/Q _34986_/Q _34922_/Q _34858_/Q _16803_/X _16804_/X VGND VGND VPWR
+ VPWR _17083_/X sky130_fd_sc_hd__mux4_1
X_31100_ _31100_/A VGND VGND VPWR VPWR _35770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16034_ _16059_/A VGND VGND VPWR VPWR _17830_/A sky130_fd_sc_hd__buf_12
XFILLER_87_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32080_ _34973_/CLK _32080_/D VGND VGND VPWR VPWR _32080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31031_ _31031_/A VGND VGND VPWR VPWR _35737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_340_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _34297_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17985_ _17769_/X _17983_/X _17984_/X _17773_/X VGND VGND VPWR VPWR _17985_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16936_ _17995_/A VGND VGND VPWR VPWR _16936_/X sky130_fd_sc_hd__clkbuf_4
X_19724_ _35764_/Q _35124_/Q _34484_/Q _33844_/Q _19440_/X _19441_/X VGND VGND VPWR
+ VPWR _19724_/X sky130_fd_sc_hd__mux4_1
X_32982_ _36052_/CLK _32982_/D VGND VGND VPWR VPWR _32982_/Q sky130_fd_sc_hd__dfxtp_1
X_35770_ _35834_/CLK _35770_/D VGND VGND VPWR VPWR _35770_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_60__f_CLK clkbuf_5_30_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_60__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34721_ _35098_/CLK _34721_/D VGND VGND VPWR VPWR _34721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31933_ _31933_/A VGND VGND VPWR VPWR _36165_/D sky130_fd_sc_hd__clkbuf_1
X_16867_ _16646_/X _16865_/X _16866_/X _16649_/X VGND VGND VPWR VPWR _16867_/X sky130_fd_sc_hd__a22o_1
X_19655_ _20165_/A VGND VGND VPWR VPWR _19655_/X sky130_fd_sc_hd__buf_4
XFILLER_37_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18606_ _18387_/X _18604_/X _18605_/X _18397_/X VGND VGND VPWR VPWR _18606_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19586_ _19299_/X _19584_/X _19585_/X _19302_/X VGND VGND VPWR VPWR _19586_/X sky130_fd_sc_hd__a22o_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34652_ _34781_/CLK _34652_/D VGND VGND VPWR VPWR _34652_/Q sky130_fd_sc_hd__dfxtp_1
X_31864_ _31864_/A VGND VGND VPWR VPWR _36132_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16798_ _35298_/Q _35234_/Q _35170_/Q _32290_/Q _16653_/X _16654_/X VGND VGND VPWR
+ VPWR _16798_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33603_ _33795_/CLK _33603_/D VGND VGND VPWR VPWR _33603_/Q sky130_fd_sc_hd__dfxtp_1
X_18537_ _18533_/X _18536_/X _18400_/X VGND VGND VPWR VPWR _18538_/D sky130_fd_sc_hd__o21ba_1
XFILLER_34_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30815_ _30815_/A VGND VGND VPWR VPWR _35635_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31795_ _36100_/Q input50/X _31805_/S VGND VGND VPWR VPWR _31796_/A sky130_fd_sc_hd__mux2_1
X_34583_ _36202_/CLK _34583_/D VGND VGND VPWR VPWR _34583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18468_ _34512_/Q _32400_/Q _34384_/Q _34320_/Q _18466_/X _18467_/X VGND VGND VPWR
+ VPWR _18468_/X sky130_fd_sc_hd__mux4_1
X_30746_ _30746_/A VGND VGND VPWR VPWR _35602_/D sky130_fd_sc_hd__clkbuf_1
X_33534_ _34303_/CLK _33534_/D VGND VGND VPWR VPWR _33534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17419_ _33012_/Q _32948_/Q _32884_/Q _32820_/Q _17342_/X _17343_/X VGND VGND VPWR
+ VPWR _17419_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_159_CLK clkbuf_6_30__f_CLK/X VGND VGND VPWR VPWR _34251_/CLK sky130_fd_sc_hd__clkbuf_16
X_33465_ _34297_/CLK _33465_/D VGND VGND VPWR VPWR _33465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18399_ input82/X input81/X VGND VGND VPWR VPWR _20167_/A sky130_fd_sc_hd__or2b_4
X_30677_ _35570_/Q _29163_/X _30683_/S VGND VGND VPWR VPWR _30678_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35204_ _35332_/CLK _35204_/D VGND VGND VPWR VPWR _35204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20430_ _20208_/X _20428_/X _20429_/X _20211_/X VGND VGND VPWR VPWR _20430_/X sky130_fd_sc_hd__a22o_1
XFILLER_165_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32416_ _35294_/CLK _32416_/D VGND VGND VPWR VPWR _32416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36184_ _36185_/CLK _36184_/D VGND VGND VPWR VPWR _36184_/Q sky130_fd_sc_hd__dfxtp_1
X_33396_ _33779_/CLK _33396_/D VGND VGND VPWR VPWR _33396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20361_ _20160_/X _20359_/X _20360_/X _20165_/X VGND VGND VPWR VPWR _20361_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35135_ _35837_/CLK _35135_/D VGND VGND VPWR VPWR _35135_/Q sky130_fd_sc_hd__dfxtp_1
X_32347_ _36121_/CLK _32347_/D VGND VGND VPWR VPWR _32347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22100_ _22453_/A VGND VGND VPWR VPWR _22100_/X sky130_fd_sc_hd__clkbuf_4
X_23080_ input88/X VGND VGND VPWR VPWR _30329_/A sky130_fd_sc_hd__buf_6
X_35066_ _35386_/CLK _35066_/D VGND VGND VPWR VPWR _35066_/Q sky130_fd_sc_hd__dfxtp_1
X_20292_ _20005_/X _20290_/X _20291_/X _20008_/X VGND VGND VPWR VPWR _20292_/X sky130_fd_sc_hd__a22o_1
X_32278_ _35286_/CLK _32278_/D VGND VGND VPWR VPWR _32278_/Q sky130_fd_sc_hd__dfxtp_1
X_22031_ _22025_/X _22030_/X _21747_/X VGND VGND VPWR VPWR _22039_/C sky130_fd_sc_hd__o21ba_1
X_34017_ _34017_/CLK _34017_/D VGND VGND VPWR VPWR _34017_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31229_ _31229_/A VGND VGND VPWR VPWR _35831_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_331_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _36023_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_1062 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26770_ _26770_/A VGND VGND VPWR VPWR _33781_/D sky130_fd_sc_hd__clkbuf_1
X_35968_ _35968_/CLK _35968_/D VGND VGND VPWR VPWR _35968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23982_ _23982_/A VGND VGND VPWR VPWR _32529_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25721_ _33286_/Q _24419_/X _25727_/S VGND VGND VPWR VPWR _25722_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34919_ _35302_/CLK _34919_/D VGND VGND VPWR VPWR _34919_/Q sky130_fd_sc_hd__dfxtp_1
X_22933_ _22932_/X _32031_/Q _22939_/S VGND VGND VPWR VPWR _22934_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35899_ _35965_/CLK _35899_/D VGND VGND VPWR VPWR _35899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28440_ _26919_/X _34541_/Q _28456_/S VGND VGND VPWR VPWR _28441_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25652_ _33253_/Q _24317_/X _25664_/S VGND VGND VPWR VPWR _25653_/A sky130_fd_sc_hd__mux2_1
X_22864_ _20597_/X _22862_/X _22863_/X _20603_/X VGND VGND VPWR VPWR _22864_/X sky130_fd_sc_hd__a22o_1
XFILLER_71_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24603_ _24603_/A VGND VGND VPWR VPWR _32791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28371_ _34509_/Q _24440_/X _28371_/S VGND VGND VPWR VPWR _28372_/A sky130_fd_sc_hd__mux2_1
X_21815_ _35822_/Q _32199_/Q _35694_/Q _35630_/Q _21560_/X _21561_/X VGND VGND VPWR
+ VPWR _21815_/X sky130_fd_sc_hd__mux4_1
X_25583_ _33222_/Q _24419_/X _25589_/S VGND VGND VPWR VPWR _25584_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_398_CLK clkbuf_6_34__f_CLK/X VGND VGND VPWR VPWR _35564_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22795_ _32523_/Q _32395_/Q _32075_/Q _36043_/Q _22582_/X _21607_/A VGND VGND VPWR
+ VPWR _22795_/X sky130_fd_sc_hd__mux4_1
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27322_ _34012_/Q _24289_/X _27332_/S VGND VGND VPWR VPWR _27323_/A sky130_fd_sc_hd__mux2_1
XPHY_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24534_ _23010_/X _32760_/Q _24548_/S VGND VGND VPWR VPWR _24535_/A sky130_fd_sc_hd__mux2_1
XPHY_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21746_ _21599_/X _21744_/X _21745_/X _21602_/X VGND VGND VPWR VPWR _21746_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27253_ _27253_/A VGND VGND VPWR VPWR _33979_/D sky130_fd_sc_hd__clkbuf_1
X_24465_ _24465_/A VGND VGND VPWR VPWR _32727_/D sky130_fd_sc_hd__clkbuf_1
X_21677_ _21599_/X _21673_/X _21676_/X _21602_/X VGND VGND VPWR VPWR _21677_/X sky130_fd_sc_hd__a22o_1
XFILLER_184_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26204_ _25078_/X _33514_/Q _26206_/S VGND VGND VPWR VPWR _26205_/A sky130_fd_sc_hd__mux2_1
X_23416_ _23416_/A VGND VGND VPWR VPWR _32266_/D sky130_fd_sc_hd__clkbuf_1
X_20628_ _22582_/A VGND VGND VPWR VPWR _20628_/X sky130_fd_sc_hd__buf_6
X_27184_ _27184_/A VGND VGND VPWR VPWR _33946_/D sky130_fd_sc_hd__clkbuf_1
X_24396_ _24396_/A VGND VGND VPWR VPWR _32702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26135_ _26135_/A VGND VGND VPWR VPWR _33481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23347_ _23347_/A VGND VGND VPWR VPWR _32233_/D sky130_fd_sc_hd__clkbuf_1
X_20559_ _35853_/Q _32233_/Q _35725_/Q _35661_/Q _18289_/X _18291_/X VGND VGND VPWR
+ VPWR _20559_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26066_ _26066_/A VGND VGND VPWR VPWR _33448_/D sky130_fd_sc_hd__clkbuf_1
X_23278_ _32210_/Q _23277_/X _23301_/S VGND VGND VPWR VPWR _23279_/A sky130_fd_sc_hd__mux2_1
X_25017_ _25016_/X _32982_/Q _25020_/S VGND VGND VPWR VPWR _25018_/A sky130_fd_sc_hd__mux2_1
X_22229_ _22582_/A VGND VGND VPWR VPWR _22229_/X sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_322_CLK clkbuf_6_38__f_CLK/X VGND VGND VPWR VPWR _35574_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29825_ _29825_/A VGND VGND VPWR VPWR _35166_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17770_ _17770_/A VGND VGND VPWR VPWR _17770_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_43_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29756_ _35134_/Q _29200_/X _29758_/S VGND VGND VPWR VPWR _29757_/A sky130_fd_sc_hd__mux2_1
X_26968_ input42/X VGND VGND VPWR VPWR _26968_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_134_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16721_ _17931_/A VGND VGND VPWR VPWR _16721_/X sky130_fd_sc_hd__buf_6
X_25919_ _25919_/A VGND VGND VPWR VPWR _33378_/D sky130_fd_sc_hd__clkbuf_1
X_28707_ _28776_/S VGND VGND VPWR VPWR _28726_/S sky130_fd_sc_hd__buf_4
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29687_ _35101_/Q _29098_/X _29695_/S VGND VGND VPWR VPWR _29688_/A sky130_fd_sc_hd__mux2_1
X_26899_ _26899_/A VGND VGND VPWR VPWR _33830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19440_ _20294_/A VGND VGND VPWR VPWR _19440_/X sky130_fd_sc_hd__buf_6
X_28638_ _28638_/A VGND VGND VPWR VPWR _34635_/D sky130_fd_sc_hd__clkbuf_1
X_16652_ _34782_/Q _34718_/Q _34654_/Q _34590_/Q _16582_/X _16583_/X VGND VGND VPWR
+ VPWR _16652_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19371_ _35754_/Q _35114_/Q _34474_/Q _33834_/Q _19087_/X _19088_/X VGND VGND VPWR
+ VPWR _19371_/X sky130_fd_sc_hd__mux4_1
XFILLER_216_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16583_ _17995_/A VGND VGND VPWR VPWR _16583_/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_389_CLK clkbuf_6_35__f_CLK/X VGND VGND VPWR VPWR _35052_/CLK sky130_fd_sc_hd__clkbuf_16
X_28569_ _28569_/A VGND VGND VPWR VPWR _34602_/D sky130_fd_sc_hd__clkbuf_1
X_30600_ _31140_/A _30600_/B VGND VGND VPWR VPWR _30733_/S sky130_fd_sc_hd__nor2_8
XFILLER_188_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18322_ _33230_/Q _36110_/Q _33102_/Q _33038_/Q _18320_/X _18321_/X VGND VGND VPWR
+ VPWR _18322_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31580_ _35998_/Q input8/X _31586_/S VGND VGND VPWR VPWR _31581_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _33293_/Q _36173_/Q _33165_/Q _33101_/Q _16028_/X _17157_/A VGND VGND VPWR
+ VPWR _18253_/X sky130_fd_sc_hd__mux4_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30531_ _30531_/A VGND VGND VPWR VPWR _35500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17204_ _34030_/Q _33966_/Q _33902_/Q _32238_/Q _17020_/X _17021_/X VGND VGND VPWR
+ VPWR _17204_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33250_ _36132_/CLK _33250_/D VGND VGND VPWR VPWR _33250_/Q sky130_fd_sc_hd__dfxtp_1
X_30462_ _30462_/A VGND VGND VPWR VPWR _35468_/D sky130_fd_sc_hd__clkbuf_1
X_18184_ _18184_/A VGND VGND VPWR VPWR _32010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32201_ _35951_/CLK _32201_/D VGND VGND VPWR VPWR _32201_/Q sky130_fd_sc_hd__dfxtp_1
X_17135_ _17063_/X _17133_/X _17134_/X _17067_/X VGND VGND VPWR VPWR _17135_/X sky130_fd_sc_hd__a22o_1
X_33181_ _35933_/CLK _33181_/D VGND VGND VPWR VPWR _33181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30393_ _30393_/A VGND VGND VPWR VPWR _35435_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32132_ _35814_/CLK _32132_/D VGND VGND VPWR VPWR _32132_/Q sky130_fd_sc_hd__dfxtp_1
X_17066_ _33002_/Q _32938_/Q _32874_/Q _32810_/Q _16989_/X _16990_/X VGND VGND VPWR
+ VPWR _17066_/X sky130_fd_sc_hd__mux4_1
X_16017_ _16059_/A VGND VGND VPWR VPWR _17762_/A sky130_fd_sc_hd__buf_12
X_32063_ _36031_/CLK _32063_/D VGND VGND VPWR VPWR _32063_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_313_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _34745_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31014_ _31014_/A VGND VGND VPWR VPWR _35729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35822_ _35822_/CLK _35822_/D VGND VGND VPWR VPWR _35822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17968_ _17964_/X _17967_/X _17867_/X VGND VGND VPWR VPWR _17969_/D sky130_fd_sc_hd__o21ba_1
XFILLER_214_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19707_ _19703_/X _19706_/X _19428_/X VGND VGND VPWR VPWR _19739_/A sky130_fd_sc_hd__o21ba_1
X_35753_ _35879_/CLK _35753_/D VGND VGND VPWR VPWR _35753_/Q sky130_fd_sc_hd__dfxtp_1
X_16919_ _17978_/A VGND VGND VPWR VPWR _16919_/X sky130_fd_sc_hd__buf_8
X_32965_ _32965_/CLK _32965_/D VGND VGND VPWR VPWR _32965_/Q sky130_fd_sc_hd__dfxtp_1
X_17899_ _17899_/A _17899_/B _17899_/C _17899_/D VGND VGND VPWR VPWR _17900_/A sky130_fd_sc_hd__or4_4
XFILLER_226_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34704_ _35280_/CLK _34704_/D VGND VGND VPWR VPWR _34704_/Q sky130_fd_sc_hd__dfxtp_1
X_31916_ _31916_/A VGND VGND VPWR VPWR _36157_/D sky130_fd_sc_hd__clkbuf_1
X_19638_ _32754_/Q _32690_/Q _32626_/Q _36082_/Q _19572_/X _19356_/X VGND VGND VPWR
+ VPWR _19638_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35684_ _35811_/CLK _35684_/D VGND VGND VPWR VPWR _35684_/Q sky130_fd_sc_hd__dfxtp_1
X_32896_ _32962_/CLK _32896_/D VGND VGND VPWR VPWR _32896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34635_ _35339_/CLK _34635_/D VGND VGND VPWR VPWR _34635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19569_ _34032_/Q _33968_/Q _33904_/Q _32240_/Q _19320_/X _19321_/X VGND VGND VPWR
+ VPWR _19569_/X sky130_fd_sc_hd__mux4_1
X_31847_ _31847_/A VGND VGND VPWR VPWR _36124_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21600_ _35560_/Q _35496_/Q _35432_/Q _35368_/Q _21497_/X _21498_/X VGND VGND VPWR
+ VPWR _21600_/X sky130_fd_sc_hd__mux4_1
X_22580_ _33284_/Q _36164_/Q _33156_/Q _33092_/Q _22364_/X _22365_/X VGND VGND VPWR
+ VPWR _22580_/X sky130_fd_sc_hd__mux4_1
XFILLER_181_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34566_ _35078_/CLK _34566_/D VGND VGND VPWR VPWR _34566_/Q sky130_fd_sc_hd__dfxtp_1
X_31778_ _36092_/Q input41/X _31784_/S VGND VGND VPWR VPWR _31779_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21531_ _35558_/Q _35494_/Q _35430_/Q _35366_/Q _21497_/X _21498_/X VGND VGND VPWR
+ VPWR _21531_/X sky130_fd_sc_hd__mux4_1
X_33517_ _34293_/CLK _33517_/D VGND VGND VPWR VPWR _33517_/Q sky130_fd_sc_hd__dfxtp_1
X_30729_ _35595_/Q _29240_/X _30733_/S VGND VGND VPWR VPWR _30730_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34497_ _36038_/CLK _34497_/D VGND VGND VPWR VPWR _34497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36236_ _36237_/CLK _36236_/D VGND VGND VPWR VPWR _36236_/Q sky130_fd_sc_hd__dfxtp_1
X_24250_ _32655_/Q _24249_/X _24274_/S VGND VGND VPWR VPWR _24251_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21462_ _35812_/Q _32188_/Q _35684_/Q _35620_/Q _21207_/X _21208_/X VGND VGND VPWR
+ VPWR _21462_/X sky130_fd_sc_hd__mux4_1
XFILLER_193_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33448_ _33512_/CLK _33448_/D VGND VGND VPWR VPWR _33448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20413_ _33224_/Q _32584_/Q _35976_/Q _35912_/Q _18375_/X _18376_/X VGND VGND VPWR
+ VPWR _20413_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23201_ _23201_/A VGND VGND VPWR VPWR _32182_/D sky130_fd_sc_hd__clkbuf_1
X_36167_ _36167_/CLK _36167_/D VGND VGND VPWR VPWR _36167_/Q sky130_fd_sc_hd__dfxtp_1
X_33379_ _33635_/CLK _33379_/D VGND VGND VPWR VPWR _33379_/Q sky130_fd_sc_hd__dfxtp_1
X_21393_ _21246_/X _21391_/X _21392_/X _21249_/X VGND VGND VPWR VPWR _21393_/X sky130_fd_sc_hd__a22o_1
X_24181_ _24181_/A VGND VGND VPWR VPWR _32623_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20344_ _20061_/X _20342_/X _20343_/X _20067_/X VGND VGND VPWR VPWR _20344_/X sky130_fd_sc_hd__a22o_1
X_35118_ _35822_/CLK _35118_/D VGND VGND VPWR VPWR _35118_/Q sky130_fd_sc_hd__dfxtp_1
X_23132_ _23132_/A VGND VGND VPWR VPWR _32156_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36098_ _36098_/CLK _36098_/D VGND VGND VPWR VPWR _36098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27940_ _34304_/Q _24400_/X _27958_/S VGND VGND VPWR VPWR _27941_/A sky130_fd_sc_hd__mux2_1
X_23063_ _23062_/X _32073_/Q _23063_/S VGND VGND VPWR VPWR _23064_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20275_ _34052_/Q _33988_/Q _33924_/Q _32260_/Q _20026_/X _20027_/X VGND VGND VPWR
+ VPWR _20275_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_1340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_304_CLK clkbuf_6_50__f_CLK/X VGND VGND VPWR VPWR _35707_/CLK sky130_fd_sc_hd__clkbuf_16
X_35049_ _35943_/CLK _35049_/D VGND VGND VPWR VPWR _35049_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22014_ _22506_/A VGND VGND VPWR VPWR _22014_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27871_ _27871_/A VGND VGND VPWR VPWR _34271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26822_ _30735_/B _31410_/A VGND VGND VPWR VPWR _27018_/S sky130_fd_sc_hd__nand2_8
XTAP_5438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29610_ _29610_/A VGND VGND VPWR VPWR _35064_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29541_ _29652_/S VGND VGND VPWR VPWR _29560_/S sky130_fd_sc_hd__buf_4
XTAP_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26753_ _33773_/Q _24342_/X _26769_/S VGND VGND VPWR VPWR _26754_/A sky130_fd_sc_hd__mux2_1
X_23965_ _23965_/A VGND VGND VPWR VPWR _32522_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25704_ _33278_/Q _24394_/X _25706_/S VGND VGND VPWR VPWR _25705_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29472_ _23274_/X _34999_/Q _29488_/S VGND VGND VPWR VPWR _29473_/A sky130_fd_sc_hd__mux2_1
X_22916_ _22916_/A VGND VGND VPWR VPWR _32025_/D sky130_fd_sc_hd__clkbuf_1
X_26684_ _26684_/A VGND VGND VPWR VPWR _33741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23896_ _23896_/A VGND VGND VPWR VPWR _32489_/D sky130_fd_sc_hd__clkbuf_1
X_28423_ _26894_/X _34533_/Q _28435_/S VGND VGND VPWR VPWR _28424_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25635_ _33245_/Q _24292_/X _25643_/S VGND VGND VPWR VPWR _25636_/A sky130_fd_sc_hd__mux2_1
X_22847_ _20614_/X _22845_/X _22846_/X _20623_/X VGND VGND VPWR VPWR _22847_/X sky130_fd_sc_hd__a22o_1
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28354_ _28354_/A VGND VGND VPWR VPWR _34500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25566_ _33214_/Q _24394_/X _25568_/S VGND VGND VPWR VPWR _25567_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22778_ _20644_/X _22776_/X _22777_/X _20654_/X VGND VGND VPWR VPWR _22778_/X sky130_fd_sc_hd__a22o_1
XFILLER_231_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27305_ _34004_/Q _24264_/X _27311_/S VGND VGND VPWR VPWR _27306_/A sky130_fd_sc_hd__mux2_1
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24517_ _22985_/X _32752_/Q _24527_/S VGND VGND VPWR VPWR _24518_/A sky130_fd_sc_hd__mux2_1
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28285_ _28285_/A VGND VGND VPWR VPWR _34467_/D sky130_fd_sc_hd__clkbuf_1
X_21729_ _21722_/X _21727_/X _21728_/X VGND VGND VPWR VPWR _21763_/A sky130_fd_sc_hd__o21ba_1
XFILLER_169_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25497_ _33181_/Q _24292_/X _25505_/S VGND VGND VPWR VPWR _25498_/A sky130_fd_sc_hd__mux2_1
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_786 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27236_ _27236_/A VGND VGND VPWR VPWR _33971_/D sky130_fd_sc_hd__clkbuf_1
X_24448_ _22883_/X _32719_/Q _24464_/S VGND VGND VPWR VPWR _24449_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27167_ _27167_/A VGND VGND VPWR VPWR _33938_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24379_ input38/X VGND VGND VPWR VPWR _24379_/X sky130_fd_sc_hd__buf_4
XFILLER_181_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26118_ _25150_/X _33473_/Q _26134_/S VGND VGND VPWR VPWR _26119_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27098_ _26934_/X _33906_/Q _27104_/S VGND VGND VPWR VPWR _27099_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18940_ _18934_/X _18939_/X _18730_/X _18731_/X VGND VGND VPWR VPWR _18961_/B sky130_fd_sc_hd__o211a_2
X_26049_ _26049_/A VGND VGND VPWR VPWR _33440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18871_ _32476_/Q _32348_/Q _32028_/Q _35996_/Q _18870_/X _18658_/X VGND VGND VPWR
+ VPWR _18871_/X sky130_fd_sc_hd__mux4_1
XTAP_6640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17822_ _17507_/X _17820_/X _17821_/X _17512_/X VGND VGND VPWR VPWR _17822_/X sky130_fd_sc_hd__a22o_1
X_29808_ _29808_/A VGND VGND VPWR VPWR _35158_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29739_ _29787_/S VGND VGND VPWR VPWR _29758_/S sky130_fd_sc_hd__buf_4
X_17753_ _17753_/A VGND VGND VPWR VPWR _31997_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_207_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16704_ _32736_/Q _32672_/Q _32608_/Q _36064_/Q _16566_/X _16703_/X VGND VGND VPWR
+ VPWR _16704_/X sky130_fd_sc_hd__mux4_1
X_17684_ _33788_/Q _33724_/Q _33660_/Q _33596_/Q _17549_/X _17550_/X VGND VGND VPWR
+ VPWR _17684_/X sky130_fd_sc_hd__mux4_1
X_32750_ _36078_/CLK _32750_/D VGND VGND VPWR VPWR _32750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31701_ _31701_/A VGND VGND VPWR VPWR _36055_/D sky130_fd_sc_hd__clkbuf_1
X_19423_ _20129_/A VGND VGND VPWR VPWR _19423_/X sky130_fd_sc_hd__buf_4
X_16635_ _32478_/Q _32350_/Q _32030_/Q _35998_/Q _16570_/X _16358_/X VGND VGND VPWR
+ VPWR _16635_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32681_ _36137_/CLK _32681_/D VGND VGND VPWR VPWR _32681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34420_ _35250_/CLK _34420_/D VGND VGND VPWR VPWR _34420_/Q sky130_fd_sc_hd__dfxtp_1
X_31632_ _31632_/A VGND VGND VPWR VPWR _36022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16566_ _17978_/A VGND VGND VPWR VPWR _16566_/X sky130_fd_sc_hd__buf_6
X_19354_ _19350_/X _19353_/X _19075_/X VGND VGND VPWR VPWR _19386_/A sky130_fd_sc_hd__o21ba_1
XFILLER_210_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18305_ _20256_/A VGND VGND VPWR VPWR _18305_/X sky130_fd_sc_hd__buf_6
X_31563_ _35990_/Q input63/X _31565_/S VGND VGND VPWR VPWR _31564_/A sky130_fd_sc_hd__mux2_1
X_34351_ _35758_/CLK _34351_/D VGND VGND VPWR VPWR _34351_/Q sky130_fd_sc_hd__dfxtp_1
X_19285_ _32744_/Q _32680_/Q _32616_/Q _36072_/Q _19219_/X _19003_/X VGND VGND VPWR
+ VPWR _19285_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16497_ _33498_/Q _33434_/Q _33370_/Q _33306_/Q _16417_/X _16418_/X VGND VGND VPWR
+ VPWR _16497_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18236_ _34828_/Q _34764_/Q _34700_/Q _34636_/Q _17994_/X _17995_/X VGND VGND VPWR
+ VPWR _18236_/X sky130_fd_sc_hd__mux4_1
X_33302_ _36228_/CLK _33302_/D VGND VGND VPWR VPWR _33302_/Q sky130_fd_sc_hd__dfxtp_1
X_30514_ _30514_/A VGND VGND VPWR VPWR _35492_/D sky130_fd_sc_hd__clkbuf_1
X_34282_ _34282_/CLK _34282_/D VGND VGND VPWR VPWR _34282_/Q sky130_fd_sc_hd__dfxtp_1
X_31494_ _31494_/A VGND VGND VPWR VPWR _35957_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33233_ _36114_/CLK _33233_/D VGND VGND VPWR VPWR _33233_/Q sky130_fd_sc_hd__dfxtp_1
X_36021_ _36021_/CLK _36021_/D VGND VGND VPWR VPWR _36021_/Q sky130_fd_sc_hd__dfxtp_1
X_30445_ _23316_/X _35460_/Q _30455_/S VGND VGND VPWR VPWR _30446_/A sky130_fd_sc_hd__mux2_1
X_18167_ _17154_/A _18165_/X _18166_/X _17159_/A VGND VGND VPWR VPWR _18167_/X sky130_fd_sc_hd__a22o_1
XFILLER_15_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_90_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _35284_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17118_ _17118_/A _17118_/B _17118_/C _17118_/D VGND VGND VPWR VPWR _17119_/A sky130_fd_sc_hd__or4_4
XFILLER_209_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33164_ _36173_/CLK _33164_/D VGND VGND VPWR VPWR _33164_/Q sky130_fd_sc_hd__dfxtp_1
X_18098_ _33544_/Q _33480_/Q _33416_/Q _33352_/Q _17829_/X _17830_/X VGND VGND VPWR
+ VPWR _18098_/X sky130_fd_sc_hd__mux4_1
X_30376_ _23152_/X _35427_/Q _30392_/S VGND VGND VPWR VPWR _30377_/A sky130_fd_sc_hd__mux2_1
XFILLER_239_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32115_ _35555_/CLK _32115_/D VGND VGND VPWR VPWR _32115_/Q sky130_fd_sc_hd__dfxtp_1
X_17049_ _34282_/Q _34218_/Q _34154_/Q _34090_/Q _16736_/X _16737_/X VGND VGND VPWR
+ VPWR _17049_/X sky130_fd_sc_hd__mux4_1
XFILLER_217_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33095_ _36167_/CLK _33095_/D VGND VGND VPWR VPWR _33095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20060_ _20056_/X _20059_/X _19781_/X VGND VGND VPWR VPWR _20092_/A sky130_fd_sc_hd__o21ba_1
XFILLER_131_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32046_ _36013_/CLK _32046_/D VGND VGND VPWR VPWR _32046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1062 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_959 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35805_ _35809_/CLK _35805_/D VGND VGND VPWR VPWR _35805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33997_ _34060_/CLK _33997_/D VGND VGND VPWR VPWR _33997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35736_ _35738_/CLK _35736_/D VGND VGND VPWR VPWR _35736_/Q sky130_fd_sc_hd__dfxtp_1
X_23750_ _23750_/A VGND VGND VPWR VPWR _32420_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20962_ _20957_/X _20959_/X _20960_/X _20961_/X VGND VGND VPWR VPWR _20962_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32948_ _33013_/CLK _32948_/D VGND VGND VPWR VPWR _32948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22701_ _22697_/X _22700_/X _22434_/X VGND VGND VPWR VPWR _22723_/A sky130_fd_sc_hd__o21ba_2
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23681_ _23681_/A VGND VGND VPWR VPWR _32389_/D sky130_fd_sc_hd__clkbuf_1
X_35667_ _35667_/CLK _35667_/D VGND VGND VPWR VPWR _35667_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20893_ _22460_/A VGND VGND VPWR VPWR _20893_/X sky130_fd_sc_hd__buf_4
X_32879_ _33007_/CLK _32879_/D VGND VGND VPWR VPWR _32879_/Q sky130_fd_sc_hd__dfxtp_1
X_25420_ _25420_/A VGND VGND VPWR VPWR _33146_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22632_ _22628_/X _22631_/X _22467_/X VGND VGND VPWR VPWR _22633_/D sky130_fd_sc_hd__o21ba_1
X_34618_ _35771_/CLK _34618_/D VGND VGND VPWR VPWR _34618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35598_ _35727_/CLK _35598_/D VGND VGND VPWR VPWR _35598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1041 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25351_ _25351_/A VGND VGND VPWR VPWR _33113_/D sky130_fd_sc_hd__clkbuf_1
X_22563_ _35331_/Q _35267_/Q _35203_/Q _32323_/Q _22312_/X _22313_/X VGND VGND VPWR
+ VPWR _22563_/X sky130_fd_sc_hd__mux4_1
X_34549_ _34805_/CLK _34549_/D VGND VGND VPWR VPWR _34549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24302_ _32672_/Q _24301_/X _24305_/S VGND VGND VPWR VPWR _24303_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28070_ _26971_/X _34366_/Q _28072_/S VGND VGND VPWR VPWR _28071_/A sky130_fd_sc_hd__mux2_1
X_21514_ _21442_/X _21512_/X _21513_/X _21447_/X VGND VGND VPWR VPWR _21514_/X sky130_fd_sc_hd__a22o_1
X_25282_ _25282_/A VGND VGND VPWR VPWR _33081_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22494_ _22455_/X _22492_/X _22493_/X _22458_/X VGND VGND VPWR VPWR _22494_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27021_ _27426_/A _31410_/B VGND VGND VPWR VPWR _27154_/S sky130_fd_sc_hd__nand2_8
X_36219_ _36220_/CLK _36219_/D VGND VGND VPWR VPWR _36219_/Q sky130_fd_sc_hd__dfxtp_1
X_24233_ _24233_/A VGND VGND VPWR VPWR _32648_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21445_ _33764_/Q _33700_/Q _33636_/Q _33572_/Q _21443_/X _21444_/X VGND VGND VPWR
+ VPWR _21445_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_81_CLK clkbuf_leaf_87_CLK/A VGND VGND VPWR VPWR _35667_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24164_ _24164_/A VGND VGND VPWR VPWR _32615_/D sky130_fd_sc_hd__clkbuf_1
X_21376_ _21369_/X _21374_/X _21375_/X VGND VGND VPWR VPWR _21410_/A sky130_fd_sc_hd__o21ba_1
XFILLER_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20327_ _35333_/Q _35269_/Q _35205_/Q _32325_/Q _20012_/X _20013_/X VGND VGND VPWR
+ VPWR _20327_/X sky130_fd_sc_hd__mux4_1
X_23115_ _32151_/Q _23114_/X _23115_/S VGND VGND VPWR VPWR _23116_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24095_ _24095_/A VGND VGND VPWR VPWR _32583_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28972_ _28972_/A VGND VGND VPWR VPWR _34793_/D sky130_fd_sc_hd__clkbuf_1
X_20258_ _35587_/Q _35523_/Q _35459_/Q _35395_/Q _20256_/X _20257_/X VGND VGND VPWR
+ VPWR _20258_/X sky130_fd_sc_hd__mux4_1
X_23046_ _23046_/A VGND VGND VPWR VPWR _32067_/D sky130_fd_sc_hd__clkbuf_1
X_27923_ _34296_/Q _24376_/X _27937_/S VGND VGND VPWR VPWR _27924_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27854_ _27854_/A VGND VGND VPWR VPWR _34263_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20189_ _33217_/Q _32577_/Q _35969_/Q _35905_/Q _20080_/X _20081_/X VGND VGND VPWR
+ VPWR _20189_/X sky130_fd_sc_hd__mux4_1
XTAP_5235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26805_ _33798_/Q _24419_/X _26811_/S VGND VGND VPWR VPWR _26806_/A sky130_fd_sc_hd__mux2_1
XTAP_5268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27785_ _27785_/A VGND VGND VPWR VPWR _34230_/D sky130_fd_sc_hd__clkbuf_1
X_24997_ _24997_/A VGND VGND VPWR VPWR _32975_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29524_ _29524_/A VGND VGND VPWR VPWR _35023_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26736_ _33765_/Q _24317_/X _26748_/S VGND VGND VPWR VPWR _26737_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23948_ _23041_/X _32514_/Q _23962_/S VGND VGND VPWR VPWR _23949_/A sky130_fd_sc_hd__mux2_1
XTAP_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_800 _23075_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_811 _22910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29455_ _23247_/X _34991_/Q _29467_/S VGND VGND VPWR VPWR _29456_/A sky130_fd_sc_hd__mux2_1
XANTENNA_822 _23421_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26667_ _25162_/X _33733_/Q _26675_/S VGND VGND VPWR VPWR _26668_/A sky130_fd_sc_hd__mux2_1
XTAP_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_833 _23136_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23879_ _23879_/A VGND VGND VPWR VPWR _32481_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_844 _23333_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16420_ _34008_/Q _33944_/Q _33880_/Q _32152_/Q _16314_/X _16315_/X VGND VGND VPWR
+ VPWR _16420_/X sky130_fd_sc_hd__mux4_1
XANTENNA_855 _24342_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_866 _24428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25618_ _33237_/Q _24267_/X _25622_/S VGND VGND VPWR VPWR _25619_/A sky130_fd_sc_hd__mux2_1
X_28406_ _26869_/X _34525_/Q _28414_/S VGND VGND VPWR VPWR _28407_/A sky130_fd_sc_hd__mux2_1
X_29386_ _23077_/X _34958_/Q _29404_/S VGND VGND VPWR VPWR _29387_/A sky130_fd_sc_hd__mux2_1
XANTENNA_877 _25187_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26598_ _25060_/X _33700_/Q _26612_/S VGND VGND VPWR VPWR _26599_/A sky130_fd_sc_hd__mux2_1
XANTENNA_888 _25322_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_899 _26007_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28337_ _28337_/A VGND VGND VPWR VPWR _34492_/D sky130_fd_sc_hd__clkbuf_1
X_16351_ _32726_/Q _32662_/Q _32598_/Q _36054_/Q _16213_/X _16350_/X VGND VGND VPWR
+ VPWR _16351_/X sky130_fd_sc_hd__mux4_1
X_25549_ _25597_/S VGND VGND VPWR VPWR _25568_/S sky130_fd_sc_hd__buf_4
XFILLER_158_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19070_ _20129_/A VGND VGND VPWR VPWR _19070_/X sky130_fd_sc_hd__buf_4
X_16282_ _32468_/Q _32340_/Q _32020_/Q _35988_/Q _16217_/X _17863_/A VGND VGND VPWR
+ VPWR _16282_/X sky130_fd_sc_hd__mux4_1
X_28268_ _28268_/A VGND VGND VPWR VPWR _34459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18021_ _17700_/X _18019_/X _18020_/X _17703_/X VGND VGND VPWR VPWR _18021_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27219_ _27219_/A VGND VGND VPWR VPWR _33963_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28199_ _26962_/X _34427_/Q _28207_/S VGND VGND VPWR VPWR _28200_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_CLK clkbuf_leaf_73_CLK/A VGND VGND VPWR VPWR _36115_/CLK sky130_fd_sc_hd__clkbuf_16
X_30230_ _30230_/A VGND VGND VPWR VPWR _35358_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_1_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_9_0_CLK/A sky130_fd_sc_hd__clkbuf_8
XFILLER_99_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30161_ _35326_/Q _29200_/X _30163_/S VGND VGND VPWR VPWR _30162_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19972_ _33211_/Q _32571_/Q _35963_/Q _35899_/Q _19727_/X _19728_/X VGND VGND VPWR
+ VPWR _19972_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18923_ _18923_/A _18923_/B _18923_/C _18923_/D VGND VGND VPWR VPWR _18924_/A sky130_fd_sc_hd__or4_2
X_30092_ _35293_/Q _29098_/X _30100_/S VGND VGND VPWR VPWR _30093_/A sky130_fd_sc_hd__mux2_1
XANTENNA_1210 _23319_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1221 _24283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1232 _24425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1243 _26007_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33920_ _33922_/CLK _33920_/D VGND VGND VPWR VPWR _33920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18854_ _35035_/Q _34971_/Q _34907_/Q _34843_/Q _18750_/X _18751_/X VGND VGND VPWR
+ VPWR _18854_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1254 _26922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1265 _29234_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1276 _17903_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17805_ _17761_/X _17803_/X _17804_/X _17767_/X VGND VGND VPWR VPWR _17805_/X sky130_fd_sc_hd__a22o_1
XANTENNA_1287 _17858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33851_ _35707_/CLK _33851_/D VGND VGND VPWR VPWR _33851_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1298 _17157_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15997_ _17860_/A VGND VGND VPWR VPWR _15997_/X sky130_fd_sc_hd__buf_4
X_18785_ _18748_/X _18783_/X _18784_/X _18753_/X VGND VGND VPWR VPWR _18785_/X sky130_fd_sc_hd__a22o_1
XTAP_5780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32802_ _32994_/CLK _32802_/D VGND VGND VPWR VPWR _32802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17736_ _17416_/X _17734_/X _17735_/X _17420_/X VGND VGND VPWR VPWR _17736_/X sky130_fd_sc_hd__a22o_1
X_30994_ _30994_/A VGND VGND VPWR VPWR _35720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33782_ _34039_/CLK _33782_/D VGND VGND VPWR VPWR _33782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35521_ _35585_/CLK _35521_/D VGND VGND VPWR VPWR _35521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32733_ _36127_/CLK _32733_/D VGND VGND VPWR VPWR _32733_/Q sky130_fd_sc_hd__dfxtp_1
X_17667_ _17796_/A VGND VGND VPWR VPWR _17667_/X sky130_fd_sc_hd__buf_4
XFILLER_51_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19406_ _19294_/X _19404_/X _19405_/X _19297_/X VGND VGND VPWR VPWR _19406_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35452_ _35517_/CLK _35452_/D VGND VGND VPWR VPWR _35452_/Q sky130_fd_sc_hd__dfxtp_1
X_16618_ _16443_/X _16616_/X _16617_/X _16446_/X VGND VGND VPWR VPWR _16618_/X sky130_fd_sc_hd__a22o_1
X_17598_ _17416_/X _17596_/X _17597_/X _17420_/X VGND VGND VPWR VPWR _17598_/X sky130_fd_sc_hd__a22o_1
X_32664_ _34265_/CLK _32664_/D VGND VGND VPWR VPWR _32664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34403_ _35932_/CLK _34403_/D VGND VGND VPWR VPWR _34403_/Q sky130_fd_sc_hd__dfxtp_1
X_19337_ _19299_/X _19335_/X _19336_/X _19302_/X VGND VGND VPWR VPWR _19337_/X sky130_fd_sc_hd__a22o_1
X_31615_ _31615_/A VGND VGND VPWR VPWR _36014_/D sky130_fd_sc_hd__clkbuf_1
X_16549_ _16543_/X _16548_/X _16441_/X VGND VGND VPWR VPWR _16557_/C sky130_fd_sc_hd__o21ba_1
XFILLER_149_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35383_ _35638_/CLK _35383_/D VGND VGND VPWR VPWR _35383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32595_ _36050_/CLK _32595_/D VGND VGND VPWR VPWR _32595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34334_ _35036_/CLK _34334_/D VGND VGND VPWR VPWR _34334_/Q sky130_fd_sc_hd__dfxtp_1
X_31546_ _31678_/S VGND VGND VPWR VPWR _31565_/S sky130_fd_sc_hd__buf_4
X_19268_ _19264_/X _19267_/X _19094_/X VGND VGND VPWR VPWR _19276_/C sky130_fd_sc_hd__o21ba_1
XFILLER_206_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18219_ _34060_/Q _33996_/Q _33932_/Q _32268_/Q _16058_/X _16060_/X VGND VGND VPWR
+ VPWR _18219_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34265_ _34265_/CLK _34265_/D VGND VGND VPWR VPWR _34265_/Q sky130_fd_sc_hd__dfxtp_1
X_19199_ _35557_/Q _35493_/Q _35429_/Q _35365_/Q _19197_/X _19198_/X VGND VGND VPWR
+ VPWR _19199_/X sky130_fd_sc_hd__mux4_1
X_31477_ _23241_/X _35949_/Q _31493_/S VGND VGND VPWR VPWR _31478_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_63_CLK clkbuf_leaf_66_CLK/A VGND VGND VPWR VPWR _35991_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36004_ _36004_/CLK _36004_/D VGND VGND VPWR VPWR _36004_/Q sky130_fd_sc_hd__dfxtp_1
X_21230_ _21096_/X _21228_/X _21229_/X _21099_/X VGND VGND VPWR VPWR _21230_/X sky130_fd_sc_hd__a22o_1
XFILLER_191_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33216_ _35906_/CLK _33216_/D VGND VGND VPWR VPWR _33216_/Q sky130_fd_sc_hd__dfxtp_1
X_30428_ _23289_/X _35452_/Q _30434_/S VGND VGND VPWR VPWR _30429_/A sky130_fd_sc_hd__mux2_1
X_34196_ _34260_/CLK _34196_/D VGND VGND VPWR VPWR _34196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21161_ _21089_/X _21159_/X _21160_/X _21094_/X VGND VGND VPWR VPWR _21161_/X sky130_fd_sc_hd__a22o_1
X_33147_ _36156_/CLK _33147_/D VGND VGND VPWR VPWR _33147_/Q sky130_fd_sc_hd__dfxtp_1
X_30359_ _23127_/X _35419_/Q _30371_/S VGND VGND VPWR VPWR _30360_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20112_ _20000_/X _20110_/X _20111_/X _20003_/X VGND VGND VPWR VPWR _20112_/X sky130_fd_sc_hd__a22o_1
XFILLER_236_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33078_ _36150_/CLK _33078_/D VGND VGND VPWR VPWR _33078_/Q sky130_fd_sc_hd__dfxtp_1
X_21092_ _33754_/Q _33690_/Q _33626_/Q _33562_/Q _21090_/X _21091_/X VGND VGND VPWR
+ VPWR _21092_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20043_ _20005_/X _20041_/X _20042_/X _20008_/X VGND VGND VPWR VPWR _20043_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24920_ _24920_/A VGND VGND VPWR VPWR _32940_/D sky130_fd_sc_hd__clkbuf_1
X_32029_ _36129_/CLK _32029_/D VGND VGND VPWR VPWR _32029_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24851_ _24851_/A VGND VGND VPWR VPWR _32908_/D sky130_fd_sc_hd__clkbuf_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23802_ _23802_/A VGND VGND VPWR VPWR _32445_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27570_ _27570_/A VGND VGND VPWR VPWR _34128_/D sky130_fd_sc_hd__clkbuf_1
X_24782_ _24782_/A VGND VGND VPWR VPWR _32875_/D sky130_fd_sc_hd__clkbuf_1
X_21994_ _21749_/X _21992_/X _21993_/X _21752_/X VGND VGND VPWR VPWR _21994_/X sky130_fd_sc_hd__a22o_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_107 _32129_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26521_ _25146_/X _33664_/Q _26539_/S VGND VGND VPWR VPWR _26522_/A sky130_fd_sc_hd__mux2_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35719_ _35848_/CLK _35719_/D VGND VGND VPWR VPWR _35719_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_118 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23733_ _23733_/A VGND VGND VPWR VPWR _32412_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20945_ _33494_/Q _33430_/Q _33366_/Q _33302_/Q _20598_/X _20599_/X VGND VGND VPWR
+ VPWR _20945_/X sky130_fd_sc_hd__mux4_1
XANTENNA_129 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_984 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29240_ input58/X VGND VGND VPWR VPWR _29240_/X sky130_fd_sc_hd__buf_2
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1019 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26452_ _26452_/A VGND VGND VPWR VPWR _33631_/D sky130_fd_sc_hd__clkbuf_1
X_23664_ _23664_/A VGND VGND VPWR VPWR _32381_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20876_ _34004_/Q _33940_/Q _33876_/Q _32148_/Q _20708_/X _20709_/X VGND VGND VPWR
+ VPWR _20876_/X sky130_fd_sc_hd__mux4_1
XFILLER_161_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25403_ _25403_/A VGND VGND VPWR VPWR _33138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22615_ _32517_/Q _32389_/Q _32069_/Q _36037_/Q _22582_/X _22370_/X VGND VGND VPWR
+ VPWR _22615_/X sky130_fd_sc_hd__mux4_1
X_29171_ _29171_/A VGND VGND VPWR VPWR _34868_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26383_ _25143_/X _33599_/Q _26383_/S VGND VGND VPWR VPWR _26384_/A sky130_fd_sc_hd__mux2_1
X_23595_ _23595_/A VGND VGND VPWR VPWR _32348_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28122_ _28122_/A VGND VGND VPWR VPWR _34390_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_37__f_CLK clkbuf_5_18_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_37__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25334_ _25334_/A VGND VGND VPWR VPWR _33105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22546_ _32771_/Q _32707_/Q _32643_/Q _36099_/Q _22225_/X _22362_/X VGND VGND VPWR
+ VPWR _22546_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28053_ _28101_/S VGND VGND VPWR VPWR _28072_/S sky130_fd_sc_hd__buf_4
X_25265_ _25265_/A VGND VGND VPWR VPWR _33073_/D sky130_fd_sc_hd__clkbuf_1
X_22477_ _22473_/X _22476_/X _22434_/X VGND VGND VPWR VPWR _22499_/A sky130_fd_sc_hd__o21ba_1
XFILLER_120_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_54_CLK clkbuf_leaf_57_CLK/A VGND VGND VPWR VPWR _35995_/CLK sky130_fd_sc_hd__clkbuf_16
X_27004_ _27004_/A VGND VGND VPWR VPWR _33864_/D sky130_fd_sc_hd__clkbuf_1
X_24216_ _23034_/X _32640_/Q _24234_/S VGND VGND VPWR VPWR _24217_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21428_ _21241_/X _21426_/X _21427_/X _21244_/X VGND VGND VPWR VPWR _21428_/X sky130_fd_sc_hd__a22o_1
X_25196_ _25196_/A VGND VGND VPWR VPWR _33040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24147_ _24147_/A VGND VGND VPWR VPWR _32607_/D sky130_fd_sc_hd__clkbuf_1
X_21359_ _35297_/Q _35233_/Q _35169_/Q _32289_/Q _21253_/X _21254_/X VGND VGND VPWR
+ VPWR _21359_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24078_ _24078_/A VGND VGND VPWR VPWR _32575_/D sky130_fd_sc_hd__clkbuf_1
X_28955_ _28955_/A VGND VGND VPWR VPWR _34785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23029_ _23028_/X _32062_/Q _23032_/S VGND VGND VPWR VPWR _23030_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27906_ _34288_/Q _24351_/X _27916_/S VGND VGND VPWR VPWR _27907_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28886_ _28886_/A VGND VGND VPWR VPWR _34752_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27837_ _34255_/Q _24249_/X _27853_/S VGND VGND VPWR VPWR _27838_/A sky130_fd_sc_hd__mux2_1
XFILLER_188_1003 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18570_ _18570_/A _18570_/B _18570_/C _18570_/D VGND VGND VPWR VPWR _18571_/A sky130_fd_sc_hd__or4_4
XTAP_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27768_ _27768_/A VGND VGND VPWR VPWR _34222_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29507_ _23330_/X _35016_/Q _29509_/S VGND VGND VPWR VPWR _29508_/A sky130_fd_sc_hd__mux2_1
XTAP_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17521_ _33527_/Q _33463_/Q _33399_/Q _33335_/Q _17476_/X _17477_/X VGND VGND VPWR
+ VPWR _17521_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26719_ _33757_/Q _24292_/X _26727_/S VGND VGND VPWR VPWR _26720_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27699_ _27831_/S VGND VGND VPWR VPWR _27718_/S sky130_fd_sc_hd__buf_6
XFILLER_45_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_630 _18857_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_641 _19355_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_652 _20211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _17408_/X _17450_/X _17451_/X _17414_/X VGND VGND VPWR VPWR _17452_/X sky130_fd_sc_hd__a22o_1
X_29438_ _23220_/X _34983_/Q _29446_/S VGND VGND VPWR VPWR _29439_/A sky130_fd_sc_hd__mux2_1
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_663 _20580_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_674 _20597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16403_ _16293_/X _16401_/X _16402_/X _16296_/X VGND VGND VPWR VPWR _16403_/X sky130_fd_sc_hd__a22o_1
XANTENNA_685 _22501_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_696 _22595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17383_ _17063_/X _17381_/X _17382_/X _17067_/X VGND VGND VPWR VPWR _17383_/X sky130_fd_sc_hd__a22o_1
X_29369_ _29369_/A VGND VGND VPWR VPWR _34950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31400_ _35913_/Q input55/X _31400_/S VGND VGND VPWR VPWR _31401_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16334_ _35285_/Q _35221_/Q _35157_/Q _32277_/Q _16300_/X _16301_/X VGND VGND VPWR
+ VPWR _16334_/X sky130_fd_sc_hd__mux4_1
X_19122_ _32483_/Q _32355_/Q _32035_/Q _36003_/Q _18870_/X _19011_/X VGND VGND VPWR
+ VPWR _19122_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32380_ _36028_/CLK _32380_/D VGND VGND VPWR VPWR _32380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31331_ _35880_/Q input19/X _31337_/S VGND VGND VPWR VPWR _31332_/A sky130_fd_sc_hd__mux2_1
X_19053_ _18941_/X _19051_/X _19052_/X _18944_/X VGND VGND VPWR VPWR _19053_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16265_ _16074_/X _16263_/X _16264_/X _16084_/X VGND VGND VPWR VPWR _16265_/X sky130_fd_sc_hd__a22o_1
XFILLER_12_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_45_CLK clkbuf_6_6__f_CLK/X VGND VGND VPWR VPWR _36062_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18004_ _18004_/A VGND VGND VPWR VPWR _32004_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_127_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31262_ _31262_/A VGND VGND VPWR VPWR _35847_/D sky130_fd_sc_hd__clkbuf_1
X_34050_ _34050_/CLK _34050_/D VGND VGND VPWR VPWR _34050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16196_ _16190_/X _16195_/X _16071_/X VGND VGND VPWR VPWR _16204_/C sky130_fd_sc_hd__o21ba_1
XFILLER_177_1430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30213_ _30213_/A VGND VGND VPWR VPWR _35350_/D sky130_fd_sc_hd__clkbuf_1
X_33001_ _36137_/CLK _33001_/D VGND VGND VPWR VPWR _33001_/Q sky130_fd_sc_hd__dfxtp_1
X_31193_ _31193_/A VGND VGND VPWR VPWR _35814_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30144_ _30192_/S VGND VGND VPWR VPWR _30163_/S sky130_fd_sc_hd__clkbuf_8
X_19955_ _33531_/Q _33467_/Q _33403_/Q _33339_/Q _19776_/X _19777_/X VGND VGND VPWR
+ VPWR _19955_/X sky130_fd_sc_hd__mux4_1
XFILLER_218_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18906_ _18902_/X _18905_/X _18730_/X _18731_/X VGND VGND VPWR VPWR _18923_/B sky130_fd_sc_hd__o211a_1
X_34952_ _35847_/CLK _34952_/D VGND VGND VPWR VPWR _34952_/Q sky130_fd_sc_hd__dfxtp_1
X_30075_ _35285_/Q _29073_/X _30079_/S VGND VGND VPWR VPWR _30076_/A sky130_fd_sc_hd__mux2_1
X_19886_ _33785_/Q _33721_/Q _33657_/Q _33593_/Q _19849_/X _19850_/X VGND VGND VPWR
+ VPWR _19886_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1040 _17152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1051 _16103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1062 _16765_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33903_ _34032_/CLK _33903_/D VGND VGND VPWR VPWR _33903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18837_ _32475_/Q _32347_/Q _32027_/Q _35995_/Q _18517_/X _18658_/X VGND VGND VPWR
+ VPWR _18837_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1073 _17164_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_34883_ _34947_/CLK _34883_/D VGND VGND VPWR VPWR _34883_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1084 _17232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1095 _17264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33834_ _35944_/CLK _33834_/D VGND VGND VPWR VPWR _33834_/Q sky130_fd_sc_hd__dfxtp_1
X_18768_ _18649_/X _18766_/X _18767_/X _18655_/X VGND VGND VPWR VPWR _18768_/X sky130_fd_sc_hd__a22o_1
XFILLER_208_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17719_ _17715_/X _17718_/X _17514_/X VGND VGND VPWR VPWR _17720_/D sky130_fd_sc_hd__o21ba_1
X_33765_ _34277_/CLK _33765_/D VGND VGND VPWR VPWR _33765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30977_ _35712_/Q _29206_/X _30995_/S VGND VGND VPWR VPWR _30978_/A sky130_fd_sc_hd__mux2_1
X_18699_ _35735_/Q _35095_/Q _34455_/Q _33815_/Q _18349_/X _18351_/X VGND VGND VPWR
+ VPWR _18699_/X sky130_fd_sc_hd__mux4_1
X_35504_ _36077_/CLK _35504_/D VGND VGND VPWR VPWR _35504_/Q sky130_fd_sc_hd__dfxtp_1
X_20730_ _34511_/Q _32399_/Q _34383_/Q _34319_/Q _20688_/X _20690_/X VGND VGND VPWR
+ VPWR _20730_/X sky130_fd_sc_hd__mux4_1
X_32716_ _36109_/CLK _32716_/D VGND VGND VPWR VPWR _32716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33696_ _34010_/CLK _33696_/D VGND VGND VPWR VPWR _33696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35435_ _35819_/CLK _35435_/D VGND VGND VPWR VPWR _35435_/Q sky130_fd_sc_hd__dfxtp_1
X_32647_ _36103_/CLK _32647_/D VGND VGND VPWR VPWR _32647_/Q sky130_fd_sc_hd__dfxtp_1
X_20661_ _35534_/Q _35470_/Q _35406_/Q _35342_/Q _20658_/X _20660_/X VGND VGND VPWR
+ VPWR _20661_/X sky130_fd_sc_hd__mux4_1
X_22400_ _34047_/Q _33983_/Q _33919_/Q _32255_/Q _22326_/X _22327_/X VGND VGND VPWR
+ VPWR _22400_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20592_ _34254_/Q _34190_/Q _34126_/Q _34062_/Q _20589_/X _20591_/X VGND VGND VPWR
+ VPWR _20592_/X sky130_fd_sc_hd__mux4_1
XFILLER_188_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23380_ _32249_/Q _23280_/X _23392_/S VGND VGND VPWR VPWR _23381_/A sky130_fd_sc_hd__mux2_1
X_35366_ _35750_/CLK _35366_/D VGND VGND VPWR VPWR _35366_/Q sky130_fd_sc_hd__dfxtp_1
X_32578_ _35903_/CLK _32578_/D VGND VGND VPWR VPWR _32578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34317_ _34317_/CLK _34317_/D VGND VGND VPWR VPWR _34317_/Q sky130_fd_sc_hd__dfxtp_1
X_22331_ _32765_/Q _32701_/Q _32637_/Q _36093_/Q _22225_/X _22009_/X VGND VGND VPWR
+ VPWR _22331_/X sky130_fd_sc_hd__mux4_1
X_31529_ _23322_/X _35974_/Q _31535_/S VGND VGND VPWR VPWR _31530_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_CLK clkbuf_6_7__f_CLK/X VGND VGND VPWR VPWR _34265_/CLK sky130_fd_sc_hd__clkbuf_16
X_35297_ _35743_/CLK _35297_/D VGND VGND VPWR VPWR _35297_/Q sky130_fd_sc_hd__dfxtp_1
X_25050_ input11/X VGND VGND VPWR VPWR _25050_/X sky130_fd_sc_hd__clkbuf_4
X_34248_ _34312_/CLK _34248_/D VGND VGND VPWR VPWR _34248_/Q sky130_fd_sc_hd__dfxtp_1
X_22262_ _32507_/Q _32379_/Q _32059_/Q _36027_/Q _22229_/X _22017_/X VGND VGND VPWR
+ VPWR _22262_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24001_ _24001_/A VGND VGND VPWR VPWR _32538_/D sky130_fd_sc_hd__clkbuf_1
X_21213_ _33181_/Q _32541_/Q _35933_/Q _35869_/Q _20968_/X _20969_/X VGND VGND VPWR
+ VPWR _21213_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22193_ _32761_/Q _32697_/Q _32633_/Q _36089_/Q _21872_/X _22009_/X VGND VGND VPWR
+ VPWR _22193_/X sky130_fd_sc_hd__mux4_1
X_34179_ _34243_/CLK _34179_/D VGND VGND VPWR VPWR _34179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21144_ _22556_/A VGND VGND VPWR VPWR _21144_/X sky130_fd_sc_hd__buf_4
XFILLER_105_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28740_ _28740_/A VGND VGND VPWR VPWR _34683_/D sky130_fd_sc_hd__clkbuf_1
X_25952_ _25952_/A VGND VGND VPWR VPWR _33394_/D sky130_fd_sc_hd__clkbuf_1
X_21075_ _20888_/X _21073_/X _21074_/X _20891_/X VGND VGND VPWR VPWR _21075_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20026_ _20146_/A VGND VGND VPWR VPWR _20026_/X sky130_fd_sc_hd__buf_4
XFILLER_150_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24903_ _24903_/A VGND VGND VPWR VPWR _32932_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28671_ _28671_/A VGND VGND VPWR VPWR _34650_/D sky130_fd_sc_hd__clkbuf_1
X_25883_ _25883_/A VGND VGND VPWR VPWR _33361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_918 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24834_ _23047_/X _32900_/Q _24844_/S VGND VGND VPWR VPWR _24835_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27622_ _27622_/A VGND VGND VPWR VPWR _34153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27553_ _27008_/X _34122_/Q _27559_/S VGND VGND VPWR VPWR _27554_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24765_ _22945_/X _32867_/Q _24781_/S VGND VGND VPWR VPWR _24766_/A sky130_fd_sc_hd__mux2_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21977_ _21971_/X _21976_/X _21728_/X VGND VGND VPWR VPWR _21999_/A sky130_fd_sc_hd__o21ba_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26504_ _25122_/X _33656_/Q _26518_/S VGND VGND VPWR VPWR _26505_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23716_ _23716_/A VGND VGND VPWR VPWR _32404_/D sky130_fd_sc_hd__clkbuf_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20928_ _20888_/X _20926_/X _20927_/X _20891_/X VGND VGND VPWR VPWR _20928_/X sky130_fd_sc_hd__a22o_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27484_ _26906_/X _34089_/Q _27488_/S VGND VGND VPWR VPWR _27485_/A sky130_fd_sc_hd__mux2_1
X_24696_ _24696_/A VGND VGND VPWR VPWR _32835_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29223_ _34885_/Q _29222_/X _29235_/S VGND VGND VPWR VPWR _29224_/A sky130_fd_sc_hd__mux2_1
X_26435_ _26435_/A VGND VGND VPWR VPWR _33623_/D sky130_fd_sc_hd__clkbuf_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23647_ _23647_/A VGND VGND VPWR VPWR _32373_/D sky130_fd_sc_hd__clkbuf_1
X_20859_ _35539_/Q _35475_/Q _35411_/Q _35347_/Q _20791_/X _20792_/X VGND VGND VPWR
+ VPWR _20859_/X sky130_fd_sc_hd__mux4_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29154_ input27/X VGND VGND VPWR VPWR _29154_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_35_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26366_ _26366_/A VGND VGND VPWR VPWR _33590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23578_ _23578_/A VGND VGND VPWR VPWR _32340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28105_ _26821_/X _34382_/Q _28123_/S VGND VGND VPWR VPWR _28106_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_812 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25317_ _25317_/A VGND VGND VPWR VPWR _33098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22529_ _35330_/Q _35266_/Q _35202_/Q _32322_/Q _22312_/X _22313_/X VGND VGND VPWR
+ VPWR _22529_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29085_ _29085_/A VGND VGND VPWR VPWR _34840_/D sky130_fd_sc_hd__clkbuf_1
X_26297_ _25016_/X _33558_/Q _26299_/S VGND VGND VPWR VPWR _26298_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _34074_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16050_ _17762_/A VGND VGND VPWR VPWR _17995_/A sky130_fd_sc_hd__buf_12
X_28036_ _28036_/A VGND VGND VPWR VPWR _34349_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25248_ _25248_/A VGND VGND VPWR VPWR _33065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25179_ _25179_/A VGND VGND VPWR VPWR _33034_/D sky130_fd_sc_hd__clkbuf_1
X_29987_ _29987_/A VGND VGND VPWR VPWR _35243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19740_ _19740_/A VGND VGND VPWR VPWR _32116_/D sky130_fd_sc_hd__buf_2
XFILLER_173_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28938_ _34777_/Q _24280_/X _28954_/S VGND VGND VPWR VPWR _28939_/A sky130_fd_sc_hd__mux2_1
X_16952_ _16948_/X _16951_/X _16775_/X VGND VGND VPWR VPWR _16976_/A sky130_fd_sc_hd__o21ba_1
XFILLER_238_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19671_ _19495_/X _19669_/X _19670_/X _19500_/X VGND VGND VPWR VPWR _19671_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16883_ _33509_/Q _33445_/Q _33381_/Q _33317_/Q _16770_/X _16771_/X VGND VGND VPWR
+ VPWR _16883_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28869_ _28869_/A VGND VGND VPWR VPWR _34744_/D sky130_fd_sc_hd__clkbuf_1
X_18622_ _32469_/Q _32341_/Q _32021_/Q _35989_/Q _18517_/X _20163_/A VGND VGND VPWR
+ VPWR _18622_/X sky130_fd_sc_hd__mux4_1
X_30900_ _30900_/A VGND VGND VPWR VPWR _35675_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31880_ _23237_/X _36140_/Q _31898_/S VGND VGND VPWR VPWR _31881_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18553_ _18549_/X _18552_/X _18340_/X _18342_/X VGND VGND VPWR VPWR _18570_/B sky130_fd_sc_hd__o211a_2
X_30831_ _23286_/X _35643_/Q _30839_/S VGND VGND VPWR VPWR _30832_/A sky130_fd_sc_hd__mux2_1
XTAP_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17504_ _35318_/Q _35254_/Q _35190_/Q _32310_/Q _17359_/X _17360_/X VGND VGND VPWR
+ VPWR _17504_/X sky130_fd_sc_hd__mux4_1
X_33550_ _35277_/CLK _33550_/D VGND VGND VPWR VPWR _33550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18484_ _32465_/Q _32337_/Q _32017_/Q _35985_/Q _18328_/X _20163_/A VGND VGND VPWR
+ VPWR _18484_/X sky130_fd_sc_hd__mux4_1
X_30762_ _23124_/X _35610_/Q _30776_/S VGND VGND VPWR VPWR _30763_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_460 _31991_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_471 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32501_ _33013_/CLK _32501_/D VGND VGND VPWR VPWR _32501_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17435_ _34548_/Q _32436_/Q _34420_/Q _34356_/Q _17225_/X _17226_/X VGND VGND VPWR
+ VPWR _17435_/X sky130_fd_sc_hd__mux4_1
XANTENNA_482 _31994_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33481_ _33545_/CLK _33481_/D VGND VGND VPWR VPWR _33481_/Q sky130_fd_sc_hd__dfxtp_1
X_30693_ _30693_/A VGND VGND VPWR VPWR _35577_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_493 _31994_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35220_ _35284_/CLK _35220_/D VGND VGND VPWR VPWR _35220_/Q sky130_fd_sc_hd__dfxtp_1
X_32432_ _35758_/CLK _32432_/D VGND VGND VPWR VPWR _32432_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_18 _32115_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_29 _32116_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17366_ _17362_/X _17365_/X _17161_/X VGND VGND VPWR VPWR _17367_/D sky130_fd_sc_hd__o21ba_1
XFILLER_144_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_20__f_CLK clkbuf_5_10_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_20__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_19105_ _35042_/Q _34978_/Q _34914_/Q _34850_/Q _19103_/X _19104_/X VGND VGND VPWR
+ VPWR _19105_/X sky130_fd_sc_hd__mux4_1
X_16317_ _16143_/X _16313_/X _16316_/X _16146_/X VGND VGND VPWR VPWR _16317_/X sky130_fd_sc_hd__a22o_1
X_35151_ _35215_/CLK _35151_/D VGND VGND VPWR VPWR _35151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17297_ _17297_/A _17297_/B _17297_/C _17297_/D VGND VGND VPWR VPWR _17298_/A sky130_fd_sc_hd__or4_4
X_32363_ _35242_/CLK _32363_/D VGND VGND VPWR VPWR _32363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _34080_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_220_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34102_ _36150_/CLK _34102_/D VGND VGND VPWR VPWR _34102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16248_ _33235_/Q _36115_/Q _33107_/Q _33043_/Q _16020_/X _16021_/X VGND VGND VPWR
+ VPWR _16248_/X sky130_fd_sc_hd__mux4_1
X_31314_ _35872_/Q input10/X _31316_/S VGND VGND VPWR VPWR _31315_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_1080 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19036_ _20256_/A VGND VGND VPWR VPWR _19036_/X sky130_fd_sc_hd__clkbuf_8
X_35082_ _35788_/CLK _35082_/D VGND VGND VPWR VPWR _35082_/Q sky130_fd_sc_hd__dfxtp_1
X_32294_ _35239_/CLK _32294_/D VGND VGND VPWR VPWR _32294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31245_ _31245_/A VGND VGND VPWR VPWR _35839_/D sky130_fd_sc_hd__clkbuf_1
Xoutput103 _31971_/Q VGND VGND VPWR VPWR D1[21] sky130_fd_sc_hd__buf_2
X_34033_ _34033_/CLK _34033_/D VGND VGND VPWR VPWR _34033_/Q sky130_fd_sc_hd__dfxtp_1
X_16179_ _16143_/X _16177_/X _16178_/X _16146_/X VGND VGND VPWR VPWR _16179_/X sky130_fd_sc_hd__a22o_1
Xoutput114 _31981_/Q VGND VGND VPWR VPWR D1[31] sky130_fd_sc_hd__buf_2
Xoutput125 _31991_/Q VGND VGND VPWR VPWR D1[41] sky130_fd_sc_hd__buf_2
XFILLER_126_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput136 _32001_/Q VGND VGND VPWR VPWR D1[51] sky130_fd_sc_hd__buf_2
XFILLER_217_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput147 _32011_/Q VGND VGND VPWR VPWR D1[61] sky130_fd_sc_hd__buf_2
XFILLER_142_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput158 _36187_/Q VGND VGND VPWR VPWR D2[13] sky130_fd_sc_hd__buf_2
X_31176_ _31176_/A VGND VGND VPWR VPWR _35806_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput169 _36197_/Q VGND VGND VPWR VPWR D2[23] sky130_fd_sc_hd__buf_2
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30127_ _30127_/A VGND VGND VPWR VPWR _35309_/D sky130_fd_sc_hd__clkbuf_1
X_19938_ _33210_/Q _32570_/Q _35962_/Q _35898_/Q _19727_/X _19728_/X VGND VGND VPWR
+ VPWR _19938_/X sky130_fd_sc_hd__mux4_1
X_35984_ _35984_/CLK _35984_/D VGND VGND VPWR VPWR _35984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30058_ _30058_/A VGND VGND VPWR VPWR _35277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34935_ _35257_/CLK _34935_/D VGND VGND VPWR VPWR _34935_/Q sky130_fd_sc_hd__dfxtp_1
X_19869_ _35768_/Q _35128_/Q _34488_/Q _33848_/Q _19793_/X _19794_/X VGND VGND VPWR
+ VPWR _19869_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21900_ _34289_/Q _34225_/Q _34161_/Q _34097_/Q _21689_/X _21690_/X VGND VGND VPWR
+ VPWR _21900_/X sky130_fd_sc_hd__mux4_1
X_22880_ _23075_/S VGND VGND VPWR VPWR _22908_/S sky130_fd_sc_hd__buf_4
XFILLER_110_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34866_ _34866_/CLK _34866_/D VGND VGND VPWR VPWR _34866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21831_ _21831_/A _21831_/B _21831_/C _21831_/D VGND VGND VPWR VPWR _21832_/A sky130_fd_sc_hd__or4_1
X_33817_ _35803_/CLK _33817_/D VGND VGND VPWR VPWR _33817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34797_ _34797_/CLK _34797_/D VGND VGND VPWR VPWR _34797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_984 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24550_ _24577_/S VGND VGND VPWR VPWR _24569_/S sky130_fd_sc_hd__clkbuf_8
X_33748_ _34259_/CLK _33748_/D VGND VGND VPWR VPWR _33748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21762_ _21753_/X _21760_/X _21761_/X VGND VGND VPWR VPWR _21763_/D sky130_fd_sc_hd__o21ba_1
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23501_ _22988_/X _32305_/Q _23509_/S VGND VGND VPWR VPWR _23502_/A sky130_fd_sc_hd__mux2_1
X_20713_ _32719_/Q _32655_/Q _32591_/Q _36047_/Q _22462_/A _22313_/A VGND VGND VPWR
+ VPWR _20713_/X sky130_fd_sc_hd__mux4_1
XFILLER_212_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24481_ _22932_/X _32735_/Q _24485_/S VGND VGND VPWR VPWR _24482_/A sky130_fd_sc_hd__mux2_1
X_33679_ _35341_/CLK _33679_/D VGND VGND VPWR VPWR _33679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21693_ _33515_/Q _33451_/Q _33387_/Q _33323_/Q _21370_/X _21371_/X VGND VGND VPWR
+ VPWR _21693_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26220_ _26220_/A VGND VGND VPWR VPWR _33521_/D sky130_fd_sc_hd__clkbuf_1
X_23432_ _22886_/X _32272_/Q _23446_/S VGND VGND VPWR VPWR _23433_/A sky130_fd_sc_hd__mux2_1
X_35418_ _35929_/CLK _35418_/D VGND VGND VPWR VPWR _35418_/Q sky130_fd_sc_hd__dfxtp_1
X_20644_ _22455_/A VGND VGND VPWR VPWR _20644_/X sky130_fd_sc_hd__buf_4
X_26151_ _26151_/A VGND VGND VPWR VPWR _33488_/D sky130_fd_sc_hd__clkbuf_1
X_35349_ _35925_/CLK _35349_/D VGND VGND VPWR VPWR _35349_/Q sky130_fd_sc_hd__dfxtp_1
X_23363_ _32241_/Q _23253_/X _23371_/S VGND VGND VPWR VPWR _23364_/A sky130_fd_sc_hd__mux2_1
X_20575_ input73/X input74/X VGND VGND VPWR VPWR _22361_/A sky130_fd_sc_hd__nor2b_4
XFILLER_20_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25102_ _25102_/A VGND VGND VPWR VPWR _33009_/D sky130_fd_sc_hd__clkbuf_1
X_22314_ _35324_/Q _35260_/Q _35196_/Q _32316_/Q _22312_/X _22313_/X VGND VGND VPWR
+ VPWR _22314_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26082_ _25097_/X _33456_/Q _26092_/S VGND VGND VPWR VPWR _26083_/A sky130_fd_sc_hd__mux2_1
X_23294_ input42/X VGND VGND VPWR VPWR _23294_/X sky130_fd_sc_hd__buf_4
XFILLER_11_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29910_ _35207_/Q _29228_/X _29914_/S VGND VGND VPWR VPWR _29911_/A sky130_fd_sc_hd__mux2_1
X_25033_ _25032_/X _32987_/Q _25051_/S VGND VGND VPWR VPWR _25034_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22245_ _22102_/X _22243_/X _22244_/X _22105_/X VGND VGND VPWR VPWR _22245_/X sky130_fd_sc_hd__a22o_1
XFILLER_191_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29841_ _35174_/Q _29126_/X _29851_/S VGND VGND VPWR VPWR _29842_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22176_ _35320_/Q _35256_/Q _35192_/Q _32312_/Q _21959_/X _21960_/X VGND VGND VPWR
+ VPWR _22176_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21127_ _33755_/Q _33691_/Q _33627_/Q _33563_/Q _21090_/X _21091_/X VGND VGND VPWR
+ VPWR _21127_/X sky130_fd_sc_hd__mux4_1
X_29772_ _29772_/A VGND VGND VPWR VPWR _35141_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26984_ input48/X VGND VGND VPWR VPWR _26984_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_247_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28723_ _28723_/A VGND VGND VPWR VPWR _34675_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21058_ _21058_/A VGND VGND VPWR VPWR _36184_/D sky130_fd_sc_hd__clkbuf_1
X_25935_ _25935_/A VGND VGND VPWR VPWR _33386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20009_ _20005_/X _20006_/X _20007_/X _20008_/X VGND VGND VPWR VPWR _20009_/X sky130_fd_sc_hd__a22o_1
XFILLER_235_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25866_ _25177_/X _33354_/Q _25872_/S VGND VGND VPWR VPWR _25867_/A sky130_fd_sc_hd__mux2_1
X_28654_ _28654_/A VGND VGND VPWR VPWR _34642_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24817_ _23022_/X _32892_/Q _24823_/S VGND VGND VPWR VPWR _24818_/A sky130_fd_sc_hd__mux2_1
X_27605_ _27605_/A VGND VGND VPWR VPWR _34145_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25797_ _25075_/X _33321_/Q _25801_/S VGND VGND VPWR VPWR _25798_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28585_ _26934_/X _34610_/Q _28591_/S VGND VGND VPWR VPWR _28586_/A sky130_fd_sc_hd__mux2_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27536_ _27536_/A VGND VGND VPWR VPWR _34113_/D sky130_fd_sc_hd__clkbuf_1
X_24748_ _22920_/X _32859_/Q _24760_/S VGND VGND VPWR VPWR _24749_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27467_ _26881_/X _34081_/Q _27467_/S VGND VGND VPWR VPWR _27468_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_959 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24679_ _24679_/A VGND VGND VPWR VPWR _32827_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29206_ input46/X VGND VGND VPWR VPWR _29206_/X sky130_fd_sc_hd__buf_4
X_17220_ _16999_/X _17218_/X _17219_/X _17002_/X VGND VGND VPWR VPWR _17220_/X sky130_fd_sc_hd__a22o_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26418_ _24995_/X _33615_/Q _26434_/S VGND VGND VPWR VPWR _26419_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27398_ _34048_/Q _24400_/X _27416_/S VGND VGND VPWR VPWR _27399_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17151_ _35308_/Q _35244_/Q _35180_/Q _32300_/Q _17006_/X _17007_/X VGND VGND VPWR
+ VPWR _17151_/X sky130_fd_sc_hd__mux4_1
X_29137_ _29137_/A VGND VGND VPWR VPWR _34857_/D sky130_fd_sc_hd__clkbuf_1
X_26349_ _26349_/A VGND VGND VPWR VPWR _33582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput16 DW[23] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__buf_4
Xinput27 DW[33] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__buf_4
X_16102_ _16102_/A _16102_/B _16102_/C _16102_/D VGND VGND VPWR VPWR _16103_/A sky130_fd_sc_hd__or4_4
XFILLER_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput38 DW[43] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__buf_4
X_29068_ _34835_/Q _29067_/X _29080_/S VGND VGND VPWR VPWR _29069_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput49 DW[53] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__buf_8
X_17082_ _34538_/Q _32426_/Q _34410_/Q _34346_/Q _16872_/X _16873_/X VGND VGND VPWR
+ VPWR _17082_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16033_ _17829_/A VGND VGND VPWR VPWR _16033_/X sky130_fd_sc_hd__buf_4
XFILLER_157_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28019_ _28019_/A VGND VGND VPWR VPWR _34341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31030_ _35737_/Q _29086_/X _31046_/S VGND VGND VPWR VPWR _31031_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_948 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17984_ _33028_/Q _32964_/Q _32900_/Q _32836_/Q _17695_/X _17696_/X VGND VGND VPWR
+ VPWR _17984_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19723_ _35828_/Q _32206_/Q _35700_/Q _35636_/Q _19613_/X _19614_/X VGND VGND VPWR
+ VPWR _19723_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16935_ _17994_/A VGND VGND VPWR VPWR _16935_/X sky130_fd_sc_hd__buf_6
X_32981_ _32983_/CLK _32981_/D VGND VGND VPWR VPWR _32981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34720_ _35098_/CLK _34720_/D VGND VGND VPWR VPWR _34720_/Q sky130_fd_sc_hd__dfxtp_1
X_31932_ _23319_/X _36165_/Q _31940_/S VGND VGND VPWR VPWR _31933_/A sky130_fd_sc_hd__mux2_1
X_19654_ _33202_/Q _32562_/Q _35954_/Q _35890_/Q _19374_/X _19375_/X VGND VGND VPWR
+ VPWR _19654_/X sky130_fd_sc_hd__mux4_1
X_16866_ _33188_/Q _32548_/Q _35940_/Q _35876_/Q _16721_/X _16722_/X VGND VGND VPWR
+ VPWR _16866_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_7_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _35293_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_237_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18605_ _35028_/Q _34964_/Q _34900_/Q _34836_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _18605_/X sky130_fd_sc_hd__mux4_1
X_34651_ _36201_/CLK _34651_/D VGND VGND VPWR VPWR _34651_/Q sky130_fd_sc_hd__dfxtp_1
X_19585_ _33200_/Q _32560_/Q _35952_/Q _35888_/Q _19374_/X _19375_/X VGND VGND VPWR
+ VPWR _19585_/X sky130_fd_sc_hd__mux4_1
X_31863_ _23175_/X _36132_/Q _31877_/S VGND VGND VPWR VPWR _31864_/A sky130_fd_sc_hd__mux2_1
X_16797_ _34786_/Q _34722_/Q _34658_/Q _34594_/Q _16582_/X _16583_/X VGND VGND VPWR
+ VPWR _16797_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33602_ _33795_/CLK _33602_/D VGND VGND VPWR VPWR _33602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18536_ _18387_/X _18534_/X _18535_/X _18397_/X VGND VGND VPWR VPWR _18536_/X sky130_fd_sc_hd__a22o_1
X_30814_ _23261_/X _35635_/Q _30818_/S VGND VGND VPWR VPWR _30815_/A sky130_fd_sc_hd__mux2_1
X_34582_ _35286_/CLK _34582_/D VGND VGND VPWR VPWR _34582_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31794_ _31794_/A VGND VGND VPWR VPWR _36099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33533_ _33789_/CLK _33533_/D VGND VGND VPWR VPWR _33533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30745_ _23099_/X _35602_/Q _30755_/S VGND VGND VPWR VPWR _30746_/A sky130_fd_sc_hd__mux2_1
X_18467_ _19173_/A VGND VGND VPWR VPWR _18467_/X sky130_fd_sc_hd__buf_6
XANTENNA_290 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17418_ _32500_/Q _32372_/Q _32052_/Q _36020_/Q _17276_/X _17417_/X VGND VGND VPWR
+ VPWR _17418_/X sky130_fd_sc_hd__mux4_1
X_33464_ _34297_/CLK _33464_/D VGND VGND VPWR VPWR _33464_/Q sky130_fd_sc_hd__dfxtp_1
X_18398_ _18387_/X _18391_/X _18395_/X _18397_/X VGND VGND VPWR VPWR _18398_/X sky130_fd_sc_hd__a22o_1
X_30676_ _30676_/A VGND VGND VPWR VPWR _35569_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35203_ _35331_/CLK _35203_/D VGND VGND VPWR VPWR _35203_/Q sky130_fd_sc_hd__dfxtp_1
X_32415_ _35296_/CLK _32415_/D VGND VGND VPWR VPWR _32415_/Q sky130_fd_sc_hd__dfxtp_1
X_36183_ _36202_/CLK _36183_/D VGND VGND VPWR VPWR _36183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17349_ _35762_/Q _35122_/Q _34482_/Q _33842_/Q _17140_/X _17141_/X VGND VGND VPWR
+ VPWR _17349_/X sky130_fd_sc_hd__mux4_1
X_33395_ _33779_/CLK _33395_/D VGND VGND VPWR VPWR _33395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35134_ _35711_/CLK _35134_/D VGND VGND VPWR VPWR _35134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20360_ _35078_/Q _35014_/Q _34950_/Q _34886_/Q _20162_/X _20163_/X VGND VGND VPWR
+ VPWR _20360_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32346_ _32860_/CLK _32346_/D VGND VGND VPWR VPWR _32346_/Q sky130_fd_sc_hd__dfxtp_1
X_19019_ _18941_/X _19017_/X _19018_/X _18944_/X VGND VGND VPWR VPWR _19019_/X sky130_fd_sc_hd__a22o_1
X_20291_ _33220_/Q _32580_/Q _35972_/Q _35908_/Q _20080_/X _20081_/X VGND VGND VPWR
+ VPWR _20291_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35065_ _35386_/CLK _35065_/D VGND VGND VPWR VPWR _35065_/Q sky130_fd_sc_hd__dfxtp_1
X_32277_ _36202_/CLK _32277_/D VGND VGND VPWR VPWR _32277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22030_ _21952_/X _22026_/X _22029_/X _21955_/X VGND VGND VPWR VPWR _22030_/X sky130_fd_sc_hd__a22o_1
X_34016_ _34016_/CLK _34016_/D VGND VGND VPWR VPWR _34016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31228_ _35831_/Q input36/X _31244_/S VGND VGND VPWR VPWR _31229_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31159_ _31159_/A VGND VGND VPWR VPWR _35798_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23981_ _22889_/X _32529_/Q _23993_/S VGND VGND VPWR VPWR _23982_/A sky130_fd_sc_hd__mux2_1
X_35967_ _35970_/CLK _35967_/D VGND VGND VPWR VPWR _35967_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25720_ _25720_/A VGND VGND VPWR VPWR _33285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22932_ input9/X VGND VGND VPWR VPWR _22932_/X sky130_fd_sc_hd__clkbuf_4
X_34918_ _35942_/CLK _34918_/D VGND VGND VPWR VPWR _34918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35898_ _36027_/CLK _35898_/D VGND VGND VPWR VPWR _35898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25651_ _25651_/A VGND VGND VPWR VPWR _33252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22863_ _33229_/Q _32589_/Q _35981_/Q _35917_/Q _20675_/X _20676_/X VGND VGND VPWR
+ VPWR _22863_/X sky130_fd_sc_hd__mux4_1
X_34849_ _35040_/CLK _34849_/D VGND VGND VPWR VPWR _34849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24602_ _22907_/X _32791_/Q _24602_/S VGND VGND VPWR VPWR _24603_/A sky130_fd_sc_hd__mux2_1
X_28370_ _28370_/A VGND VGND VPWR VPWR _34508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21814_ _21810_/X _21813_/X _21736_/X _21737_/X VGND VGND VPWR VPWR _21831_/B sky130_fd_sc_hd__o211a_1
X_25582_ _25582_/A VGND VGND VPWR VPWR _33221_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22794_ _21749_/A _22792_/X _22793_/X _21752_/A VGND VGND VPWR VPWR _22794_/X sky130_fd_sc_hd__a22o_1
XFILLER_225_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27321_ _27321_/A VGND VGND VPWR VPWR _34011_/D sky130_fd_sc_hd__clkbuf_1
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24533_ _24533_/A VGND VGND VPWR VPWR _32759_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21745_ _33196_/Q _32556_/Q _35948_/Q _35884_/Q _21674_/X _21675_/X VGND VGND VPWR
+ VPWR _21745_/X sky130_fd_sc_hd__mux4_1
XPHY_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27252_ _26962_/X _33979_/Q _27260_/S VGND VGND VPWR VPWR _27253_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24464_ _22907_/X _32727_/Q _24464_/S VGND VGND VPWR VPWR _24465_/A sky130_fd_sc_hd__mux2_1
X_21676_ _33194_/Q _32554_/Q _35946_/Q _35882_/Q _21674_/X _21675_/X VGND VGND VPWR
+ VPWR _21676_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26203_ _26203_/A VGND VGND VPWR VPWR _33513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23415_ _32266_/Q _23336_/X _23421_/S VGND VGND VPWR VPWR _23416_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20627_ _20657_/A VGND VGND VPWR VPWR _22582_/A sky130_fd_sc_hd__buf_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27183_ _26860_/X _33946_/Q _27197_/S VGND VGND VPWR VPWR _27184_/A sky130_fd_sc_hd__mux2_1
X_24395_ _32702_/Q _24394_/X _24398_/S VGND VGND VPWR VPWR _24396_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26134_ _25174_/X _33481_/Q _26134_/S VGND VGND VPWR VPWR _26135_/A sky130_fd_sc_hd__mux2_1
X_23346_ _32233_/Q _23345_/X _23346_/S VGND VGND VPWR VPWR _23347_/A sky130_fd_sc_hd__mux2_1
X_20558_ _20554_/X _20557_/X _20142_/A _20143_/A VGND VGND VPWR VPWR _20573_/B sky130_fd_sc_hd__o211a_1
XFILLER_164_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26065_ _25072_/X _33448_/Q _26071_/S VGND VGND VPWR VPWR _26066_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23277_ input37/X VGND VGND VPWR VPWR _23277_/X sky130_fd_sc_hd__buf_4
X_20489_ _34059_/Q _33995_/Q _33931_/Q _32267_/Q _18358_/X _18360_/X VGND VGND VPWR
+ VPWR _20489_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25016_ input63/X VGND VGND VPWR VPWR _25016_/X sky130_fd_sc_hd__buf_6
X_22228_ _22008_/X _22226_/X _22227_/X _22014_/X VGND VGND VPWR VPWR _22228_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29824_ _35166_/Q _29101_/X _29830_/S VGND VGND VPWR VPWR _29825_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22159_ _22155_/X _22156_/X _22157_/X _22158_/X VGND VGND VPWR VPWR _22159_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29755_ _29755_/A VGND VGND VPWR VPWR _35133_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26967_ _26967_/A VGND VGND VPWR VPWR _33852_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16720_ _35552_/Q _35488_/Q _35424_/Q _35360_/Q _16544_/X _16545_/X VGND VGND VPWR
+ VPWR _16720_/X sky130_fd_sc_hd__mux4_1
X_28706_ _28706_/A VGND VGND VPWR VPWR _34667_/D sky130_fd_sc_hd__clkbuf_1
X_25918_ _25053_/X _33378_/Q _25936_/S VGND VGND VPWR VPWR _25919_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29686_ _29686_/A VGND VGND VPWR VPWR _35100_/D sky130_fd_sc_hd__clkbuf_1
X_26898_ _26897_/X _33830_/Q _26913_/S VGND VGND VPWR VPWR _26899_/A sky130_fd_sc_hd__mux2_1
XFILLER_247_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28637_ _27011_/X _34635_/Q _28641_/S VGND VGND VPWR VPWR _28638_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16651_ _16645_/X _16650_/X _16441_/X VGND VGND VPWR VPWR _16661_/C sky130_fd_sc_hd__o21ba_1
XFILLER_78_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25849_ _25849_/A VGND VGND VPWR VPWR _33345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19370_ _35818_/Q _32195_/Q _35690_/Q _35626_/Q _19260_/X _19261_/X VGND VGND VPWR
+ VPWR _19370_/X sky130_fd_sc_hd__mux4_1
X_16582_ _17994_/A VGND VGND VPWR VPWR _16582_/X sky130_fd_sc_hd__buf_6
X_28568_ _26909_/X _34602_/Q _28570_/S VGND VGND VPWR VPWR _28569_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18321_ _20203_/A VGND VGND VPWR VPWR _18321_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_231_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27519_ _27519_/A VGND VGND VPWR VPWR _34105_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28499_ _28499_/A VGND VGND VPWR VPWR _34569_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ _32781_/Q _32717_/Q _32653_/Q _36109_/Q _17978_/X _16873_/A VGND VGND VPWR
+ VPWR _18252_/X sky130_fd_sc_hd__mux4_1
XFILLER_188_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30530_ _23237_/X _35500_/Q _30548_/S VGND VGND VPWR VPWR _30531_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17203_ _33518_/Q _33454_/Q _33390_/Q _33326_/Q _17123_/X _17124_/X VGND VGND VPWR
+ VPWR _17203_/X sky130_fd_sc_hd__mux4_1
X_30461_ _23342_/X _35468_/Q _30463_/S VGND VGND VPWR VPWR _30462_/A sky130_fd_sc_hd__mux2_1
X_18183_ _18183_/A _18183_/B _18183_/C _18183_/D VGND VGND VPWR VPWR _18184_/A sky130_fd_sc_hd__or4_4
XFILLER_30_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32200_ _35951_/CLK _32200_/D VGND VGND VPWR VPWR _32200_/Q sky130_fd_sc_hd__dfxtp_1
X_17134_ _33004_/Q _32940_/Q _32876_/Q _32812_/Q _16989_/X _16990_/X VGND VGND VPWR
+ VPWR _17134_/X sky130_fd_sc_hd__mux4_1
X_30392_ _23234_/X _35435_/Q _30392_/S VGND VGND VPWR VPWR _30393_/A sky130_fd_sc_hd__mux2_1
X_33180_ _35928_/CLK _33180_/D VGND VGND VPWR VPWR _33180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_7_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_7_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_7_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32131_ _35750_/CLK _32131_/D VGND VGND VPWR VPWR _32131_/Q sky130_fd_sc_hd__dfxtp_1
X_17065_ _32490_/Q _32362_/Q _32042_/Q _36010_/Q _16923_/X _17064_/X VGND VGND VPWR
+ VPWR _17065_/X sky130_fd_sc_hd__mux4_1
XFILLER_170_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16016_ _17978_/A VGND VGND VPWR VPWR _17862_/A sky130_fd_sc_hd__buf_12
X_32062_ _36033_/CLK _32062_/D VGND VGND VPWR VPWR _32062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31013_ _35729_/Q _29061_/X _31025_/S VGND VGND VPWR VPWR _31014_/A sky130_fd_sc_hd__mux2_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35821_ _35885_/CLK _35821_/D VGND VGND VPWR VPWR _35821_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _17860_/X _17965_/X _17966_/X _17865_/X VGND VGND VPWR VPWR _17967_/X sky130_fd_sc_hd__a22o_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19706_ _19502_/X _19704_/X _19705_/X _19505_/X VGND VGND VPWR VPWR _19706_/X sky130_fd_sc_hd__a22o_1
XFILLER_239_985 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35752_ _35879_/CLK _35752_/D VGND VGND VPWR VPWR _35752_/Q sky130_fd_sc_hd__dfxtp_1
X_16918_ _16914_/X _16917_/X _16775_/X VGND VGND VPWR VPWR _16944_/A sky130_fd_sc_hd__o21ba_1
XFILLER_211_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32964_ _36100_/CLK _32964_/D VGND VGND VPWR VPWR _32964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17898_ _17894_/X _17897_/X _17867_/X VGND VGND VPWR VPWR _17899_/D sky130_fd_sc_hd__o21ba_1
XFILLER_238_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34703_ _35215_/CLK _34703_/D VGND VGND VPWR VPWR _34703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31915_ _23294_/X _36157_/Q _31919_/S VGND VGND VPWR VPWR _31916_/A sky130_fd_sc_hd__mux2_1
X_19637_ _19633_/X _19636_/X _19428_/X VGND VGND VPWR VPWR _19667_/A sky130_fd_sc_hd__o21ba_1
XFILLER_93_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35683_ _35811_/CLK _35683_/D VGND VGND VPWR VPWR _35683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16849_ _17908_/A VGND VGND VPWR VPWR _16849_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_214_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32895_ _32959_/CLK _32895_/D VGND VGND VPWR VPWR _32895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34634_ _35338_/CLK _34634_/D VGND VGND VPWR VPWR _34634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_871 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19568_ _33520_/Q _33456_/Q _33392_/Q _33328_/Q _19423_/X _19424_/X VGND VGND VPWR
+ VPWR _19568_/X sky130_fd_sc_hd__mux4_1
X_31846_ _23130_/X _36124_/Q _31856_/S VGND VGND VPWR VPWR _31847_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18519_ _32978_/Q _32914_/Q _32850_/Q _32786_/Q _18333_/X _18335_/X VGND VGND VPWR
+ VPWR _18519_/X sky130_fd_sc_hd__mux4_1
X_34565_ _35779_/CLK _34565_/D VGND VGND VPWR VPWR _34565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31777_ _31777_/A VGND VGND VPWR VPWR _36091_/D sky130_fd_sc_hd__clkbuf_1
X_19499_ _34286_/Q _34222_/Q _34158_/Q _34094_/Q _19389_/X _19390_/X VGND VGND VPWR
+ VPWR _19499_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21530_ _21241_/X _21528_/X _21529_/X _21244_/X VGND VGND VPWR VPWR _21530_/X sky130_fd_sc_hd__a22o_1
X_33516_ _34293_/CLK _33516_/D VGND VGND VPWR VPWR _33516_/Q sky130_fd_sc_hd__dfxtp_1
X_30728_ _30728_/A VGND VGND VPWR VPWR _35594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34496_ _35777_/CLK _34496_/D VGND VGND VPWR VPWR _34496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36235_ _36237_/CLK _36235_/D VGND VGND VPWR VPWR _36235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33447_ _35991_/CLK _33447_/D VGND VGND VPWR VPWR _33447_/Q sky130_fd_sc_hd__dfxtp_1
X_21461_ _21457_/X _21460_/X _21383_/X _21384_/X VGND VGND VPWR VPWR _21478_/B sky130_fd_sc_hd__o211a_1
X_30659_ _30659_/A VGND VGND VPWR VPWR _35561_/D sky130_fd_sc_hd__clkbuf_1
X_23200_ _32182_/Q _23199_/X _23350_/S VGND VGND VPWR VPWR _23201_/A sky130_fd_sc_hd__mux2_1
X_20412_ _35592_/Q _35528_/Q _35464_/Q _35400_/Q _20256_/X _20257_/X VGND VGND VPWR
+ VPWR _20412_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36166_ _36166_/CLK _36166_/D VGND VGND VPWR VPWR _36166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24180_ _22982_/X _32623_/Q _24192_/S VGND VGND VPWR VPWR _24181_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33378_ _33635_/CLK _33378_/D VGND VGND VPWR VPWR _33378_/Q sky130_fd_sc_hd__dfxtp_1
X_21392_ _33186_/Q _32546_/Q _35938_/Q _35874_/Q _21321_/X _21322_/X VGND VGND VPWR
+ VPWR _21392_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35117_ _35564_/CLK _35117_/D VGND VGND VPWR VPWR _35117_/Q sky130_fd_sc_hd__dfxtp_1
X_23131_ _32156_/Q _23130_/X _23146_/S VGND VGND VPWR VPWR _23132_/A sky130_fd_sc_hd__mux2_1
X_32329_ _35273_/CLK _32329_/D VGND VGND VPWR VPWR _32329_/Q sky130_fd_sc_hd__dfxtp_1
X_20343_ _33286_/Q _36166_/Q _33158_/Q _33094_/Q _20064_/X _20065_/X VGND VGND VPWR
+ VPWR _20343_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36097_ _36097_/CLK _36097_/D VGND VGND VPWR VPWR _36097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23062_ input55/X VGND VGND VPWR VPWR _23062_/X sky130_fd_sc_hd__clkbuf_4
X_35048_ _35050_/CLK _35048_/D VGND VGND VPWR VPWR _35048_/Q sky130_fd_sc_hd__dfxtp_1
X_20274_ _33540_/Q _33476_/Q _33412_/Q _33348_/Q _20129_/X _20130_/X VGND VGND VPWR
+ VPWR _20274_/X sky130_fd_sc_hd__mux4_1
XTAP_6107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22013_ _33268_/Q _36148_/Q _33140_/Q _33076_/Q _22011_/X _22012_/X VGND VGND VPWR
+ VPWR _22013_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27870_ _34271_/Q _24298_/X _27874_/S VGND VGND VPWR VPWR _27871_/A sky130_fd_sc_hd__mux2_1
XTAP_5406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26821_ input1/X VGND VGND VPWR VPWR _26821_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1030 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29540_ _29540_/A VGND VGND VPWR VPWR _35031_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23964_ _23065_/X _32522_/Q _23970_/S VGND VGND VPWR VPWR _23965_/A sky130_fd_sc_hd__mux2_1
X_26752_ _26752_/A VGND VGND VPWR VPWR _33772_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25703_ _25703_/A VGND VGND VPWR VPWR _33277_/D sky130_fd_sc_hd__clkbuf_1
X_22915_ _22914_/X _32025_/Q _22939_/S VGND VGND VPWR VPWR _22916_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26683_ _25186_/X _33741_/Q _26683_/S VGND VGND VPWR VPWR _26684_/A sky130_fd_sc_hd__mux2_1
X_29471_ _29471_/A VGND VGND VPWR VPWR _34998_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23895_ _22963_/X _32489_/Q _23899_/S VGND VGND VPWR VPWR _23896_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28422_ _28422_/A VGND VGND VPWR VPWR _34532_/D sky130_fd_sc_hd__clkbuf_1
X_22846_ _34317_/Q _34253_/Q _34189_/Q _34125_/Q _20645_/X _20646_/X VGND VGND VPWR
+ VPWR _22846_/X sky130_fd_sc_hd__mux4_1
X_25634_ _25634_/A VGND VGND VPWR VPWR _33244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28353_ _34500_/Q _24413_/X _28363_/S VGND VGND VPWR VPWR _28354_/A sky130_fd_sc_hd__mux2_1
X_25565_ _25565_/A VGND VGND VPWR VPWR _33213_/D sky130_fd_sc_hd__clkbuf_1
X_22777_ _35338_/Q _35274_/Q _35210_/Q _32330_/Q _20688_/X _20690_/X VGND VGND VPWR
+ VPWR _22777_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_240_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _34312_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_169_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27304_ _27304_/A VGND VGND VPWR VPWR _34003_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24516_ _24516_/A VGND VGND VPWR VPWR _32751_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21728_ _22434_/A VGND VGND VPWR VPWR _21728_/X sky130_fd_sc_hd__clkbuf_4
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28284_ _34467_/Q _24311_/X _28300_/S VGND VGND VPWR VPWR _28285_/A sky130_fd_sc_hd__mux2_1
X_25496_ _25496_/A VGND VGND VPWR VPWR _33180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24447_ _24447_/A VGND VGND VPWR VPWR _32718_/D sky130_fd_sc_hd__clkbuf_1
X_27235_ _26937_/X _33971_/Q _27239_/S VGND VGND VPWR VPWR _27236_/A sky130_fd_sc_hd__mux2_1
X_21659_ _22370_/A VGND VGND VPWR VPWR _21659_/X sky130_fd_sc_hd__buf_4
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27166_ _26835_/X _33938_/Q _27176_/S VGND VGND VPWR VPWR _27167_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24378_ _24378_/A VGND VGND VPWR VPWR _32696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26117_ _26117_/A VGND VGND VPWR VPWR _33472_/D sky130_fd_sc_hd__clkbuf_1
X_23329_ _23329_/A VGND VGND VPWR VPWR _32227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27097_ _27097_/A VGND VGND VPWR VPWR _33905_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26048_ _25047_/X _33440_/Q _26050_/S VGND VGND VPWR VPWR _26049_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18870_ _20282_/A VGND VGND VPWR VPWR _18870_/X sky130_fd_sc_hd__buf_6
XTAP_6630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17821_ _35071_/Q _35007_/Q _34943_/Q _34879_/Q _17509_/X _17510_/X VGND VGND VPWR
+ VPWR _17821_/X sky130_fd_sc_hd__mux4_1
X_29807_ _35158_/Q _29076_/X _29809_/S VGND VGND VPWR VPWR _29808_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27999_ _26866_/X _34332_/Q _28009_/S VGND VGND VPWR VPWR _28000_/A sky130_fd_sc_hd__mux2_1
XTAP_6696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17752_ _17752_/A _17752_/B _17752_/C _17752_/D VGND VGND VPWR VPWR _17753_/A sky130_fd_sc_hd__or4_2
X_29738_ _29738_/A VGND VGND VPWR VPWR _35125_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16703_ _17762_/A VGND VGND VPWR VPWR _16703_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_236_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29669_ _29669_/A VGND VGND VPWR VPWR _35092_/D sky130_fd_sc_hd__clkbuf_1
X_17683_ _17683_/A VGND VGND VPWR VPWR _31995_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31700_ _36055_/Q input64/X _31700_/S VGND VGND VPWR VPWR _31701_/A sky130_fd_sc_hd__mux2_1
X_19422_ _19142_/X _19420_/X _19421_/X _19147_/X VGND VGND VPWR VPWR _19422_/X sky130_fd_sc_hd__a22o_1
X_16634_ _16349_/X _16632_/X _16633_/X _16355_/X VGND VGND VPWR VPWR _16634_/X sky130_fd_sc_hd__a22o_1
X_32680_ _33255_/CLK _32680_/D VGND VGND VPWR VPWR _32680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31631_ _36022_/Q input35/X _31649_/S VGND VGND VPWR VPWR _31632_/A sky130_fd_sc_hd__mux2_1
X_19353_ _19149_/X _19351_/X _19352_/X _19152_/X VGND VGND VPWR VPWR _19353_/X sky130_fd_sc_hd__a22o_1
X_16565_ _16561_/X _16564_/X _16422_/X VGND VGND VPWR VPWR _16591_/A sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_231_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _36039_/CLK sky130_fd_sc_hd__clkbuf_16
X_18304_ _18357_/A VGND VGND VPWR VPWR _20256_/A sky130_fd_sc_hd__buf_12
X_34350_ _35052_/CLK _34350_/D VGND VGND VPWR VPWR _34350_/Q sky130_fd_sc_hd__dfxtp_1
X_31562_ _31562_/A VGND VGND VPWR VPWR _35989_/D sky130_fd_sc_hd__clkbuf_1
X_19284_ _19280_/X _19283_/X _19075_/X VGND VGND VPWR VPWR _19314_/A sky130_fd_sc_hd__o21ba_1
X_16496_ _17908_/A VGND VGND VPWR VPWR _16496_/X sky130_fd_sc_hd__buf_4
XFILLER_241_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33301_ _34001_/CLK _33301_/D VGND VGND VPWR VPWR _33301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18235_ _18231_/X _18234_/X _17853_/A VGND VGND VPWR VPWR _18243_/C sky130_fd_sc_hd__o21ba_1
X_30513_ _23175_/X _35492_/Q _30527_/S VGND VGND VPWR VPWR _30514_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34281_ _34281_/CLK _34281_/D VGND VGND VPWR VPWR _34281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31493_ _23267_/X _35957_/Q _31493_/S VGND VGND VPWR VPWR _31494_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36020_ _36149_/CLK _36020_/D VGND VGND VPWR VPWR _36020_/Q sky130_fd_sc_hd__dfxtp_1
X_33232_ _36114_/CLK _33232_/D VGND VGND VPWR VPWR _33232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18166_ _33034_/Q _32970_/Q _32906_/Q _32842_/Q _15980_/X _15983_/X VGND VGND VPWR
+ VPWR _18166_/X sky130_fd_sc_hd__mux4_1
X_30444_ _30444_/A VGND VGND VPWR VPWR _35459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17117_ _17113_/X _17116_/X _16808_/X VGND VGND VPWR VPWR _17118_/D sky130_fd_sc_hd__o21ba_1
X_33163_ _36172_/CLK _33163_/D VGND VGND VPWR VPWR _33163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18097_ _17901_/X _18095_/X _18096_/X _17906_/X VGND VGND VPWR VPWR _18097_/X sky130_fd_sc_hd__a22o_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30375_ _30375_/A VGND VGND VPWR VPWR _35426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32114_ _35555_/CLK _32114_/D VGND VGND VPWR VPWR _32114_/Q sky130_fd_sc_hd__dfxtp_1
X_17048_ _33770_/Q _33706_/Q _33642_/Q _33578_/Q _16843_/X _16844_/X VGND VGND VPWR
+ VPWR _17048_/X sky130_fd_sc_hd__mux4_1
X_33094_ _36166_/CLK _33094_/D VGND VGND VPWR VPWR _33094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_298_CLK clkbuf_6_50__f_CLK/X VGND VGND VPWR VPWR _35772_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32045_ _36013_/CLK _32045_/D VGND VGND VPWR VPWR _32045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1074 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18999_ _34016_/Q _33952_/Q _33888_/Q _32160_/Q _18967_/X _18968_/X VGND VGND VPWR
+ VPWR _18999_/X sky130_fd_sc_hd__mux4_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35804_ _35929_/CLK _35804_/D VGND VGND VPWR VPWR _35804_/Q sky130_fd_sc_hd__dfxtp_1
X_33996_ _34316_/CLK _33996_/D VGND VGND VPWR VPWR _33996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_960 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35735_ _35925_/CLK _35735_/D VGND VGND VPWR VPWR _35735_/Q sky130_fd_sc_hd__dfxtp_1
X_20961_ _22511_/A VGND VGND VPWR VPWR _20961_/X sky130_fd_sc_hd__buf_4
XFILLER_39_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32947_ _35765_/CLK _32947_/D VGND VGND VPWR VPWR _32947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22700_ _22508_/X _22698_/X _22699_/X _22511_/X VGND VGND VPWR VPWR _22700_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_470_CLK clkbuf_6_8__f_CLK/X VGND VGND VPWR VPWR _35811_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23680_ _32389_/Q _23319_/X _23688_/S VGND VGND VPWR VPWR _23681_/A sky130_fd_sc_hd__mux2_1
X_35666_ _35666_/CLK _35666_/D VGND VGND VPWR VPWR _35666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20892_ _20888_/X _20889_/X _20890_/X _20891_/X VGND VGND VPWR VPWR _20892_/X sky130_fd_sc_hd__a22o_1
X_32878_ _33007_/CLK _32878_/D VGND VGND VPWR VPWR _32878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22631_ _22460_/X _22629_/X _22630_/X _22465_/X VGND VGND VPWR VPWR _22631_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34617_ _34745_/CLK _34617_/D VGND VGND VPWR VPWR _34617_/Q sky130_fd_sc_hd__dfxtp_1
X_31829_ _23105_/X _36116_/Q _31835_/S VGND VGND VPWR VPWR _31830_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35597_ _35597_/CLK _35597_/D VGND VGND VPWR VPWR _35597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_222_CLK clkbuf_6_55__f_CLK/X VGND VGND VPWR VPWR _34562_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_224_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25350_ _25026_/X _33113_/Q _25366_/S VGND VGND VPWR VPWR _25351_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22562_ _34819_/Q _34755_/Q _34691_/Q _34627_/Q _22241_/X _22242_/X VGND VGND VPWR
+ VPWR _22562_/X sky130_fd_sc_hd__mux4_1
X_34548_ _34805_/CLK _34548_/D VGND VGND VPWR VPWR _34548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24301_ input10/X VGND VGND VPWR VPWR _24301_/X sky130_fd_sc_hd__buf_4
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21513_ _34278_/Q _34214_/Q _34150_/Q _34086_/Q _21336_/X _21337_/X VGND VGND VPWR
+ VPWR _21513_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25281_ _25125_/X _33081_/Q _25293_/S VGND VGND VPWR VPWR _25282_/A sky130_fd_sc_hd__mux2_1
X_22493_ _35329_/Q _35265_/Q _35201_/Q _32321_/Q _22312_/X _22313_/X VGND VGND VPWR
+ VPWR _22493_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34479_ _35822_/CLK _34479_/D VGND VGND VPWR VPWR _34479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27020_ _30329_/B _29049_/B _30329_/A VGND VGND VPWR VPWR _27426_/A sky130_fd_sc_hd__nor3b_4
X_36218_ _36220_/CLK _36218_/D VGND VGND VPWR VPWR _36218_/Q sky130_fd_sc_hd__dfxtp_1
X_24232_ _23059_/X _32648_/Q _24234_/S VGND VGND VPWR VPWR _24233_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21444_ _22503_/A VGND VGND VPWR VPWR _21444_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_147_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24163_ _22957_/X _32615_/Q _24171_/S VGND VGND VPWR VPWR _24164_/A sky130_fd_sc_hd__mux2_1
X_36149_ _36149_/CLK _36149_/D VGND VGND VPWR VPWR _36149_/Q sky130_fd_sc_hd__dfxtp_1
X_21375_ _22434_/A VGND VGND VPWR VPWR _21375_/X sky130_fd_sc_hd__buf_2
X_23114_ input64/X VGND VGND VPWR VPWR _23114_/X sky130_fd_sc_hd__buf_4
X_20326_ _34821_/Q _34757_/Q _34693_/Q _34629_/Q _20294_/X _20295_/X VGND VGND VPWR
+ VPWR _20326_/X sky130_fd_sc_hd__mux4_1
X_24094_ _23056_/X _32583_/Q _24098_/S VGND VGND VPWR VPWR _24095_/A sky130_fd_sc_hd__mux2_1
X_28971_ _34793_/Q _24329_/X _28975_/S VGND VGND VPWR VPWR _28972_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_289_CLK clkbuf_6_57__f_CLK/X VGND VGND VPWR VPWR _36095_/CLK sky130_fd_sc_hd__clkbuf_16
X_23045_ _23044_/X _32067_/Q _23063_/S VGND VGND VPWR VPWR _23046_/A sky130_fd_sc_hd__mux2_1
X_27922_ _27922_/A VGND VGND VPWR VPWR _34295_/D sky130_fd_sc_hd__clkbuf_1
X_20257_ _20257_/A VGND VGND VPWR VPWR _20257_/X sky130_fd_sc_hd__buf_4
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27853_ _34263_/Q _24273_/X _27853_/S VGND VGND VPWR VPWR _27854_/A sky130_fd_sc_hd__mux2_1
XTAP_5225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20188_ _35585_/Q _35521_/Q _35457_/Q _35393_/Q _19903_/X _19904_/X VGND VGND VPWR
+ VPWR _20188_/X sky130_fd_sc_hd__mux4_1
XTAP_5236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26804_ _26804_/A VGND VGND VPWR VPWR _33797_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27784_ _34230_/Q _24369_/X _27802_/S VGND VGND VPWR VPWR _27785_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24996_ _24995_/X _32975_/Q _25020_/S VGND VGND VPWR VPWR _24997_/A sky130_fd_sc_hd__mux2_1
XTAP_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29523_ _35023_/Q _29055_/X _29539_/S VGND VGND VPWR VPWR _29524_/A sky130_fd_sc_hd__mux2_1
XTAP_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26735_ _26735_/A VGND VGND VPWR VPWR _33764_/D sky130_fd_sc_hd__clkbuf_1
X_23947_ _23947_/A VGND VGND VPWR VPWR _32513_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_801 _22889_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_461_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _35943_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29454_ _29454_/A VGND VGND VPWR VPWR _34990_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_812 _22914_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26666_ _26666_/A VGND VGND VPWR VPWR _33732_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_823 _23099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23878_ _22938_/X _32481_/Q _23878_/S VGND VGND VPWR VPWR _23879_/A sky130_fd_sc_hd__mux2_1
XTAP_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_834 _23346_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_845 _23696_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28405_ _28405_/A VGND VGND VPWR VPWR _34524_/D sky130_fd_sc_hd__clkbuf_1
X_22829_ _35852_/Q _32232_/Q _35724_/Q _35660_/Q _20589_/X _20591_/X VGND VGND VPWR
+ VPWR _22829_/X sky130_fd_sc_hd__mux4_1
X_25617_ _25617_/A VGND VGND VPWR VPWR _33236_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_856 _24342_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_867 _24428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29385_ _29517_/S VGND VGND VPWR VPWR _29404_/S sky130_fd_sc_hd__buf_4
X_26597_ _26597_/A VGND VGND VPWR VPWR _33699_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_878 _25041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_213_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _35080_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_889 _25458_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_241_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28336_ _34492_/Q _24388_/X _28342_/S VGND VGND VPWR VPWR _28337_/A sky130_fd_sc_hd__mux2_1
X_16350_ _17762_/A VGND VGND VPWR VPWR _16350_/X sky130_fd_sc_hd__buf_4
XFILLER_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25548_ _25548_/A VGND VGND VPWR VPWR _33205_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16281_ _16014_/X _16279_/X _16280_/X _16023_/X VGND VGND VPWR VPWR _16281_/X sky130_fd_sc_hd__a22o_1
XFILLER_73_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25479_ _25479_/A VGND VGND VPWR VPWR _33172_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28267_ _34459_/Q _24286_/X _28279_/S VGND VGND VPWR VPWR _28268_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18020_ _35781_/Q _35141_/Q _34501_/Q _33861_/Q _17846_/X _17847_/X VGND VGND VPWR
+ VPWR _18020_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27218_ _26912_/X _33963_/Q _27218_/S VGND VGND VPWR VPWR _27219_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28198_ _28198_/A VGND VGND VPWR VPWR _34426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27149_ _27149_/A VGND VGND VPWR VPWR _33930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30160_ _30160_/A VGND VGND VPWR VPWR _35325_/D sky130_fd_sc_hd__clkbuf_1
X_19971_ _35579_/Q _35515_/Q _35451_/Q _35387_/Q _19903_/X _19904_/X VGND VGND VPWR
+ VPWR _19971_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_1066 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18922_ _18918_/X _18921_/X _18755_/X VGND VGND VPWR VPWR _18923_/D sky130_fd_sc_hd__o21ba_1
X_30091_ _30091_/A VGND VGND VPWR VPWR _35292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1200 _23077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1211 _23319_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1222 _24295_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1233 _24425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18853_ _34523_/Q _32411_/Q _34395_/Q _34331_/Q _18819_/X _18820_/X VGND VGND VPWR
+ VPWR _18853_/X sky130_fd_sc_hd__mux4_1
XTAP_6460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1244 _26142_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1255 _26953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1266 _29652_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17804_ _33279_/Q _36159_/Q _33151_/Q _33087_/Q _17764_/X _17765_/X VGND VGND VPWR
+ VPWR _17804_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1277 _17903_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33850_ _35771_/CLK _33850_/D VGND VGND VPWR VPWR _33850_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1288 _17846_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18784_ _35033_/Q _34969_/Q _34905_/Q _34841_/Q _18750_/X _18751_/X VGND VGND VPWR
+ VPWR _18784_/X sky130_fd_sc_hd__mux4_1
XTAP_5770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15996_ _17769_/A VGND VGND VPWR VPWR _17860_/A sky130_fd_sc_hd__buf_12
XANTENNA_1299 _17157_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32801_ _35481_/CLK _32801_/D VGND VGND VPWR VPWR _32801_/Q sky130_fd_sc_hd__dfxtp_1
X_17735_ _33021_/Q _32957_/Q _32893_/Q _32829_/Q _17695_/X _17696_/X VGND VGND VPWR
+ VPWR _17735_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33781_ _34292_/CLK _33781_/D VGND VGND VPWR VPWR _33781_/Q sky130_fd_sc_hd__dfxtp_1
X_30993_ _35720_/Q _29231_/X _30995_/S VGND VGND VPWR VPWR _30994_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_1315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35520_ _35585_/CLK _35520_/D VGND VGND VPWR VPWR _35520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_452_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _35042_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32732_ _36127_/CLK _32732_/D VGND VGND VPWR VPWR _32732_/Q sky130_fd_sc_hd__dfxtp_1
X_17666_ _17795_/A VGND VGND VPWR VPWR _17666_/X sky130_fd_sc_hd__buf_6
XFILLER_39_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19405_ _35755_/Q _35115_/Q _34475_/Q _33835_/Q _19087_/X _19088_/X VGND VGND VPWR
+ VPWR _19405_/X sky130_fd_sc_hd__mux4_1
XFILLER_211_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35451_ _35515_/CLK _35451_/D VGND VGND VPWR VPWR _35451_/Q sky130_fd_sc_hd__dfxtp_1
X_16617_ _35293_/Q _35229_/Q _35165_/Q _32285_/Q _16300_/X _16301_/X VGND VGND VPWR
+ VPWR _16617_/X sky130_fd_sc_hd__mux4_1
X_32663_ _36116_/CLK _32663_/D VGND VGND VPWR VPWR _32663_/Q sky130_fd_sc_hd__dfxtp_1
X_17597_ _33017_/Q _32953_/Q _32889_/Q _32825_/Q _17342_/X _17343_/X VGND VGND VPWR
+ VPWR _17597_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_204_CLK clkbuf_6_52__f_CLK/X VGND VGND VPWR VPWR _35973_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_189_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34402_ _35932_/CLK _34402_/D VGND VGND VPWR VPWR _34402_/Q sky130_fd_sc_hd__dfxtp_1
X_19336_ _33193_/Q _32553_/Q _35945_/Q _35881_/Q _19021_/X _19022_/X VGND VGND VPWR
+ VPWR _19336_/X sky130_fd_sc_hd__mux4_1
X_31614_ _36014_/Q input26/X _31628_/S VGND VGND VPWR VPWR _31615_/A sky130_fd_sc_hd__mux2_1
X_16548_ _16293_/X _16546_/X _16547_/X _16296_/X VGND VGND VPWR VPWR _16548_/X sky130_fd_sc_hd__a22o_1
X_35382_ _35638_/CLK _35382_/D VGND VGND VPWR VPWR _35382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32594_ _36050_/CLK _32594_/D VGND VGND VPWR VPWR _32594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34333_ _35036_/CLK _34333_/D VGND VGND VPWR VPWR _34333_/Q sky130_fd_sc_hd__dfxtp_1
X_31545_ _31545_/A _31680_/B VGND VGND VPWR VPWR _31678_/S sky130_fd_sc_hd__nor2_8
X_19267_ _18946_/X _19265_/X _19266_/X _18949_/X VGND VGND VPWR VPWR _19267_/X sky130_fd_sc_hd__a22o_1
X_16479_ _16475_/X _16478_/X _16441_/X VGND VGND VPWR VPWR _16487_/C sky130_fd_sc_hd__o21ba_1
XFILLER_223_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18218_ _33548_/Q _33484_/Q _33420_/Q _33356_/Q _16033_/X _16035_/X VGND VGND VPWR
+ VPWR _18218_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34264_ _34265_/CLK _34264_/D VGND VGND VPWR VPWR _34264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19198_ _20257_/A VGND VGND VPWR VPWR _19198_/X sky130_fd_sc_hd__buf_4
X_31476_ _31476_/A VGND VGND VPWR VPWR _35948_/D sky130_fd_sc_hd__clkbuf_1
X_36003_ _36003_/CLK _36003_/D VGND VGND VPWR VPWR _36003_/Q sky130_fd_sc_hd__dfxtp_1
X_33215_ _36032_/CLK _33215_/D VGND VGND VPWR VPWR _33215_/Q sky130_fd_sc_hd__dfxtp_1
X_18149_ _34569_/Q _32457_/Q _34441_/Q _34377_/Q _17931_/X _17932_/X VGND VGND VPWR
+ VPWR _18149_/X sky130_fd_sc_hd__mux4_1
X_30427_ _30427_/A VGND VGND VPWR VPWR _35451_/D sky130_fd_sc_hd__clkbuf_1
X_34195_ _34259_/CLK _34195_/D VGND VGND VPWR VPWR _34195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33146_ _36090_/CLK _33146_/D VGND VGND VPWR VPWR _33146_/Q sky130_fd_sc_hd__dfxtp_1
X_21160_ _34268_/Q _34204_/Q _34140_/Q _34076_/Q _20983_/X _20984_/X VGND VGND VPWR
+ VPWR _21160_/X sky130_fd_sc_hd__mux4_1
X_30358_ _30358_/A VGND VGND VPWR VPWR _35418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20111_ _35775_/Q _35135_/Q _34495_/Q _33855_/Q _19793_/X _19794_/X VGND VGND VPWR
+ VPWR _20111_/X sky130_fd_sc_hd__mux4_1
XFILLER_217_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21091_ _22503_/A VGND VGND VPWR VPWR _21091_/X sky130_fd_sc_hd__buf_4
X_33077_ _34229_/CLK _33077_/D VGND VGND VPWR VPWR _33077_/Q sky130_fd_sc_hd__dfxtp_1
X_30289_ _30289_/A VGND VGND VPWR VPWR _35386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20042_ _33213_/Q _32573_/Q _35965_/Q _35901_/Q _19727_/X _19728_/X VGND VGND VPWR
+ VPWR _20042_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32028_ _32860_/CLK _32028_/D VGND VGND VPWR VPWR _32028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24850_ _23071_/X _32908_/Q _24852_/S VGND VGND VPWR VPWR _24851_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23801_ _23025_/X _32445_/Q _23805_/S VGND VGND VPWR VPWR _23802_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24781_ _22969_/X _32875_/Q _24781_/S VGND VGND VPWR VPWR _24782_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33979_ _34171_/CLK _33979_/D VGND VGND VPWR VPWR _33979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21993_ _35315_/Q _35251_/Q _35187_/Q _32307_/Q _21959_/X _21960_/X VGND VGND VPWR
+ VPWR _21993_/X sky130_fd_sc_hd__mux4_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_443_CLK clkbuf_6_14__f_CLK/X VGND VGND VPWR VPWR _36069_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_215_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26520_ _26547_/S VGND VGND VPWR VPWR _26539_/S sky130_fd_sc_hd__buf_6
XFILLER_187_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_108 _32129_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23732_ _22923_/X _32412_/Q _23742_/S VGND VGND VPWR VPWR _23733_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20944_ _20736_/X _20942_/X _20943_/X _20741_/X VGND VGND VPWR VPWR _20944_/X sky130_fd_sc_hd__a22o_1
X_35718_ _35849_/CLK _35718_/D VGND VGND VPWR VPWR _35718_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_119 _32131_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23663_ _32381_/Q _23294_/X _23667_/S VGND VGND VPWR VPWR _23664_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26451_ _25044_/X _33631_/Q _26455_/S VGND VGND VPWR VPWR _26452_/A sky130_fd_sc_hd__mux2_1
X_20875_ _33492_/Q _33428_/Q _33364_/Q _33300_/Q _20598_/X _20599_/X VGND VGND VPWR
+ VPWR _20875_/X sky130_fd_sc_hd__mux4_1
X_35649_ _35715_/CLK _35649_/D VGND VGND VPWR VPWR _35649_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22614_ _22361_/X _22612_/X _22613_/X _22367_/X VGND VGND VPWR VPWR _22614_/X sky130_fd_sc_hd__a22o_1
X_25402_ _25103_/X _33138_/Q _25408_/S VGND VGND VPWR VPWR _25403_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26382_ _26382_/A VGND VGND VPWR VPWR _33598_/D sky130_fd_sc_hd__clkbuf_1
X_29170_ _34868_/Q _29169_/X _29173_/S VGND VGND VPWR VPWR _29171_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23594_ _32348_/Q _23130_/X _23604_/S VGND VGND VPWR VPWR _23595_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25333_ _25001_/X _33105_/Q _25345_/S VGND VGND VPWR VPWR _25334_/A sky130_fd_sc_hd__mux2_1
X_28121_ _26847_/X _34390_/Q _28123_/S VGND VGND VPWR VPWR _28122_/A sky130_fd_sc_hd__mux2_1
X_22545_ _22541_/X _22544_/X _22434_/X VGND VGND VPWR VPWR _22569_/A sky130_fd_sc_hd__o21ba_1
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25264_ _25100_/X _33073_/Q _25272_/S VGND VGND VPWR VPWR _25265_/A sky130_fd_sc_hd__mux2_1
X_28052_ _28052_/A VGND VGND VPWR VPWR _34357_/D sky130_fd_sc_hd__clkbuf_1
X_22476_ _22155_/X _22474_/X _22475_/X _22158_/X VGND VGND VPWR VPWR _22476_/X sky130_fd_sc_hd__a22o_1
XFILLER_6_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27003_ _27002_/X _33864_/Q _27006_/S VGND VGND VPWR VPWR _27004_/A sky130_fd_sc_hd__mux2_1
X_24215_ _24242_/S VGND VGND VPWR VPWR _24234_/S sky130_fd_sc_hd__buf_6
XFILLER_154_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21427_ _35747_/Q _35107_/Q _34467_/Q _33827_/Q _21387_/X _21388_/X VGND VGND VPWR
+ VPWR _21427_/X sky130_fd_sc_hd__mux4_1
X_25195_ _24998_/X _33040_/Q _25209_/S VGND VGND VPWR VPWR _25196_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24146_ _22932_/X _32607_/Q _24150_/S VGND VGND VPWR VPWR _24147_/A sky130_fd_sc_hd__mux2_1
X_21358_ _34785_/Q _34721_/Q _34657_/Q _34593_/Q _21182_/X _21183_/X VGND VGND VPWR
+ VPWR _21358_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20309_ _34053_/Q _33989_/Q _33925_/Q _32261_/Q _20026_/X _20027_/X VGND VGND VPWR
+ VPWR _20309_/X sky130_fd_sc_hd__mux4_1
X_24077_ _23031_/X _32575_/Q _24077_/S VGND VGND VPWR VPWR _24078_/A sky130_fd_sc_hd__mux2_1
X_28954_ _34785_/Q _24304_/X _28954_/S VGND VGND VPWR VPWR _28955_/A sky130_fd_sc_hd__mux2_1
X_21289_ _34527_/Q _32415_/Q _34399_/Q _34335_/Q _21119_/X _21120_/X VGND VGND VPWR
+ VPWR _21289_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23028_ input43/X VGND VGND VPWR VPWR _23028_/X sky130_fd_sc_hd__clkbuf_4
X_27905_ _27905_/A VGND VGND VPWR VPWR _34287_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28885_ _26977_/X _34752_/Q _28903_/S VGND VGND VPWR VPWR _28886_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27836_ _27836_/A VGND VGND VPWR VPWR _34254_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27767_ _34222_/Q _24345_/X _27781_/S VGND VGND VPWR VPWR _27768_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24979_ _23062_/X _32969_/Q _24979_/S VGND VGND VPWR VPWR _24980_/A sky130_fd_sc_hd__mux2_1
XTAP_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_434_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _34870_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_73_930 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29506_ _29506_/A VGND VGND VPWR VPWR _35015_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17520_ _17195_/X _17518_/X _17519_/X _17200_/X VGND VGND VPWR VPWR _17520_/X sky130_fd_sc_hd__a22o_1
XTAP_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26718_ _26718_/A VGND VGND VPWR VPWR _33756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27698_ _27833_/A _29924_/A VGND VGND VPWR VPWR _27831_/S sky130_fd_sc_hd__nor2_8
XTAP_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_620 _18571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_631 _18891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29437_ _29437_/A VGND VGND VPWR VPWR _34982_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_642 _19356_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _33269_/Q _36149_/Q _33141_/Q _33077_/Q _17411_/X _17412_/X VGND VGND VPWR
+ VPWR _17451_/X sky130_fd_sc_hd__mux4_1
X_26649_ _26649_/A VGND VGND VPWR VPWR _33724_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_653 _20238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_664 _22395_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_675 _22511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16402_ _33175_/Q _32535_/Q _35927_/Q _35863_/Q _16368_/X _16369_/X VGND VGND VPWR
+ VPWR _16402_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_686 _22501_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29368_ _23322_/X _34950_/Q _29374_/S VGND VGND VPWR VPWR _29369_/A sky130_fd_sc_hd__mux2_1
XANTENNA_697 _22458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17382_ _33011_/Q _32947_/Q _32883_/Q _32819_/Q _17342_/X _17343_/X VGND VGND VPWR
+ VPWR _17382_/X sky130_fd_sc_hd__mux4_1
XFILLER_186_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19121_ _19002_/X _19119_/X _19120_/X _19008_/X VGND VGND VPWR VPWR _19121_/X sky130_fd_sc_hd__a22o_1
X_16333_ _34773_/Q _34709_/Q _34645_/Q _34581_/Q _16229_/X _16230_/X VGND VGND VPWR
+ VPWR _16333_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28319_ _34484_/Q _24363_/X _28321_/S VGND VGND VPWR VPWR _28320_/A sky130_fd_sc_hd__mux2_1
X_29299_ _23199_/X _34917_/Q _29311_/S VGND VGND VPWR VPWR _29300_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31330_ _31330_/A VGND VGND VPWR VPWR _35879_/D sky130_fd_sc_hd__clkbuf_1
X_19052_ _35745_/Q _35105_/Q _34465_/Q _33825_/Q _18734_/X _18735_/X VGND VGND VPWR
+ VPWR _19052_/X sky130_fd_sc_hd__mux4_1
X_16264_ _35283_/Q _35219_/Q _35155_/Q _32275_/Q _16079_/X _16081_/X VGND VGND VPWR
+ VPWR _16264_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18003_ _18003_/A _18003_/B _18003_/C _18003_/D VGND VGND VPWR VPWR _18004_/A sky130_fd_sc_hd__or4_4
XFILLER_199_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31261_ _35847_/Q input53/X _31265_/S VGND VGND VPWR VPWR _31262_/A sky130_fd_sc_hd__mux2_1
X_16195_ _16056_/X _16193_/X _16194_/X _16068_/X VGND VGND VPWR VPWR _16195_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33000_ _36009_/CLK _33000_/D VGND VGND VPWR VPWR _33000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30212_ _35350_/Q _29076_/X _30214_/S VGND VGND VPWR VPWR _30213_/A sky130_fd_sc_hd__mux2_1
X_31192_ _35814_/Q input17/X _31202_/S VGND VGND VPWR VPWR _31193_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19954_ _19848_/X _19952_/X _19953_/X _19853_/X VGND VGND VPWR VPWR _19954_/X sky130_fd_sc_hd__a22o_1
X_30143_ _30143_/A VGND VGND VPWR VPWR _35317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18905_ _18657_/X _18903_/X _18904_/X _18661_/X VGND VGND VPWR VPWR _18905_/X sky130_fd_sc_hd__a22o_1
X_34951_ _35079_/CLK _34951_/D VGND VGND VPWR VPWR _34951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30074_ _30074_/A VGND VGND VPWR VPWR _35284_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_1030 _17865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19885_ _19885_/A VGND VGND VPWR VPWR _32120_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA_1041 _17154_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1052 _16135_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18836_ _18649_/X _18834_/X _18835_/X _18655_/X VGND VGND VPWR VPWR _18836_/X sky130_fd_sc_hd__a22o_1
XANTENNA_1063 _16765_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33902_ _34032_/CLK _33902_/D VGND VGND VPWR VPWR _33902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34882_ _34947_/CLK _34882_/D VGND VGND VPWR VPWR _34882_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1074 _17164_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1085 _17232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1096 _17264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33833_ _34859_/CLK _33833_/D VGND VGND VPWR VPWR _33833_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_43__f_CLK clkbuf_5_21_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_43__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_18767_ _33241_/Q _36121_/Q _33113_/Q _33049_/Q _18652_/X _18653_/X VGND VGND VPWR
+ VPWR _18767_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15979_ _16057_/A VGND VGND VPWR VPWR _17902_/A sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_425_CLK clkbuf_6_36__f_CLK/X VGND VGND VPWR VPWR _36075_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_209_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17718_ _17507_/X _17716_/X _17717_/X _17512_/X VGND VGND VPWR VPWR _17718_/X sky130_fd_sc_hd__a22o_1
XFILLER_236_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33764_ _34277_/CLK _33764_/D VGND VGND VPWR VPWR _33764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30976_ _31003_/S VGND VGND VPWR VPWR _30995_/S sky130_fd_sc_hd__buf_4
X_18698_ _35799_/Q _32174_/Q _35671_/Q _35607_/Q _18554_/X _18555_/X VGND VGND VPWR
+ VPWR _18698_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32715_ _36171_/CLK _32715_/D VGND VGND VPWR VPWR _32715_/Q sky130_fd_sc_hd__dfxtp_1
X_35503_ _35951_/CLK _35503_/D VGND VGND VPWR VPWR _35503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17649_ _17645_/X _17648_/X _17514_/X VGND VGND VPWR VPWR _17650_/D sky130_fd_sc_hd__o21ba_1
XFILLER_36_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33695_ _34016_/CLK _33695_/D VGND VGND VPWR VPWR _33695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35434_ _35562_/CLK _35434_/D VGND VGND VPWR VPWR _35434_/Q sky130_fd_sc_hd__dfxtp_1
X_20660_ _22447_/A VGND VGND VPWR VPWR _20660_/X sky130_fd_sc_hd__buf_6
X_32646_ _36103_/CLK _32646_/D VGND VGND VPWR VPWR _32646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19319_ _33513_/Q _33449_/Q _33385_/Q _33321_/Q _19070_/X _19071_/X VGND VGND VPWR
+ VPWR _19319_/X sky130_fd_sc_hd__mux4_1
X_35365_ _35749_/CLK _35365_/D VGND VGND VPWR VPWR _35365_/Q sky130_fd_sc_hd__dfxtp_1
X_20591_ _22396_/A VGND VGND VPWR VPWR _20591_/X sky130_fd_sc_hd__buf_4
X_32577_ _35906_/CLK _32577_/D VGND VGND VPWR VPWR _32577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34316_ _34316_/CLK _34316_/D VGND VGND VPWR VPWR _34316_/Q sky130_fd_sc_hd__dfxtp_1
X_22330_ _22324_/X _22329_/X _22081_/X VGND VGND VPWR VPWR _22352_/A sky130_fd_sc_hd__o21ba_1
XFILLER_109_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31528_ _31528_/A VGND VGND VPWR VPWR _35973_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35296_ _35296_/CLK _35296_/D VGND VGND VPWR VPWR _35296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34247_ _34819_/CLK _34247_/D VGND VGND VPWR VPWR _34247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22261_ _22008_/X _22259_/X _22260_/X _22014_/X VGND VGND VPWR VPWR _22261_/X sky130_fd_sc_hd__a22o_1
X_31459_ _31459_/A VGND VGND VPWR VPWR _35940_/D sky130_fd_sc_hd__clkbuf_1
X_24000_ _22917_/X _32538_/Q _24014_/S VGND VGND VPWR VPWR _24001_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21212_ _35549_/Q _35485_/Q _35421_/Q _35357_/Q _21144_/X _21145_/X VGND VGND VPWR
+ VPWR _21212_/X sky130_fd_sc_hd__mux4_1
X_34178_ _34243_/CLK _34178_/D VGND VGND VPWR VPWR _34178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22192_ _22188_/X _22191_/X _22081_/X VGND VGND VPWR VPWR _22216_/A sky130_fd_sc_hd__o21ba_1
XFILLER_183_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21143_ _20888_/X _21141_/X _21142_/X _20891_/X VGND VGND VPWR VPWR _21143_/X sky130_fd_sc_hd__a22o_1
X_33129_ _33255_/CLK _33129_/D VGND VGND VPWR VPWR _33129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21074_ _35737_/Q _35097_/Q _34457_/Q _33817_/Q _21034_/X _21035_/X VGND VGND VPWR
+ VPWR _21074_/X sky130_fd_sc_hd__mux4_1
X_25951_ _25103_/X _33394_/Q _25957_/S VGND VGND VPWR VPWR _25952_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20025_ _33533_/Q _33469_/Q _33405_/Q _33341_/Q _19776_/X _19777_/X VGND VGND VPWR
+ VPWR _20025_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24902_ _22948_/X _32932_/Q _24916_/S VGND VGND VPWR VPWR _24903_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28670_ _26860_/X _34650_/Q _28684_/S VGND VGND VPWR VPWR _28671_/A sky130_fd_sc_hd__mux2_1
X_25882_ _25001_/X _33361_/Q _25894_/S VGND VGND VPWR VPWR _25883_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27621_ _34153_/Q _24329_/X _27625_/S VGND VGND VPWR VPWR _27622_/A sky130_fd_sc_hd__mux2_1
X_24833_ _24833_/A VGND VGND VPWR VPWR _32899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_416_CLK clkbuf_6_35__f_CLK/X VGND VGND VPWR VPWR _34797_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_132_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27552_ _27552_/A VGND VGND VPWR VPWR _34121_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24764_ _24764_/A VGND VGND VPWR VPWR _32866_/D sky130_fd_sc_hd__clkbuf_1
X_21976_ _21802_/X _21972_/X _21975_/X _21805_/X VGND VGND VPWR VPWR _21976_/X sky130_fd_sc_hd__a22o_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26503_ _26503_/A VGND VGND VPWR VPWR _33655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20927_ _35733_/Q _35093_/Q _34453_/Q _33813_/Q _20649_/X _20651_/X VGND VGND VPWR
+ VPWR _20927_/X sky130_fd_sc_hd__mux4_1
X_23715_ _22898_/X _32404_/Q _23721_/S VGND VGND VPWR VPWR _23716_/A sky130_fd_sc_hd__mux2_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24695_ _23044_/X _32835_/Q _24707_/S VGND VGND VPWR VPWR _24696_/A sky130_fd_sc_hd__mux2_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_7_0_CLK/A sky130_fd_sc_hd__clkbuf_8
X_27483_ _27483_/A VGND VGND VPWR VPWR _34088_/D sky130_fd_sc_hd__clkbuf_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29222_ input51/X VGND VGND VPWR VPWR _29222_/X sky130_fd_sc_hd__clkbuf_4
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26434_ _25019_/X _33623_/Q _26434_/S VGND VGND VPWR VPWR _26435_/A sky130_fd_sc_hd__mux2_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20858_ _20644_/X _20856_/X _20857_/X _20654_/X VGND VGND VPWR VPWR _20858_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23646_ _32373_/Q _23267_/X _23646_/S VGND VGND VPWR VPWR _23647_/A sky130_fd_sc_hd__mux2_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29153_ _29153_/A VGND VGND VPWR VPWR _34862_/D sky130_fd_sc_hd__clkbuf_1
X_23577_ _32340_/Q _23105_/X _23583_/S VGND VGND VPWR VPWR _23578_/A sky130_fd_sc_hd__mux2_1
X_26365_ _25115_/X _33590_/Q _26383_/S VGND VGND VPWR VPWR _26366_/A sky130_fd_sc_hd__mux2_1
X_20789_ _35729_/Q _35089_/Q _34449_/Q _33809_/Q _20649_/X _20651_/X VGND VGND VPWR
+ VPWR _20789_/X sky130_fd_sc_hd__mux4_1
XFILLER_210_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28104_ _28236_/S VGND VGND VPWR VPWR _28123_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_167_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22528_ _34818_/Q _34754_/Q _34690_/Q _34626_/Q _22241_/X _22242_/X VGND VGND VPWR
+ VPWR _22528_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25316_ _25177_/X _33098_/Q _25322_/S VGND VGND VPWR VPWR _25317_/A sky130_fd_sc_hd__mux2_1
X_26296_ _26296_/A VGND VGND VPWR VPWR _33557_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29084_ _34840_/Q _29082_/X _29111_/S VGND VGND VPWR VPWR _29085_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28035_ _26919_/X _34349_/Q _28051_/S VGND VGND VPWR VPWR _28036_/A sky130_fd_sc_hd__mux2_1
X_22459_ _22455_/X _22456_/X _22457_/X _22458_/X VGND VGND VPWR VPWR _22459_/X sky130_fd_sc_hd__a22o_1
X_25247_ _25075_/X _33065_/Q _25251_/S VGND VGND VPWR VPWR _25248_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25178_ _25177_/X _33034_/Q _25187_/S VGND VGND VPWR VPWR _25179_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24129_ _22907_/X _32599_/Q _24129_/S VGND VGND VPWR VPWR _24130_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29986_ _35243_/Q _29141_/X _29986_/S VGND VGND VPWR VPWR _29987_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28937_ _28937_/A VGND VGND VPWR VPWR _34776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16951_ _16849_/X _16949_/X _16950_/X _16852_/X VGND VGND VPWR VPWR _16951_/X sky130_fd_sc_hd__a22o_1
XFILLER_1_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_836 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19670_ _34291_/Q _34227_/Q _34163_/Q _34099_/Q _19389_/X _19390_/X VGND VGND VPWR
+ VPWR _19670_/X sky130_fd_sc_hd__mux4_1
X_16882_ _16842_/X _16880_/X _16881_/X _16847_/X VGND VGND VPWR VPWR _16882_/X sky130_fd_sc_hd__a22o_1
X_28868_ _26953_/X _34744_/Q _28882_/S VGND VGND VPWR VPWR _28869_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18621_ _18314_/X _18619_/X _18620_/X _18323_/X VGND VGND VPWR VPWR _18621_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27819_ _34247_/Q _24422_/X _27823_/S VGND VGND VPWR VPWR _27820_/A sky130_fd_sc_hd__mux2_1
XTAP_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28799_ _28799_/A VGND VGND VPWR VPWR _34711_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_407_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _35307_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18552_ _18326_/X _18550_/X _18551_/X _18337_/X VGND VGND VPWR VPWR _18552_/X sky130_fd_sc_hd__a22o_1
XTAP_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30830_ _30830_/A VGND VGND VPWR VPWR _35642_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ _34806_/Q _34742_/Q _34678_/Q _34614_/Q _17288_/X _17289_/X VGND VGND VPWR
+ VPWR _17503_/X sky130_fd_sc_hd__mux4_1
XTAP_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18483_ _18314_/X _18481_/X _18482_/X _18323_/X VGND VGND VPWR VPWR _18483_/X sky130_fd_sc_hd__a22o_1
XTAP_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30761_ _30761_/A VGND VGND VPWR VPWR _35609_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_450 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32500_ _33013_/CLK _32500_/D VGND VGND VPWR VPWR _32500_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_461 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17434_ _17149_/X _17432_/X _17433_/X _17152_/X VGND VGND VPWR VPWR _17434_/X sky130_fd_sc_hd__a22o_1
XANTENNA_472 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33480_ _33795_/CLK _33480_/D VGND VGND VPWR VPWR _33480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_483 _31994_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30692_ _35577_/Q _29185_/X _30704_/S VGND VGND VPWR VPWR _30693_/A sky130_fd_sc_hd__mux2_1
XANTENNA_494 _31995_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_221_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32431_ _35758_/CLK _32431_/D VGND VGND VPWR VPWR _32431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_19 _32115_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17365_ _17154_/X _17363_/X _17364_/X _17159_/X VGND VGND VPWR VPWR _17365_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19104_ _19457_/A VGND VGND VPWR VPWR _19104_/X sky130_fd_sc_hd__buf_4
X_16316_ _34005_/Q _33941_/Q _33877_/Q _32149_/Q _16314_/X _16315_/X VGND VGND VPWR
+ VPWR _16316_/X sky130_fd_sc_hd__mux4_1
X_35150_ _36216_/CLK _35150_/D VGND VGND VPWR VPWR _35150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32362_ _34739_/CLK _32362_/D VGND VGND VPWR VPWR _32362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17296_ _17292_/X _17295_/X _17161_/X VGND VGND VPWR VPWR _17297_/D sky130_fd_sc_hd__o21ba_1
XFILLER_174_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34101_ _34229_/CLK _34101_/D VGND VGND VPWR VPWR _34101_/Q sky130_fd_sc_hd__dfxtp_1
X_19035_ _33761_/Q _33697_/Q _33633_/Q _33569_/Q _18790_/X _18791_/X VGND VGND VPWR
+ VPWR _19035_/X sky130_fd_sc_hd__mux4_1
X_31313_ _31313_/A VGND VGND VPWR VPWR _35871_/D sky130_fd_sc_hd__clkbuf_1
X_35081_ _35781_/CLK _35081_/D VGND VGND VPWR VPWR _35081_/Q sky130_fd_sc_hd__dfxtp_1
X_16247_ _32723_/Q _32659_/Q _32595_/Q _36051_/Q _16213_/X _17713_/A VGND VGND VPWR
+ VPWR _16247_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32293_ _36005_/CLK _32293_/D VGND VGND VPWR VPWR _32293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34032_ _34032_/CLK _34032_/D VGND VGND VPWR VPWR _34032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31244_ _35839_/Q input44/X _31244_/S VGND VGND VPWR VPWR _31245_/A sky130_fd_sc_hd__mux2_1
Xoutput104 _31972_/Q VGND VGND VPWR VPWR D1[22] sky130_fd_sc_hd__buf_2
X_16178_ _34001_/Q _33937_/Q _33873_/Q _32145_/Q _16108_/X _16109_/X VGND VGND VPWR
+ VPWR _16178_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput115 _31982_/Q VGND VGND VPWR VPWR D1[32] sky130_fd_sc_hd__buf_2
XFILLER_47_1106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput126 _31992_/Q VGND VGND VPWR VPWR D1[42] sky130_fd_sc_hd__buf_2
Xoutput137 _32002_/Q VGND VGND VPWR VPWR D1[52] sky130_fd_sc_hd__buf_2
Xoutput148 _32012_/Q VGND VGND VPWR VPWR D1[62] sky130_fd_sc_hd__buf_2
Xoutput159 _36188_/Q VGND VGND VPWR VPWR D2[14] sky130_fd_sc_hd__buf_2
X_31175_ _35806_/Q input8/X _31181_/S VGND VGND VPWR VPWR _31176_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30126_ _35309_/Q _29148_/X _30142_/S VGND VGND VPWR VPWR _30127_/A sky130_fd_sc_hd__mux2_1
X_19937_ _35578_/Q _35514_/Q _35450_/Q _35386_/Q _19903_/X _19904_/X VGND VGND VPWR
+ VPWR _19937_/X sky130_fd_sc_hd__mux4_2
X_35983_ _36041_/CLK _35983_/D VGND VGND VPWR VPWR _35983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30057_ _35277_/Q _29246_/X _30057_/S VGND VGND VPWR VPWR _30058_/A sky130_fd_sc_hd__mux2_1
X_34934_ _35257_/CLK _34934_/D VGND VGND VPWR VPWR _34934_/Q sky130_fd_sc_hd__dfxtp_1
X_19868_ _35832_/Q _32210_/Q _35704_/Q _35640_/Q _19613_/X _19614_/X VGND VGND VPWR
+ VPWR _19868_/X sky130_fd_sc_hd__mux4_1
XFILLER_112_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18819_ _20012_/A VGND VGND VPWR VPWR _18819_/X sky130_fd_sc_hd__buf_6
X_34865_ _34866_/CLK _34865_/D VGND VGND VPWR VPWR _34865_/Q sky130_fd_sc_hd__dfxtp_1
X_19799_ _19652_/X _19797_/X _19798_/X _19655_/X VGND VGND VPWR VPWR _19799_/X sky130_fd_sc_hd__a22o_1
X_21830_ _21824_/X _21829_/X _21761_/X VGND VGND VPWR VPWR _21831_/D sky130_fd_sc_hd__o21ba_1
XFILLER_209_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33816_ _35738_/CLK _33816_/D VGND VGND VPWR VPWR _33816_/Q sky130_fd_sc_hd__dfxtp_1
X_34796_ _34797_/CLK _34796_/D VGND VGND VPWR VPWR _34796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33747_ _34259_/CLK _33747_/D VGND VGND VPWR VPWR _33747_/Q sky130_fd_sc_hd__dfxtp_1
X_21761_ _22467_/A VGND VGND VPWR VPWR _21761_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_97_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30959_ _30959_/A VGND VGND VPWR VPWR _35703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20712_ _20706_/X _20711_/X _20611_/X VGND VGND VPWR VPWR _20734_/A sky130_fd_sc_hd__o21ba_1
X_23500_ _23500_/A VGND VGND VPWR VPWR _32304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24480_ _24480_/A VGND VGND VPWR VPWR _32734_/D sky130_fd_sc_hd__clkbuf_1
X_33678_ _35277_/CLK _33678_/D VGND VGND VPWR VPWR _33678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21692_ _21442_/X _21688_/X _21691_/X _21447_/X VGND VGND VPWR VPWR _21692_/X sky130_fd_sc_hd__a22o_1
XFILLER_197_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23431_ _23431_/A VGND VGND VPWR VPWR _32271_/D sky130_fd_sc_hd__clkbuf_1
X_20643_ _20624_/X _20638_/X _20640_/X _20642_/X VGND VGND VPWR VPWR _20702_/B sky130_fd_sc_hd__o211a_1
X_35417_ _35801_/CLK _35417_/D VGND VGND VPWR VPWR _35417_/Q sky130_fd_sc_hd__dfxtp_1
X_32629_ _36085_/CLK _32629_/D VGND VGND VPWR VPWR _32629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26150_ _24998_/X _33488_/Q _26164_/S VGND VGND VPWR VPWR _26151_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35348_ _35797_/CLK _35348_/D VGND VGND VPWR VPWR _35348_/Q sky130_fd_sc_hd__dfxtp_1
X_23362_ _23362_/A VGND VGND VPWR VPWR _32240_/D sky130_fd_sc_hd__clkbuf_1
X_20574_ _20574_/A VGND VGND VPWR VPWR _32141_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_164_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1014 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22313_ _22313_/A VGND VGND VPWR VPWR _22313_/X sky130_fd_sc_hd__buf_6
X_25101_ _25100_/X _33009_/Q _25113_/S VGND VGND VPWR VPWR _25102_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26081_ _26081_/A VGND VGND VPWR VPWR _33455_/D sky130_fd_sc_hd__clkbuf_1
X_35279_ _35279_/CLK _35279_/D VGND VGND VPWR VPWR _35279_/Q sky130_fd_sc_hd__dfxtp_1
X_23293_ _23293_/A VGND VGND VPWR VPWR _32215_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25032_ input5/X VGND VGND VPWR VPWR _25032_/X sky130_fd_sc_hd__buf_2
X_22244_ _35322_/Q _35258_/Q _35194_/Q _32314_/Q _21959_/X _21960_/X VGND VGND VPWR
+ VPWR _22244_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29840_ _29840_/A VGND VGND VPWR VPWR _35173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22175_ _34808_/Q _34744_/Q _34680_/Q _34616_/Q _21888_/X _21889_/X VGND VGND VPWR
+ VPWR _22175_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21126_ _21126_/A VGND VGND VPWR VPWR _36186_/D sky130_fd_sc_hd__clkbuf_1
X_29771_ _35141_/Q _29222_/X _29779_/S VGND VGND VPWR VPWR _29772_/A sky130_fd_sc_hd__mux2_1
X_26983_ _26983_/A VGND VGND VPWR VPWR _33857_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28722_ _26937_/X _34675_/Q _28726_/S VGND VGND VPWR VPWR _28723_/A sky130_fd_sc_hd__mux2_1
X_25934_ _25078_/X _33386_/Q _25936_/S VGND VGND VPWR VPWR _25935_/A sky130_fd_sc_hd__mux2_1
X_21057_ _21057_/A _21057_/B _21057_/C _21057_/D VGND VGND VPWR VPWR _21058_/A sky130_fd_sc_hd__or4_2
XFILLER_232_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20008_ _20165_/A VGND VGND VPWR VPWR _20008_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28653_ _26835_/X _34642_/Q _28663_/S VGND VGND VPWR VPWR _28654_/A sky130_fd_sc_hd__mux2_1
X_25865_ _25865_/A VGND VGND VPWR VPWR _33353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27604_ _34145_/Q _24304_/X _27604_/S VGND VGND VPWR VPWR _27605_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24816_ _24816_/A VGND VGND VPWR VPWR _32891_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_963 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28584_ _28584_/A VGND VGND VPWR VPWR _34609_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_1029 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25796_ _25796_/A VGND VGND VPWR VPWR _33320_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27535_ _26981_/X _34113_/Q _27551_/S VGND VGND VPWR VPWR _27536_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24747_ _24747_/A VGND VGND VPWR VPWR _32858_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21959_ _22312_/A VGND VGND VPWR VPWR _21959_/X sky130_fd_sc_hd__buf_6
XFILLER_203_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27466_ _27466_/A VGND VGND VPWR VPWR _34080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24678_ _23019_/X _32827_/Q _24686_/S VGND VGND VPWR VPWR _24679_/A sky130_fd_sc_hd__mux2_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29205_ _29205_/A VGND VGND VPWR VPWR _34879_/D sky130_fd_sc_hd__clkbuf_1
X_26417_ _26417_/A VGND VGND VPWR VPWR _33614_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23629_ _23629_/A VGND VGND VPWR VPWR _32364_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27397_ _27424_/S VGND VGND VPWR VPWR _27416_/S sky130_fd_sc_hd__buf_4
XFILLER_208_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29136_ _34857_/Q _29135_/X _29142_/S VGND VGND VPWR VPWR _29137_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17150_ _34796_/Q _34732_/Q _34668_/Q _34604_/Q _16935_/X _16936_/X VGND VGND VPWR
+ VPWR _17150_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26348_ _25091_/X _33582_/Q _26362_/S VGND VGND VPWR VPWR _26349_/A sky130_fd_sc_hd__mux2_1
Xinput17 DW[24] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__buf_4
X_16101_ _16085_/X _16098_/X _16100_/X VGND VGND VPWR VPWR _16102_/D sky130_fd_sc_hd__o21ba_1
XFILLER_168_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput28 DW[34] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__buf_4
Xinput39 DW[44] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__clkbuf_8
X_29067_ input56/X VGND VGND VPWR VPWR _29067_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_122_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17081_ _16796_/X _17079_/X _17080_/X _16799_/X VGND VGND VPWR VPWR _17081_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_6_7__f_CLK clkbuf_5_3_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_7__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_26279_ _30735_/B _26685_/B VGND VGND VPWR VPWR _26412_/S sky130_fd_sc_hd__nand2_8
XFILLER_155_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16032_ _16057_/A VGND VGND VPWR VPWR _17829_/A sky130_fd_sc_hd__buf_12
XFILLER_171_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28018_ _26894_/X _34341_/Q _28030_/S VGND VGND VPWR VPWR _28019_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17983_ _32516_/Q _32388_/Q _32068_/Q _36036_/Q _17982_/X _17770_/X VGND VGND VPWR
+ VPWR _17983_/X sky130_fd_sc_hd__mux4_1
X_29969_ _29969_/A VGND VGND VPWR VPWR _35234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19722_ _19715_/X _19721_/X _19436_/X _19437_/X VGND VGND VPWR VPWR _19739_/B sky130_fd_sc_hd__o211a_1
X_16934_ _16930_/X _16933_/X _16794_/X VGND VGND VPWR VPWR _16944_/C sky130_fd_sc_hd__o21ba_1
XFILLER_238_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32980_ _32983_/CLK _32980_/D VGND VGND VPWR VPWR _32980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31931_ _31931_/A VGND VGND VPWR VPWR _36164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19653_ _35570_/Q _35506_/Q _35442_/Q _35378_/Q _19550_/X _19551_/X VGND VGND VPWR
+ VPWR _19653_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16865_ _35556_/Q _35492_/Q _35428_/Q _35364_/Q _16544_/X _16545_/X VGND VGND VPWR
+ VPWR _16865_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18604_ _34516_/Q _32404_/Q _34388_/Q _34324_/Q _18466_/X _18467_/X VGND VGND VPWR
+ VPWR _18604_/X sky130_fd_sc_hd__mux4_1
X_34650_ _36201_/CLK _34650_/D VGND VGND VPWR VPWR _34650_/Q sky130_fd_sc_hd__dfxtp_1
X_19584_ _35568_/Q _35504_/Q _35440_/Q _35376_/Q _19550_/X _19551_/X VGND VGND VPWR
+ VPWR _19584_/X sky130_fd_sc_hd__mux4_1
X_31862_ _31862_/A VGND VGND VPWR VPWR _36131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_237_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16796_ _17149_/A VGND VGND VPWR VPWR _16796_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_168_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33601_ _33729_/CLK _33601_/D VGND VGND VPWR VPWR _33601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18535_ _35026_/Q _34962_/Q _34898_/Q _34834_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _18535_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30813_ _30813_/A VGND VGND VPWR VPWR _35634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34581_ _36189_/CLK _34581_/D VGND VGND VPWR VPWR _34581_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31793_ _36099_/Q input49/X _31805_/S VGND VGND VPWR VPWR _31794_/A sky130_fd_sc_hd__mux2_1
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33532_ _33723_/CLK _33532_/D VGND VGND VPWR VPWR _33532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30744_ _30744_/A VGND VGND VPWR VPWR _35601_/D sky130_fd_sc_hd__clkbuf_1
X_18466_ _20012_/A VGND VGND VPWR VPWR _18466_/X sky130_fd_sc_hd__buf_6
XFILLER_34_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_280 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_291 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17417_ _17770_/A VGND VGND VPWR VPWR _17417_/X sky130_fd_sc_hd__clkbuf_4
X_33463_ _34297_/CLK _33463_/D VGND VGND VPWR VPWR _33463_/Q sky130_fd_sc_hd__dfxtp_1
X_18397_ _19459_/A VGND VGND VPWR VPWR _18397_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_159_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30675_ _35569_/Q _29160_/X _30683_/S VGND VGND VPWR VPWR _30676_/A sky130_fd_sc_hd__mux2_1
X_35202_ _35330_/CLK _35202_/D VGND VGND VPWR VPWR _35202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32414_ _35294_/CLK _32414_/D VGND VGND VPWR VPWR _32414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36182_ _36202_/CLK _36182_/D VGND VGND VPWR VPWR _36182_/Q sky130_fd_sc_hd__dfxtp_1
X_17348_ _35826_/Q _32203_/Q _35698_/Q _35634_/Q _17313_/X _17314_/X VGND VGND VPWR
+ VPWR _17348_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33394_ _33775_/CLK _33394_/D VGND VGND VPWR VPWR _33394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35133_ _35711_/CLK _35133_/D VGND VGND VPWR VPWR _35133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32345_ _33635_/CLK _32345_/D VGND VGND VPWR VPWR _32345_/Q sky130_fd_sc_hd__dfxtp_1
X_17279_ _17063_/X _17277_/X _17278_/X _17067_/X VGND VGND VPWR VPWR _17279_/X sky130_fd_sc_hd__a22o_1
XFILLER_101_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19018_ _35744_/Q _35104_/Q _34464_/Q _33824_/Q _18734_/X _18735_/X VGND VGND VPWR
+ VPWR _19018_/X sky130_fd_sc_hd__mux4_1
X_35064_ _35577_/CLK _35064_/D VGND VGND VPWR VPWR _35064_/Q sky130_fd_sc_hd__dfxtp_1
X_20290_ _35588_/Q _35524_/Q _35460_/Q _35396_/Q _20256_/X _20257_/X VGND VGND VPWR
+ VPWR _20290_/X sky130_fd_sc_hd__mux4_1
XFILLER_161_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32276_ _36191_/CLK _32276_/D VGND VGND VPWR VPWR _32276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34015_ _34016_/CLK _34015_/D VGND VGND VPWR VPWR _34015_/Q sky130_fd_sc_hd__dfxtp_1
X_31227_ _31227_/A VGND VGND VPWR VPWR _35830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31158_ _35798_/Q input63/X _31160_/S VGND VGND VPWR VPWR _31159_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30109_ _35301_/Q _29123_/X _30121_/S VGND VGND VPWR VPWR _30110_/A sky130_fd_sc_hd__mux2_1
X_23980_ _23980_/A VGND VGND VPWR VPWR _32528_/D sky130_fd_sc_hd__clkbuf_1
X_35966_ _35966_/CLK _35966_/D VGND VGND VPWR VPWR _35966_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31089_ _31089_/A VGND VGND VPWR VPWR _35765_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34917_ _35042_/CLK _34917_/D VGND VGND VPWR VPWR _34917_/Q sky130_fd_sc_hd__dfxtp_1
X_22931_ _22931_/A VGND VGND VPWR VPWR _32030_/D sky130_fd_sc_hd__clkbuf_1
X_35897_ _36025_/CLK _35897_/D VGND VGND VPWR VPWR _35897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25650_ _33252_/Q _24314_/X _25664_/S VGND VGND VPWR VPWR _25651_/A sky130_fd_sc_hd__mux2_1
X_22862_ _35597_/Q _35533_/Q _35469_/Q _35405_/Q _20605_/X _20607_/X VGND VGND VPWR
+ VPWR _22862_/X sky130_fd_sc_hd__mux4_1
X_34848_ _35038_/CLK _34848_/D VGND VGND VPWR VPWR _34848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24601_ _24601_/A VGND VGND VPWR VPWR _32790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21813_ _21663_/X _21811_/X _21812_/X _21667_/X VGND VGND VPWR VPWR _21813_/X sky130_fd_sc_hd__a22o_1
X_25581_ _33221_/Q _24416_/X _25589_/S VGND VGND VPWR VPWR _25582_/A sky130_fd_sc_hd__mux2_1
X_22793_ _33291_/Q _36171_/Q _33163_/Q _33099_/Q _20628_/X _21757_/A VGND VGND VPWR
+ VPWR _22793_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34779_ _34779_/CLK _34779_/D VGND VGND VPWR VPWR _34779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27320_ _34011_/Q _24286_/X _27332_/S VGND VGND VPWR VPWR _27321_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24532_ _23007_/X _32759_/Q _24548_/S VGND VGND VPWR VPWR _24533_/A sky130_fd_sc_hd__mux2_1
X_21744_ _35564_/Q _35500_/Q _35436_/Q _35372_/Q _21497_/X _21498_/X VGND VGND VPWR
+ VPWR _21744_/X sky130_fd_sc_hd__mux4_1
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27251_ _27251_/A VGND VGND VPWR VPWR _33978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24463_ _24463_/A VGND VGND VPWR VPWR _32726_/D sky130_fd_sc_hd__clkbuf_1
X_21675_ _22532_/A VGND VGND VPWR VPWR _21675_/X sky130_fd_sc_hd__buf_4
XFILLER_184_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26202_ _25075_/X _33513_/Q _26206_/S VGND VGND VPWR VPWR _26203_/A sky130_fd_sc_hd__mux2_1
X_23414_ _23414_/A VGND VGND VPWR VPWR _32265_/D sky130_fd_sc_hd__clkbuf_1
X_20626_ _22508_/A VGND VGND VPWR VPWR _20626_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24394_ input43/X VGND VGND VPWR VPWR _24394_/X sky130_fd_sc_hd__clkbuf_4
X_27182_ _27182_/A VGND VGND VPWR VPWR _33945_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26133_ _26133_/A VGND VGND VPWR VPWR _33480_/D sky130_fd_sc_hd__clkbuf_1
X_23345_ input60/X VGND VGND VPWR VPWR _23345_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_22_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20557_ _19454_/A _20555_/X _20556_/X _19459_/A VGND VGND VPWR VPWR _20557_/X sky130_fd_sc_hd__a22o_1
XFILLER_123_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26064_ _26064_/A VGND VGND VPWR VPWR _33447_/D sky130_fd_sc_hd__clkbuf_1
X_23276_ _23276_/A VGND VGND VPWR VPWR _32209_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20488_ _33547_/Q _33483_/Q _33419_/Q _33355_/Q _18333_/X _18335_/X VGND VGND VPWR
+ VPWR _20488_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25015_ _25015_/A VGND VGND VPWR VPWR _32981_/D sky130_fd_sc_hd__clkbuf_1
X_22227_ _33274_/Q _36154_/Q _33146_/Q _33082_/Q _22011_/X _22012_/X VGND VGND VPWR
+ VPWR _22227_/X sky130_fd_sc_hd__mux4_1
XTAP_6801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29823_ _29823_/A VGND VGND VPWR VPWR _35165_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22158_ _22511_/A VGND VGND VPWR VPWR _22158_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21109_ _35802_/Q _32177_/Q _35674_/Q _35610_/Q _20854_/X _20855_/X VGND VGND VPWR
+ VPWR _21109_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29754_ _35133_/Q _29197_/X _29758_/S VGND VGND VPWR VPWR _29755_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22089_ _22442_/A VGND VGND VPWR VPWR _22089_/X sky130_fd_sc_hd__clkbuf_4
X_26966_ _26965_/X _33852_/Q _26975_/S VGND VGND VPWR VPWR _26967_/A sky130_fd_sc_hd__mux2_1
XTAP_6889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28705_ _26912_/X _34667_/Q _28705_/S VGND VGND VPWR VPWR _28706_/A sky130_fd_sc_hd__mux2_1
X_25917_ _26007_/S VGND VGND VPWR VPWR _25936_/S sky130_fd_sc_hd__buf_4
XFILLER_130_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29685_ _35100_/Q _29095_/X _29695_/S VGND VGND VPWR VPWR _29686_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26897_ input17/X VGND VGND VPWR VPWR _26897_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_207_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28636_ _28636_/A VGND VGND VPWR VPWR _34634_/D sky130_fd_sc_hd__clkbuf_1
X_16650_ _16646_/X _16647_/X _16648_/X _16649_/X VGND VGND VPWR VPWR _16650_/X sky130_fd_sc_hd__a22o_1
XFILLER_75_866 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25848_ _25150_/X _33345_/Q _25864_/S VGND VGND VPWR VPWR _25849_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16581_ _16577_/X _16580_/X _16441_/X VGND VGND VPWR VPWR _16591_/C sky130_fd_sc_hd__o21ba_1
X_28567_ _28567_/A VGND VGND VPWR VPWR _34601_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25779_ _25779_/A VGND VGND VPWR VPWR _33312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18320_ _20202_/A VGND VGND VPWR VPWR _18320_/X sky130_fd_sc_hd__buf_4
X_27518_ _26956_/X _34105_/Q _27530_/S VGND VGND VPWR VPWR _27519_/A sky130_fd_sc_hd__mux2_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28498_ _27005_/X _34569_/Q _28498_/S VGND VGND VPWR VPWR _28499_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18251_ _18247_/X _18250_/X _17834_/A VGND VGND VPWR VPWR _18273_/A sky130_fd_sc_hd__o21ba_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27449_ _26853_/X _34072_/Q _27467_/S VGND VGND VPWR VPWR _27450_/A sky130_fd_sc_hd__mux2_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17202_ _17908_/A VGND VGND VPWR VPWR _17202_/X sky130_fd_sc_hd__clkbuf_4
X_18182_ _18178_/X _18181_/X _17867_/A VGND VGND VPWR VPWR _18183_/D sky130_fd_sc_hd__o21ba_1
X_30460_ _30460_/A VGND VGND VPWR VPWR _35467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17133_ _32492_/Q _32364_/Q _32044_/Q _36012_/Q _16923_/X _17064_/X VGND VGND VPWR
+ VPWR _17133_/X sky130_fd_sc_hd__mux4_1
X_29119_ _29119_/A VGND VGND VPWR VPWR _34851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30391_ _30391_/A VGND VGND VPWR VPWR _35434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32130_ _35750_/CLK _32130_/D VGND VGND VPWR VPWR _32130_/Q sky130_fd_sc_hd__dfxtp_1
X_17064_ _17770_/A VGND VGND VPWR VPWR _17064_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16015_ _16057_/A VGND VGND VPWR VPWR _17978_/A sky130_fd_sc_hd__buf_12
X_32061_ _36028_/CLK _32061_/D VGND VGND VPWR VPWR _32061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31012_ _31012_/A VGND VGND VPWR VPWR _35728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35820_ _35950_/CLK _35820_/D VGND VGND VPWR VPWR _35820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17966_ _35075_/Q _35011_/Q _34947_/Q _34883_/Q _17862_/X _17863_/X VGND VGND VPWR
+ VPWR _17966_/X sky130_fd_sc_hd__mux4_1
XFILLER_112_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19705_ _34036_/Q _33972_/Q _33908_/Q _32244_/Q _19673_/X _19674_/X VGND VGND VPWR
+ VPWR _19705_/X sky130_fd_sc_hd__mux4_1
X_16917_ _16849_/X _16915_/X _16916_/X _16852_/X VGND VGND VPWR VPWR _16917_/X sky130_fd_sc_hd__a22o_1
X_32963_ _33026_/CLK _32963_/D VGND VGND VPWR VPWR _32963_/Q sky130_fd_sc_hd__dfxtp_1
X_35751_ _35879_/CLK _35751_/D VGND VGND VPWR VPWR _35751_/Q sky130_fd_sc_hd__dfxtp_1
X_17897_ _17860_/X _17895_/X _17896_/X _17865_/X VGND VGND VPWR VPWR _17897_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34702_ _35280_/CLK _34702_/D VGND VGND VPWR VPWR _34702_/Q sky130_fd_sc_hd__dfxtp_1
X_31914_ _31914_/A VGND VGND VPWR VPWR _36156_/D sky130_fd_sc_hd__clkbuf_1
X_19636_ _19502_/X _19634_/X _19635_/X _19505_/X VGND VGND VPWR VPWR _19636_/X sky130_fd_sc_hd__a22o_1
X_16848_ _16842_/X _16845_/X _16846_/X _16847_/X VGND VGND VPWR VPWR _16848_/X sky130_fd_sc_hd__a22o_1
X_32894_ _32959_/CLK _32894_/D VGND VGND VPWR VPWR _32894_/Q sky130_fd_sc_hd__dfxtp_1
X_35682_ _35811_/CLK _35682_/D VGND VGND VPWR VPWR _35682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34633_ _35337_/CLK _34633_/D VGND VGND VPWR VPWR _34633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31845_ _31845_/A VGND VGND VPWR VPWR _36123_/D sky130_fd_sc_hd__clkbuf_1
X_19567_ _19495_/X _19565_/X _19566_/X _19500_/X VGND VGND VPWR VPWR _19567_/X sky130_fd_sc_hd__a22o_1
X_16779_ _16702_/X _16777_/X _16778_/X _16708_/X VGND VGND VPWR VPWR _16779_/X sky130_fd_sc_hd__a22o_1
XFILLER_207_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18518_ _32466_/Q _32338_/Q _32018_/Q _35986_/Q _18517_/X _20163_/A VGND VGND VPWR
+ VPWR _18518_/X sky130_fd_sc_hd__mux4_1
X_34564_ _35332_/CLK _34564_/D VGND VGND VPWR VPWR _34564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31776_ _36091_/Q input40/X _31784_/S VGND VGND VPWR VPWR _31777_/A sky130_fd_sc_hd__mux2_1
X_19498_ _33774_/Q _33710_/Q _33646_/Q _33582_/Q _19496_/X _19497_/X VGND VGND VPWR
+ VPWR _19498_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30727_ _35594_/Q _29237_/X _30733_/S VGND VGND VPWR VPWR _30728_/A sky130_fd_sc_hd__mux2_1
X_18449_ _32720_/Q _32656_/Q _32592_/Q _36048_/Q _20162_/A _20013_/A VGND VGND VPWR
+ VPWR _18449_/X sky130_fd_sc_hd__mux4_1
X_33515_ _35257_/CLK _33515_/D VGND VGND VPWR VPWR _33515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34495_ _35837_/CLK _34495_/D VGND VGND VPWR VPWR _34495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36234_ _36237_/CLK _36234_/D VGND VGND VPWR VPWR _36234_/Q sky130_fd_sc_hd__dfxtp_1
X_33446_ _35991_/CLK _33446_/D VGND VGND VPWR VPWR _33446_/Q sky130_fd_sc_hd__dfxtp_1
X_21460_ _21310_/X _21458_/X _21459_/X _21314_/X VGND VGND VPWR VPWR _21460_/X sky130_fd_sc_hd__a22o_1
X_30658_ _35561_/Q _29135_/X _30662_/S VGND VGND VPWR VPWR _30659_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20411_ _18277_/X _20409_/X _20410_/X _18287_/X VGND VGND VPWR VPWR _20411_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36165_ _36165_/CLK _36165_/D VGND VGND VPWR VPWR _36165_/Q sky130_fd_sc_hd__dfxtp_1
X_33377_ _34266_/CLK _33377_/D VGND VGND VPWR VPWR _33377_/Q sky130_fd_sc_hd__dfxtp_1
X_21391_ _35554_/Q _35490_/Q _35426_/Q _35362_/Q _21144_/X _21145_/X VGND VGND VPWR
+ VPWR _21391_/X sky130_fd_sc_hd__mux4_1
X_30589_ _30589_/A VGND VGND VPWR VPWR _35528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23130_ input6/X VGND VGND VPWR VPWR _23130_/X sky130_fd_sc_hd__buf_6
X_32328_ _35334_/CLK _32328_/D VGND VGND VPWR VPWR _32328_/Q sky130_fd_sc_hd__dfxtp_1
X_20342_ _32774_/Q _32710_/Q _32646_/Q _36102_/Q _20278_/X _20062_/X VGND VGND VPWR
+ VPWR _20342_/X sky130_fd_sc_hd__mux4_1
X_35116_ _35950_/CLK _35116_/D VGND VGND VPWR VPWR _35116_/Q sky130_fd_sc_hd__dfxtp_1
X_36096_ _36098_/CLK _36096_/D VGND VGND VPWR VPWR _36096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23061_ _23061_/A VGND VGND VPWR VPWR _32072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35047_ _35943_/CLK _35047_/D VGND VGND VPWR VPWR _35047_/Q sky130_fd_sc_hd__dfxtp_1
X_20273_ _20201_/X _20271_/X _20272_/X _20206_/X VGND VGND VPWR VPWR _20273_/X sky130_fd_sc_hd__a22o_1
X_32259_ _34057_/CLK _32259_/D VGND VGND VPWR VPWR _32259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22012_ _22370_/A VGND VGND VPWR VPWR _22012_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26820_ _26820_/A VGND VGND VPWR VPWR _33805_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26751_ _33772_/Q _24338_/X _26769_/S VGND VGND VPWR VPWR _26752_/A sky130_fd_sc_hd__mux2_1
X_23963_ _23963_/A VGND VGND VPWR VPWR _32521_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35949_ _35949_/CLK _35949_/D VGND VGND VPWR VPWR _35949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25702_ _33277_/Q _24391_/X _25706_/S VGND VGND VPWR VPWR _25703_/A sky130_fd_sc_hd__mux2_1
X_29470_ _23270_/X _34998_/Q _29488_/S VGND VGND VPWR VPWR _29471_/A sky130_fd_sc_hd__mux2_1
X_22914_ input3/X VGND VGND VPWR VPWR _22914_/X sky130_fd_sc_hd__buf_4
X_26682_ _26682_/A VGND VGND VPWR VPWR _33740_/D sky130_fd_sc_hd__clkbuf_1
X_23894_ _23894_/A VGND VGND VPWR VPWR _32488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28421_ _26891_/X _34532_/Q _28435_/S VGND VGND VPWR VPWR _28422_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25633_ _33244_/Q _24289_/X _25643_/S VGND VGND VPWR VPWR _25634_/A sky130_fd_sc_hd__mux2_1
X_22845_ _33805_/Q _33741_/Q _33677_/Q _33613_/Q _20620_/X _20621_/X VGND VGND VPWR
+ VPWR _22845_/X sky130_fd_sc_hd__mux4_1
XFILLER_216_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28352_ _28352_/A VGND VGND VPWR VPWR _34499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25564_ _33213_/Q _24391_/X _25568_/S VGND VGND VPWR VPWR _25565_/A sky130_fd_sc_hd__mux2_1
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22776_ _34826_/Q _34762_/Q _34698_/Q _34634_/Q _22594_/X _22595_/X VGND VGND VPWR
+ VPWR _22776_/X sky130_fd_sc_hd__mux4_1
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27303_ _34003_/Q _24261_/X _27311_/S VGND VGND VPWR VPWR _27304_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24515_ _22982_/X _32751_/Q _24527_/S VGND VGND VPWR VPWR _24516_/A sky130_fd_sc_hd__mux2_1
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28283_ _28283_/A VGND VGND VPWR VPWR _34466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21727_ _21449_/X _21725_/X _21726_/X _21452_/X VGND VGND VPWR VPWR _21727_/X sky130_fd_sc_hd__a22o_1
XFILLER_212_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25495_ _33180_/Q _24289_/X _25505_/S VGND VGND VPWR VPWR _25496_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27234_ _27234_/A VGND VGND VPWR VPWR _33970_/D sky130_fd_sc_hd__clkbuf_1
X_24446_ _22875_/X _32718_/Q _24464_/S VGND VGND VPWR VPWR _24447_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_1171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21658_ _22582_/A VGND VGND VPWR VPWR _21658_/X sky130_fd_sc_hd__buf_6
XFILLER_32_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27165_ _27165_/A VGND VGND VPWR VPWR _33937_/D sky130_fd_sc_hd__clkbuf_1
X_20609_ _20597_/X _20600_/X _20603_/X _20608_/X VGND VGND VPWR VPWR _20609_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24377_ _32696_/Q _24376_/X _24398_/S VGND VGND VPWR VPWR _24378_/A sky130_fd_sc_hd__mux2_1
X_21589_ _22429_/A VGND VGND VPWR VPWR _21589_/X sky130_fd_sc_hd__buf_8
XFILLER_137_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26116_ _25146_/X _33472_/Q _26134_/S VGND VGND VPWR VPWR _26117_/A sky130_fd_sc_hd__mux2_1
X_23328_ _32227_/Q _23327_/X _23334_/S VGND VGND VPWR VPWR _23329_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27096_ _26931_/X _33905_/Q _27104_/S VGND VGND VPWR VPWR _27097_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26047_ _26047_/A VGND VGND VPWR VPWR _33439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23259_ _32204_/Q _23220_/X _23350_/S VGND VGND VPWR VPWR _23260_/A sky130_fd_sc_hd__mux2_1
XFILLER_238_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17820_ _34559_/Q _32447_/Q _34431_/Q _34367_/Q _17578_/X _17579_/X VGND VGND VPWR
+ VPWR _17820_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29806_ _29806_/A VGND VGND VPWR VPWR _35157_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27998_ _27998_/A VGND VGND VPWR VPWR _34331_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17751_ _17747_/X _17750_/X _17514_/X VGND VGND VPWR VPWR _17752_/D sky130_fd_sc_hd__o21ba_1
XFILLER_130_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_1445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26949_ _26949_/A VGND VGND VPWR VPWR _33846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29737_ _35125_/Q _29172_/X _29737_/S VGND VGND VPWR VPWR _29738_/A sky130_fd_sc_hd__mux2_1
XTAP_5974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16702_ _17901_/A VGND VGND VPWR VPWR _16702_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_207_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29668_ _35092_/Q _29070_/X _29674_/S VGND VGND VPWR VPWR _29669_/A sky130_fd_sc_hd__mux2_1
X_17682_ _17682_/A _17682_/B _17682_/C _17682_/D VGND VGND VPWR VPWR _17683_/A sky130_fd_sc_hd__or4_1
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19421_ _34284_/Q _34220_/Q _34156_/Q _34092_/Q _19389_/X _19390_/X VGND VGND VPWR
+ VPWR _19421_/X sky130_fd_sc_hd__mux4_1
X_28619_ _26984_/X _34626_/Q _28633_/S VGND VGND VPWR VPWR _28620_/A sky130_fd_sc_hd__mux2_1
X_16633_ _33246_/Q _36126_/Q _33118_/Q _33054_/Q _16352_/X _16353_/X VGND VGND VPWR
+ VPWR _16633_/X sky130_fd_sc_hd__mux4_1
X_29599_ _29599_/A VGND VGND VPWR VPWR _35059_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31630_ _31678_/S VGND VGND VPWR VPWR _31649_/S sky130_fd_sc_hd__buf_4
X_19352_ _34026_/Q _33962_/Q _33898_/Q _32234_/Q _19320_/X _19321_/X VGND VGND VPWR
+ VPWR _19352_/X sky130_fd_sc_hd__mux4_1
X_16564_ _16496_/X _16562_/X _16563_/X _16499_/X VGND VGND VPWR VPWR _16564_/X sky130_fd_sc_hd__a22o_1
XFILLER_222_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18303_ _20211_/A VGND VGND VPWR VPWR _18303_/X sky130_fd_sc_hd__buf_4
XFILLER_206_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31561_ _35989_/Q input62/X _31565_/S VGND VGND VPWR VPWR _31562_/A sky130_fd_sc_hd__mux2_1
X_19283_ _19149_/X _19281_/X _19282_/X _19152_/X VGND VGND VPWR VPWR _19283_/X sky130_fd_sc_hd__a22o_1
X_16495_ _16489_/X _16492_/X _16493_/X _16494_/X VGND VGND VPWR VPWR _16495_/X sky130_fd_sc_hd__a22o_1
XFILLER_241_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33300_ _36237_/CLK _33300_/D VGND VGND VPWR VPWR _33300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18234_ _15997_/X _18232_/X _18233_/X _16003_/X VGND VGND VPWR VPWR _18234_/X sky130_fd_sc_hd__a22o_1
X_30512_ _30512_/A VGND VGND VPWR VPWR _35491_/D sky130_fd_sc_hd__clkbuf_1
X_34280_ _34870_/CLK _34280_/D VGND VGND VPWR VPWR _34280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31492_ _31492_/A VGND VGND VPWR VPWR _35956_/D sky130_fd_sc_hd__clkbuf_1
X_33231_ _34124_/CLK _33231_/D VGND VGND VPWR VPWR _33231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18165_ _32522_/Q _32394_/Q _32074_/Q _36042_/Q _17982_/X _17007_/A VGND VGND VPWR
+ VPWR _18165_/X sky130_fd_sc_hd__mux4_1
X_30443_ _23313_/X _35459_/Q _30455_/S VGND VGND VPWR VPWR _30444_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17116_ _16801_/X _17114_/X _17115_/X _16806_/X VGND VGND VPWR VPWR _17116_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33162_ _36172_/CLK _33162_/D VGND VGND VPWR VPWR _33162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18096_ _34312_/Q _34248_/Q _34184_/Q _34120_/Q _17795_/X _17796_/X VGND VGND VPWR
+ VPWR _18096_/X sky130_fd_sc_hd__mux4_1
X_30374_ _23148_/X _35426_/Q _30392_/S VGND VGND VPWR VPWR _30375_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32113_ _35552_/CLK _32113_/D VGND VGND VPWR VPWR _32113_/Q sky130_fd_sc_hd__dfxtp_1
X_17047_ _17047_/A VGND VGND VPWR VPWR _31977_/D sky130_fd_sc_hd__clkbuf_1
X_33093_ _36100_/CLK _33093_/D VGND VGND VPWR VPWR _33093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32044_ _36077_/CLK _32044_/D VGND VGND VPWR VPWR _32044_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ _33504_/Q _33440_/Q _33376_/Q _33312_/Q _18717_/X _18718_/X VGND VGND VPWR
+ VPWR _18998_/X sky130_fd_sc_hd__mux4_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35803_ _35803_/CLK _35803_/D VGND VGND VPWR VPWR _35803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17949_ _32515_/Q _32387_/Q _32067_/Q _36035_/Q _17629_/X _17770_/X VGND VGND VPWR
+ VPWR _17949_/X sky130_fd_sc_hd__mux4_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33995_ _35273_/CLK _33995_/D VGND VGND VPWR VPWR _33995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35734_ _35925_/CLK _35734_/D VGND VGND VPWR VPWR _35734_/Q sky130_fd_sc_hd__dfxtp_1
X_20960_ _32982_/Q _32918_/Q _32854_/Q _32790_/Q _20883_/X _20884_/X VGND VGND VPWR
+ VPWR _20960_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_1248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32946_ _35765_/CLK _32946_/D VGND VGND VPWR VPWR _32946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19619_ _33201_/Q _32561_/Q _35953_/Q _35889_/Q _19374_/X _19375_/X VGND VGND VPWR
+ VPWR _19619_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35665_ _35666_/CLK _35665_/D VGND VGND VPWR VPWR _35665_/Q sky130_fd_sc_hd__dfxtp_1
X_20891_ _22458_/A VGND VGND VPWR VPWR _20891_/X sky130_fd_sc_hd__buf_4
X_32877_ _36015_/CLK _32877_/D VGND VGND VPWR VPWR _32877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22630_ _35077_/Q _35013_/Q _34949_/Q _34885_/Q _22462_/X _22463_/X VGND VGND VPWR
+ VPWR _22630_/X sky130_fd_sc_hd__mux4_1
XFILLER_59_1160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34616_ _35318_/CLK _34616_/D VGND VGND VPWR VPWR _34616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31828_ _31828_/A VGND VGND VPWR VPWR _36115_/D sky130_fd_sc_hd__clkbuf_1
X_35596_ _35852_/CLK _35596_/D VGND VGND VPWR VPWR _35596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22561_ _22555_/X _22560_/X _22453_/X VGND VGND VPWR VPWR _22569_/C sky130_fd_sc_hd__o21ba_1
XFILLER_34_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31759_ _36083_/Q input31/X _31763_/S VGND VGND VPWR VPWR _31760_/A sky130_fd_sc_hd__mux2_1
X_34547_ _34997_/CLK _34547_/D VGND VGND VPWR VPWR _34547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21512_ _33766_/Q _33702_/Q _33638_/Q _33574_/Q _21443_/X _21444_/X VGND VGND VPWR
+ VPWR _21512_/X sky130_fd_sc_hd__mux4_1
X_24300_ _24300_/A VGND VGND VPWR VPWR _32671_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22492_ _34817_/Q _34753_/Q _34689_/Q _34625_/Q _22241_/X _22242_/X VGND VGND VPWR
+ VPWR _22492_/X sky130_fd_sc_hd__mux4_1
XFILLER_210_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25280_ _25280_/A VGND VGND VPWR VPWR _33080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34478_ _35758_/CLK _34478_/D VGND VGND VPWR VPWR _34478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24231_ _24231_/A VGND VGND VPWR VPWR _32647_/D sky130_fd_sc_hd__clkbuf_1
X_36217_ _36220_/CLK _36217_/D VGND VGND VPWR VPWR _36217_/Q sky130_fd_sc_hd__dfxtp_1
X_21443_ _22502_/A VGND VGND VPWR VPWR _21443_/X sky130_fd_sc_hd__buf_4
X_33429_ _34001_/CLK _33429_/D VGND VGND VPWR VPWR _33429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24162_ _24162_/A VGND VGND VPWR VPWR _32614_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36148_ _36149_/CLK _36148_/D VGND VGND VPWR VPWR _36148_/Q sky130_fd_sc_hd__dfxtp_1
X_21374_ _21096_/X _21372_/X _21373_/X _21099_/X VGND VGND VPWR VPWR _21374_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23113_ _23113_/A VGND VGND VPWR VPWR _32150_/D sky130_fd_sc_hd__clkbuf_1
X_20325_ _20321_/X _20324_/X _20153_/X VGND VGND VPWR VPWR _20333_/C sky130_fd_sc_hd__o21ba_1
X_24093_ _24093_/A VGND VGND VPWR VPWR _32582_/D sky130_fd_sc_hd__clkbuf_1
X_28970_ _28970_/A VGND VGND VPWR VPWR _34792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36079_ _36080_/CLK _36079_/D VGND VGND VPWR VPWR _36079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23044_ input49/X VGND VGND VPWR VPWR _23044_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_66_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27921_ _34295_/Q _24373_/X _27937_/S VGND VGND VPWR VPWR _27922_/A sky130_fd_sc_hd__mux2_1
X_20256_ _20256_/A VGND VGND VPWR VPWR _20256_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_115_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27852_ _27852_/A VGND VGND VPWR VPWR _34262_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20187_ _20000_/X _20185_/X _20186_/X _20003_/X VGND VGND VPWR VPWR _20187_/X sky130_fd_sc_hd__a22o_1
XFILLER_27_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26803_ _33797_/Q _24416_/X _26811_/S VGND VGND VPWR VPWR _26804_/A sky130_fd_sc_hd__mux2_1
XTAP_5248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27783_ _27831_/S VGND VGND VPWR VPWR _27802_/S sky130_fd_sc_hd__buf_4
XFILLER_170_1470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24995_ input12/X VGND VGND VPWR VPWR _24995_/X sky130_fd_sc_hd__buf_4
XFILLER_217_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29522_ _29522_/A VGND VGND VPWR VPWR _35022_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26734_ _33764_/Q _24314_/X _26748_/S VGND VGND VPWR VPWR _26735_/A sky130_fd_sc_hd__mux2_1
X_23946_ _23038_/X _32513_/Q _23962_/S VGND VGND VPWR VPWR _23947_/A sky130_fd_sc_hd__mux2_1
XTAP_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_983 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_802 _22892_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29453_ _23244_/X _34990_/Q _29467_/S VGND VGND VPWR VPWR _29454_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_6_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_6_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_26665_ _25159_/X _33732_/Q _26675_/S VGND VGND VPWR VPWR _26666_/A sky130_fd_sc_hd__mux2_1
XFILLER_232_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_813 _22917_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_824 _23105_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23877_ _23877_/A VGND VGND VPWR VPWR _32480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28404_ _26866_/X _34524_/Q _28414_/S VGND VGND VPWR VPWR _28405_/A sky130_fd_sc_hd__mux2_1
XANTENNA_835 _23346_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_846 _23688_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25616_ _33236_/Q _24264_/X _25622_/S VGND VGND VPWR VPWR _25617_/A sky130_fd_sc_hd__mux2_1
X_29384_ _29384_/A _30465_/B VGND VGND VPWR VPWR _29517_/S sky130_fd_sc_hd__nand2_8
X_22828_ _22824_/X _22827_/X _22442_/A _22443_/A VGND VGND VPWR VPWR _22843_/B sky130_fd_sc_hd__o211a_1
XANTENNA_857 _24345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26596_ _25057_/X _33699_/Q _26612_/S VGND VGND VPWR VPWR _26597_/A sky130_fd_sc_hd__mux2_1
XANTENNA_868 _24577_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_879 _25084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28335_ _28335_/A VGND VGND VPWR VPWR _34491_/D sky130_fd_sc_hd__clkbuf_1
X_25547_ _33205_/Q _24366_/X _25547_/S VGND VGND VPWR VPWR _25548_/A sky130_fd_sc_hd__mux2_1
X_22759_ _34058_/Q _33994_/Q _33930_/Q _32266_/Q _20658_/X _20660_/X VGND VGND VPWR
+ VPWR _22759_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16280_ _33236_/Q _36116_/Q _33108_/Q _33044_/Q _16020_/X _16021_/X VGND VGND VPWR
+ VPWR _16280_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28266_ _28266_/A VGND VGND VPWR VPWR _34458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25478_ _33172_/Q _24264_/X _25484_/S VGND VGND VPWR VPWR _25479_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27217_ _27217_/A VGND VGND VPWR VPWR _33962_/D sky130_fd_sc_hd__clkbuf_1
X_24429_ _32713_/Q _24428_/X _24429_/S VGND VGND VPWR VPWR _24430_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28197_ _26959_/X _34426_/Q _28207_/S VGND VGND VPWR VPWR _28198_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27148_ _27008_/X _33930_/Q _27154_/S VGND VGND VPWR VPWR _27149_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19970_ _19647_/X _19968_/X _19969_/X _19650_/X VGND VGND VPWR VPWR _19970_/X sky130_fd_sc_hd__a22o_1
X_27079_ _26906_/X _33897_/Q _27083_/S VGND VGND VPWR VPWR _27080_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_860 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1078 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18921_ _18748_/X _18919_/X _18920_/X _18753_/X VGND VGND VPWR VPWR _18921_/X sky130_fd_sc_hd__a22o_1
XTAP_7140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30090_ _35292_/Q _29095_/X _30100_/S VGND VGND VPWR VPWR _30091_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_1212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1201 _23102_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1212 _23327_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1223 _24304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1234 _24577_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18852_ _18743_/X _18850_/X _18851_/X _18746_/X VGND VGND VPWR VPWR _18852_/X sky130_fd_sc_hd__a22o_1
XTAP_6450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1245 _26142_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1256 _27289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1267 _29787_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17803_ _32767_/Q _32703_/Q _32639_/Q _36095_/Q _17625_/X _17762_/X VGND VGND VPWR
+ VPWR _17803_/X sky130_fd_sc_hd__mux4_1
XTAP_6494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1278 _17860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18783_ _34521_/Q _32409_/Q _34393_/Q _34329_/Q _18466_/X _18467_/X VGND VGND VPWR
+ VPWR _18783_/X sky130_fd_sc_hd__mux4_1
XTAP_5760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15995_ _15995_/A VGND VGND VPWR VPWR _17769_/A sky130_fd_sc_hd__buf_2
XANTENNA_1289 _17847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17734_ _32509_/Q _32381_/Q _32061_/Q _36029_/Q _17629_/X _17417_/X VGND VGND VPWR
+ VPWR _17734_/X sky130_fd_sc_hd__mux4_1
X_32800_ _36065_/CLK _32800_/D VGND VGND VPWR VPWR _32800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30992_ _30992_/A VGND VGND VPWR VPWR _35719_/D sky130_fd_sc_hd__clkbuf_1
X_33780_ _33780_/CLK _33780_/D VGND VGND VPWR VPWR _33780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17665_ _17661_/X _17664_/X _17489_/X _17490_/X VGND VGND VPWR VPWR _17682_/B sky130_fd_sc_hd__o211a_1
X_32731_ _36059_/CLK _32731_/D VGND VGND VPWR VPWR _32731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19404_ _35819_/Q _32196_/Q _35691_/Q _35627_/Q _19260_/X _19261_/X VGND VGND VPWR
+ VPWR _19404_/X sky130_fd_sc_hd__mux4_1
X_16616_ _34781_/Q _34717_/Q _34653_/Q _34589_/Q _16582_/X _16583_/X VGND VGND VPWR
+ VPWR _16616_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32662_ _36119_/CLK _32662_/D VGND VGND VPWR VPWR _32662_/Q sky130_fd_sc_hd__dfxtp_1
X_35450_ _35578_/CLK _35450_/D VGND VGND VPWR VPWR _35450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17596_ _32505_/Q _32377_/Q _32057_/Q _36025_/Q _17276_/X _17417_/X VGND VGND VPWR
+ VPWR _17596_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34401_ _35039_/CLK _34401_/D VGND VGND VPWR VPWR _34401_/Q sky130_fd_sc_hd__dfxtp_1
X_31613_ _31613_/A VGND VGND VPWR VPWR _36013_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19335_ _35561_/Q _35497_/Q _35433_/Q _35369_/Q _19197_/X _19198_/X VGND VGND VPWR
+ VPWR _19335_/X sky130_fd_sc_hd__mux4_1
X_16547_ _33179_/Q _32539_/Q _35931_/Q _35867_/Q _16368_/X _16369_/X VGND VGND VPWR
+ VPWR _16547_/X sky130_fd_sc_hd__mux4_1
X_32593_ _36050_/CLK _32593_/D VGND VGND VPWR VPWR _32593_/Q sky130_fd_sc_hd__dfxtp_1
X_35381_ _36021_/CLK _35381_/D VGND VGND VPWR VPWR _35381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31544_ _31544_/A VGND VGND VPWR VPWR _35981_/D sky130_fd_sc_hd__clkbuf_1
X_34332_ _35166_/CLK _34332_/D VGND VGND VPWR VPWR _34332_/Q sky130_fd_sc_hd__dfxtp_1
X_19266_ _33191_/Q _32551_/Q _35943_/Q _35879_/Q _19021_/X _19022_/X VGND VGND VPWR
+ VPWR _19266_/X sky130_fd_sc_hd__mux4_1
X_16478_ _16293_/X _16476_/X _16477_/X _16296_/X VGND VGND VPWR VPWR _16478_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18217_ _16014_/X _18215_/X _18216_/X _16023_/X VGND VGND VPWR VPWR _18217_/X sky130_fd_sc_hd__a22o_1
X_34263_ _35664_/CLK _34263_/D VGND VGND VPWR VPWR _34263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19197_ _20256_/A VGND VGND VPWR VPWR _19197_/X sky130_fd_sc_hd__buf_4
X_31475_ _23237_/X _35948_/Q _31493_/S VGND VGND VPWR VPWR _31476_/A sky130_fd_sc_hd__mux2_1
X_33214_ _35903_/CLK _33214_/D VGND VGND VPWR VPWR _33214_/Q sky130_fd_sc_hd__dfxtp_1
X_36002_ _36003_/CLK _36002_/D VGND VGND VPWR VPWR _36002_/Q sky130_fd_sc_hd__dfxtp_1
X_18148_ _17855_/X _18146_/X _18147_/X _17858_/X VGND VGND VPWR VPWR _18148_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30426_ _23286_/X _35451_/Q _30434_/S VGND VGND VPWR VPWR _30427_/A sky130_fd_sc_hd__mux2_1
X_34194_ _34194_/CLK _34194_/D VGND VGND VPWR VPWR _34194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33145_ _36090_/CLK _33145_/D VGND VGND VPWR VPWR _33145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18079_ _35847_/Q _32227_/Q _35719_/Q _35655_/Q _15989_/X _15991_/X VGND VGND VPWR
+ VPWR _18079_/X sky130_fd_sc_hd__mux4_1
X_30357_ _23124_/X _35418_/Q _30371_/S VGND VGND VPWR VPWR _30358_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20110_ _35839_/Q _32218_/Q _35711_/Q _35647_/Q _19966_/X _19967_/X VGND VGND VPWR
+ VPWR _20110_/X sky130_fd_sc_hd__mux4_1
X_33076_ _36149_/CLK _33076_/D VGND VGND VPWR VPWR _33076_/Q sky130_fd_sc_hd__dfxtp_1
X_21090_ _22502_/A VGND VGND VPWR VPWR _21090_/X sky130_fd_sc_hd__buf_6
X_30288_ _35386_/Q _29188_/X _30298_/S VGND VGND VPWR VPWR _30289_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_1142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20041_ _35581_/Q _35517_/Q _35453_/Q _35389_/Q _19903_/X _19904_/X VGND VGND VPWR
+ VPWR _20041_/X sky130_fd_sc_hd__mux4_1
X_32027_ _35995_/CLK _32027_/D VGND VGND VPWR VPWR _32027_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_140_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _35981_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23800_ _23800_/A VGND VGND VPWR VPWR _32444_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24780_ _24780_/A VGND VGND VPWR VPWR _32874_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33978_ _36154_/CLK _33978_/D VGND VGND VPWR VPWR _33978_/Q sky130_fd_sc_hd__dfxtp_1
X_21992_ _34803_/Q _34739_/Q _34675_/Q _34611_/Q _21888_/X _21889_/X VGND VGND VPWR
+ VPWR _21992_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35717_ _35849_/CLK _35717_/D VGND VGND VPWR VPWR _35717_/Q sky130_fd_sc_hd__dfxtp_1
X_23731_ _23731_/A VGND VGND VPWR VPWR _32411_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20943_ _34262_/Q _34198_/Q _34134_/Q _34070_/Q _20605_/X _20607_/X VGND VGND VPWR
+ VPWR _20943_/X sky130_fd_sc_hd__mux4_1
XANTENNA_109 _32129_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32929_ _36001_/CLK _32929_/D VGND VGND VPWR VPWR _32929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26450_ _26450_/A VGND VGND VPWR VPWR _33630_/D sky130_fd_sc_hd__clkbuf_1
X_35648_ _35715_/CLK _35648_/D VGND VGND VPWR VPWR _35648_/Q sky130_fd_sc_hd__dfxtp_1
X_23662_ _23662_/A VGND VGND VPWR VPWR _32380_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20874_ _20736_/X _20872_/X _20873_/X _20741_/X VGND VGND VPWR VPWR _20874_/X sky130_fd_sc_hd__a22o_1
XFILLER_74_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25401_ _25401_/A VGND VGND VPWR VPWR _33137_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22613_ _33285_/Q _36165_/Q _33157_/Q _33093_/Q _22364_/X _22365_/X VGND VGND VPWR
+ VPWR _22613_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_1282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26381_ _25140_/X _33598_/Q _26383_/S VGND VGND VPWR VPWR _26382_/A sky130_fd_sc_hd__mux2_1
X_35579_ _35579_/CLK _35579_/D VGND VGND VPWR VPWR _35579_/Q sky130_fd_sc_hd__dfxtp_1
X_23593_ _23593_/A VGND VGND VPWR VPWR _32347_/D sky130_fd_sc_hd__clkbuf_1
X_28120_ _28120_/A VGND VGND VPWR VPWR _34389_/D sky130_fd_sc_hd__clkbuf_1
X_25332_ _25332_/A VGND VGND VPWR VPWR _33104_/D sky130_fd_sc_hd__clkbuf_1
X_22544_ _22508_/X _22542_/X _22543_/X _22511_/X VGND VGND VPWR VPWR _22544_/X sky130_fd_sc_hd__a22o_1
XFILLER_202_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28051_ _26943_/X _34357_/Q _28051_/S VGND VGND VPWR VPWR _28052_/A sky130_fd_sc_hd__mux2_1
X_25263_ _25263_/A VGND VGND VPWR VPWR _33072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22475_ _34049_/Q _33985_/Q _33921_/Q _32257_/Q _22326_/X _22327_/X VGND VGND VPWR
+ VPWR _22475_/X sky130_fd_sc_hd__mux4_1
XFILLER_241_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27002_ input54/X VGND VGND VPWR VPWR _27002_/X sky130_fd_sc_hd__buf_4
XFILLER_194_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24214_ _24214_/A VGND VGND VPWR VPWR _32639_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21426_ _35811_/Q _32187_/Q _35683_/Q _35619_/Q _21207_/X _21208_/X VGND VGND VPWR
+ VPWR _21426_/X sky130_fd_sc_hd__mux4_1
X_25194_ _25194_/A VGND VGND VPWR VPWR _33039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21357_ _21353_/X _21356_/X _21041_/X VGND VGND VPWR VPWR _21365_/C sky130_fd_sc_hd__o21ba_1
X_24145_ _24145_/A VGND VGND VPWR VPWR _32606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20308_ _33541_/Q _33477_/Q _33413_/Q _33349_/Q _20129_/X _20130_/X VGND VGND VPWR
+ VPWR _20308_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24076_ _24076_/A VGND VGND VPWR VPWR _32574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21288_ _21043_/X _21286_/X _21287_/X _21046_/X VGND VGND VPWR VPWR _21288_/X sky130_fd_sc_hd__a22o_1
X_28953_ _28953_/A VGND VGND VPWR VPWR _34784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20239_ _33795_/Q _33731_/Q _33667_/Q _33603_/Q _20202_/X _20203_/X VGND VGND VPWR
+ VPWR _20239_/X sky130_fd_sc_hd__mux4_1
X_23027_ _23027_/A VGND VGND VPWR VPWR _32061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27904_ _34287_/Q _24348_/X _27916_/S VGND VGND VPWR VPWR _27905_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28884_ _28911_/S VGND VGND VPWR VPWR _28903_/S sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_131_CLK clkbuf_6_23__f_CLK/X VGND VGND VPWR VPWR _34256_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_5001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27835_ _34254_/Q _24244_/X _27853_/S VGND VGND VPWR VPWR _27836_/A sky130_fd_sc_hd__mux2_1
XTAP_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27766_ _27766_/A VGND VGND VPWR VPWR _34221_/D sky130_fd_sc_hd__clkbuf_1
X_24978_ _24978_/A VGND VGND VPWR VPWR _32968_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29505_ _23327_/X _35015_/Q _29509_/S VGND VGND VPWR VPWR _29506_/A sky130_fd_sc_hd__mux2_1
XTAP_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26717_ _33756_/Q _24289_/X _26727_/S VGND VGND VPWR VPWR _26718_/A sky130_fd_sc_hd__mux2_1
XTAP_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23929_ _23013_/X _32505_/Q _23941_/S VGND VGND VPWR VPWR _23930_/A sky130_fd_sc_hd__mux2_1
XTAP_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27697_ _27697_/A VGND VGND VPWR VPWR _34189_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_610 _18504_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_621 _18571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_632 _18961_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29436_ _23217_/X _34982_/Q _29446_/S VGND VGND VPWR VPWR _29437_/A sky130_fd_sc_hd__mux2_1
X_17450_ _32757_/Q _32693_/Q _32629_/Q _36085_/Q _17272_/X _17409_/X VGND VGND VPWR
+ VPWR _17450_/X sky130_fd_sc_hd__mux4_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26648_ _25134_/X _33724_/Q _26654_/S VGND VGND VPWR VPWR _26649_/A sky130_fd_sc_hd__mux2_1
XTAP_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_643 _19387_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_654 _20270_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16401_ _35543_/Q _35479_/Q _35415_/Q _35351_/Q _16191_/X _16192_/X VGND VGND VPWR
+ VPWR _16401_/X sky130_fd_sc_hd__mux4_1
XANTENNA_665 _22396_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_676 _22556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29367_ _29367_/A VGND VGND VPWR VPWR _34949_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_687 _22508_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17381_ _32499_/Q _32371_/Q _32051_/Q _36019_/Q _17276_/X _17064_/X VGND VGND VPWR
+ VPWR _17381_/X sky130_fd_sc_hd__mux4_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_198_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _35710_/CLK sky130_fd_sc_hd__clkbuf_16
X_26579_ _25032_/X _33691_/Q _26591_/S VGND VGND VPWR VPWR _26580_/A sky130_fd_sc_hd__mux2_1
XANTENNA_698 _22458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19120_ _33251_/Q _36131_/Q _33123_/Q _33059_/Q _19005_/X _19006_/X VGND VGND VPWR
+ VPWR _19120_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16332_ _16328_/X _16331_/X _16071_/X VGND VGND VPWR VPWR _16340_/C sky130_fd_sc_hd__o21ba_1
X_28318_ _28318_/A VGND VGND VPWR VPWR _34483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29298_ _29298_/A VGND VGND VPWR VPWR _34916_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19051_ _35809_/Q _32185_/Q _35681_/Q _35617_/Q _18907_/X _18908_/X VGND VGND VPWR
+ VPWR _19051_/X sky130_fd_sc_hd__mux4_1
X_28249_ _28249_/A VGND VGND VPWR VPWR _34450_/D sky130_fd_sc_hd__clkbuf_1
X_16263_ _34771_/Q _34707_/Q _34643_/Q _34579_/Q _16229_/X _16230_/X VGND VGND VPWR
+ VPWR _16263_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18002_ _17998_/X _18001_/X _17867_/X VGND VGND VPWR VPWR _18003_/D sky130_fd_sc_hd__o21ba_1
X_31260_ _31260_/A VGND VGND VPWR VPWR _35846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16194_ _33169_/Q _32529_/Q _35921_/Q _35857_/Q _16063_/X _16065_/X VGND VGND VPWR
+ VPWR _16194_/X sky130_fd_sc_hd__mux4_1
XFILLER_126_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30211_ _30211_/A VGND VGND VPWR VPWR _35349_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_370_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _33009_/CLK sky130_fd_sc_hd__clkbuf_16
X_31191_ _31191_/A VGND VGND VPWR VPWR _35813_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30142_ _35317_/Q _29172_/X _30142_/S VGND VGND VPWR VPWR _30143_/A sky130_fd_sc_hd__mux2_1
X_19953_ _34299_/Q _34235_/Q _34171_/Q _34107_/Q _19742_/X _19743_/X VGND VGND VPWR
+ VPWR _19953_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18904_ _32989_/Q _32925_/Q _32861_/Q _32797_/Q _18583_/X _18584_/X VGND VGND VPWR
+ VPWR _18904_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_122_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _36237_/CLK sky130_fd_sc_hd__clkbuf_16
X_34950_ _35080_/CLK _34950_/D VGND VGND VPWR VPWR _34950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30073_ _35284_/Q _29070_/X _30079_/S VGND VGND VPWR VPWR _30074_/A sky130_fd_sc_hd__mux2_1
XANTENNA_1020 _17847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19884_ _19884_/A _19884_/B _19884_/C _19884_/D VGND VGND VPWR VPWR _19885_/A sky130_fd_sc_hd__or4_4
XANTENNA_1031 _17865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1042 _17154_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1053 _16135_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33901_ _35958_/CLK _33901_/D VGND VGND VPWR VPWR _33901_/Q sky130_fd_sc_hd__dfxtp_1
X_18835_ _33243_/Q _36123_/Q _33115_/Q _33051_/Q _18652_/X _18653_/X VGND VGND VPWR
+ VPWR _18835_/X sky130_fd_sc_hd__mux4_1
X_34881_ _35075_/CLK _34881_/D VGND VGND VPWR VPWR _34881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1064 _16841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1075 _17164_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1086 _17232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1097 _17298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_212_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33832_ _35943_/CLK _33832_/D VGND VGND VPWR VPWR _33832_/Q sky130_fd_sc_hd__dfxtp_1
X_15978_ input65/X VGND VGND VPWR VPWR _16057_/A sky130_fd_sc_hd__buf_8
XFILLER_222_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18766_ _32729_/Q _32665_/Q _32601_/Q _36057_/Q _18513_/X _18650_/X VGND VGND VPWR
+ VPWR _18766_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17717_ _35068_/Q _35004_/Q _34940_/Q _34876_/Q _17509_/X _17510_/X VGND VGND VPWR
+ VPWR _17717_/X sky130_fd_sc_hd__mux4_1
X_30975_ _30975_/A VGND VGND VPWR VPWR _35711_/D sky130_fd_sc_hd__clkbuf_1
X_33763_ _34276_/CLK _33763_/D VGND VGND VPWR VPWR _33763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18697_ _18693_/X _18696_/X _18340_/X _18342_/X VGND VGND VPWR VPWR _18712_/B sky130_fd_sc_hd__o211a_1
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35502_ _35949_/CLK _35502_/D VGND VGND VPWR VPWR _35502_/Q sky130_fd_sc_hd__dfxtp_1
X_32714_ _36170_/CLK _32714_/D VGND VGND VPWR VPWR _32714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17648_ _17507_/X _17646_/X _17647_/X _17512_/X VGND VGND VPWR VPWR _17648_/X sky130_fd_sc_hd__a22o_1
XFILLER_51_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33694_ _34017_/CLK _33694_/D VGND VGND VPWR VPWR _33694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35433_ _35819_/CLK _35433_/D VGND VGND VPWR VPWR _35433_/Q sky130_fd_sc_hd__dfxtp_1
X_32645_ _36103_/CLK _32645_/D VGND VGND VPWR VPWR _32645_/Q sky130_fd_sc_hd__dfxtp_1
X_17579_ _17932_/A VGND VGND VPWR VPWR _17579_/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_189_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _35580_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_189_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19318_ _19142_/X _19316_/X _19317_/X _19147_/X VGND VGND VPWR VPWR _19318_/X sky130_fd_sc_hd__a22o_1
X_20590_ _20659_/A VGND VGND VPWR VPWR _22396_/A sky130_fd_sc_hd__buf_12
X_32576_ _35906_/CLK _32576_/D VGND VGND VPWR VPWR _32576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35364_ _35555_/CLK _35364_/D VGND VGND VPWR VPWR _35364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34315_ _35273_/CLK _34315_/D VGND VGND VPWR VPWR _34315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31527_ _23319_/X _35973_/Q _31535_/S VGND VGND VPWR VPWR _31528_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19249_ _33511_/Q _33447_/Q _33383_/Q _33319_/Q _19070_/X _19071_/X VGND VGND VPWR
+ VPWR _19249_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35295_ _35296_/CLK _35295_/D VGND VGND VPWR VPWR _35295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22260_ _33275_/Q _36155_/Q _33147_/Q _33083_/Q _22011_/X _22012_/X VGND VGND VPWR
+ VPWR _22260_/X sky130_fd_sc_hd__mux4_1
X_34246_ _34310_/CLK _34246_/D VGND VGND VPWR VPWR _34246_/Q sky130_fd_sc_hd__dfxtp_1
X_31458_ _23175_/X _35940_/Q _31472_/S VGND VGND VPWR VPWR _31459_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21211_ _20888_/X _21209_/X _21210_/X _20891_/X VGND VGND VPWR VPWR _21211_/X sky130_fd_sc_hd__a22o_1
X_30409_ _23261_/X _35443_/Q _30413_/S VGND VGND VPWR VPWR _30410_/A sky130_fd_sc_hd__mux2_1
X_34177_ _36160_/CLK _34177_/D VGND VGND VPWR VPWR _34177_/Q sky130_fd_sc_hd__dfxtp_1
X_22191_ _22155_/X _22189_/X _22190_/X _22158_/X VGND VGND VPWR VPWR _22191_/X sky130_fd_sc_hd__a22o_1
X_31389_ _31389_/A VGND VGND VPWR VPWR _35907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_361_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _34286_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_219_1248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21142_ _35739_/Q _35099_/Q _34459_/Q _33819_/Q _21034_/X _21035_/X VGND VGND VPWR
+ VPWR _21142_/X sky130_fd_sc_hd__mux4_1
X_33128_ _33255_/CLK _33128_/D VGND VGND VPWR VPWR _33128_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_113_CLK clkbuf_6_20__f_CLK/X VGND VGND VPWR VPWR _35281_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_1243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25950_ _25950_/A VGND VGND VPWR VPWR _33393_/D sky130_fd_sc_hd__clkbuf_1
X_21073_ _35801_/Q _32176_/Q _35673_/Q _35609_/Q _20854_/X _20855_/X VGND VGND VPWR
+ VPWR _21073_/X sky130_fd_sc_hd__mux4_1
X_33059_ _36130_/CLK _33059_/D VGND VGND VPWR VPWR _33059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20024_ _19848_/X _20022_/X _20023_/X _19853_/X VGND VGND VPWR VPWR _20024_/X sky130_fd_sc_hd__a22o_1
X_24901_ _24901_/A VGND VGND VPWR VPWR _32931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25881_ _25881_/A VGND VGND VPWR VPWR _33360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27620_ _27620_/A VGND VGND VPWR VPWR _34152_/D sky130_fd_sc_hd__clkbuf_1
X_24832_ _23044_/X _32899_/Q _24844_/S VGND VGND VPWR VPWR _24833_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27551_ _27005_/X _34121_/Q _27551_/S VGND VGND VPWR VPWR _27552_/A sky130_fd_sc_hd__mux2_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24763_ _22941_/X _32866_/Q _24781_/S VGND VGND VPWR VPWR _24764_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21975_ _34035_/Q _33971_/Q _33907_/Q _32243_/Q _21973_/X _21974_/X VGND VGND VPWR
+ VPWR _21975_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26502_ _25119_/X _33655_/Q _26518_/S VGND VGND VPWR VPWR _26503_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23714_ _23714_/A VGND VGND VPWR VPWR _32403_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20926_ _35797_/Q _32172_/Q _35669_/Q _35605_/Q _20854_/X _20855_/X VGND VGND VPWR
+ VPWR _20926_/X sky130_fd_sc_hd__mux4_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27482_ _26903_/X _34088_/Q _27488_/S VGND VGND VPWR VPWR _27483_/A sky130_fd_sc_hd__mux2_1
X_24694_ _24694_/A VGND VGND VPWR VPWR _32834_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29221_ _29221_/A VGND VGND VPWR VPWR _34884_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26433_ _26433_/A VGND VGND VPWR VPWR _33622_/D sky130_fd_sc_hd__clkbuf_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23645_ _23645_/A VGND VGND VPWR VPWR _32372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20857_ _35731_/Q _35091_/Q _34451_/Q _33811_/Q _20649_/X _20651_/X VGND VGND VPWR
+ VPWR _20857_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29152_ _34862_/Q _29151_/X _29173_/S VGND VGND VPWR VPWR _29153_/A sky130_fd_sc_hd__mux2_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26364_ _26412_/S VGND VGND VPWR VPWR _26383_/S sky130_fd_sc_hd__buf_4
XFILLER_161_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23576_ _23576_/A VGND VGND VPWR VPWR _32339_/D sky130_fd_sc_hd__clkbuf_1
X_20788_ _35793_/Q _32167_/Q _35665_/Q _35601_/Q _20645_/X _20646_/X VGND VGND VPWR
+ VPWR _20788_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28103_ _28778_/B _31410_/B VGND VGND VPWR VPWR _28236_/S sky130_fd_sc_hd__nand2_8
XFILLER_70_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25315_ _25315_/A VGND VGND VPWR VPWR _33097_/D sky130_fd_sc_hd__clkbuf_1
X_22527_ _22523_/X _22526_/X _22453_/X VGND VGND VPWR VPWR _22537_/C sky130_fd_sc_hd__o21ba_1
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29083_ _29247_/S VGND VGND VPWR VPWR _29111_/S sky130_fd_sc_hd__buf_4
X_26295_ _25013_/X _33557_/Q _26299_/S VGND VGND VPWR VPWR _26296_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28034_ _28034_/A VGND VGND VPWR VPWR _34348_/D sky130_fd_sc_hd__clkbuf_1
X_25246_ _25246_/A VGND VGND VPWR VPWR _33064_/D sky130_fd_sc_hd__clkbuf_1
X_22458_ _22458_/A VGND VGND VPWR VPWR _22458_/X sky130_fd_sc_hd__buf_4
XFILLER_210_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21409_ _21400_/X _21407_/X _21408_/X VGND VGND VPWR VPWR _21410_/D sky130_fd_sc_hd__o21ba_1
X_25177_ input57/X VGND VGND VPWR VPWR _25177_/X sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_352_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _36149_/CLK sky130_fd_sc_hd__clkbuf_16
X_22389_ _35070_/Q _35006_/Q _34942_/Q _34878_/Q _22109_/X _22110_/X VGND VGND VPWR
+ VPWR _22389_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24128_ _24128_/A VGND VGND VPWR VPWR _32598_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29985_ _29985_/A VGND VGND VPWR VPWR _35242_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_104_CLK clkbuf_leaf_80_CLK/A VGND VGND VPWR VPWR _35729_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_1340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28936_ _34776_/Q _24276_/X _28954_/S VGND VGND VPWR VPWR _28937_/A sky130_fd_sc_hd__mux2_1
X_16950_ _34023_/Q _33959_/Q _33895_/Q _32204_/Q _16667_/X _16668_/X VGND VGND VPWR
+ VPWR _16950_/X sky130_fd_sc_hd__mux4_1
X_24059_ _23003_/X _32566_/Q _24077_/S VGND VGND VPWR VPWR _24060_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16881_ _34277_/Q _34213_/Q _34149_/Q _34085_/Q _16736_/X _16737_/X VGND VGND VPWR
+ VPWR _16881_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28867_ _28867_/A VGND VGND VPWR VPWR _34743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_238_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18620_ _33237_/Q _36117_/Q _33109_/Q _33045_/Q _18320_/X _18321_/X VGND VGND VPWR
+ VPWR _18620_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27818_ _27818_/A VGND VGND VPWR VPWR _34246_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28798_ _26850_/X _34711_/Q _28798_/S VGND VGND VPWR VPWR _28799_/A sky130_fd_sc_hd__mux2_1
XTAP_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ _32979_/Q _32915_/Q _32851_/Q _32787_/Q _18333_/X _18335_/X VGND VGND VPWR
+ VPWR _18551_/X sky130_fd_sc_hd__mux4_1
XTAP_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27749_ _27749_/A VGND VGND VPWR VPWR _34213_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17502_ _17855_/A VGND VGND VPWR VPWR _17502_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18482_ _33233_/Q _36113_/Q _33105_/Q _33041_/Q _18320_/X _18321_/X VGND VGND VPWR
+ VPWR _18482_/X sky130_fd_sc_hd__mux4_1
XTAP_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30760_ _23121_/X _35609_/Q _30776_/S VGND VGND VPWR VPWR _30761_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_440 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_451 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _35316_/Q _35252_/Q _35188_/Q _32308_/Q _17359_/X _17360_/X VGND VGND VPWR
+ VPWR _17433_/X sky130_fd_sc_hd__mux4_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_462 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29419_ _23136_/X _34974_/Q _29425_/S VGND VGND VPWR VPWR _29420_/A sky130_fd_sc_hd__mux2_1
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_473 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30691_ _30691_/A VGND VGND VPWR VPWR _35576_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_484 _31994_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_495 _31997_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32430_ _35054_/CLK _32430_/D VGND VGND VPWR VPWR _32430_/Q sky130_fd_sc_hd__dfxtp_1
X_17364_ _35058_/Q _34994_/Q _34930_/Q _34866_/Q _17156_/X _17157_/X VGND VGND VPWR
+ VPWR _17364_/X sky130_fd_sc_hd__mux4_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16315_ _17847_/A VGND VGND VPWR VPWR _16315_/X sky130_fd_sc_hd__buf_6
X_19103_ _20162_/A VGND VGND VPWR VPWR _19103_/X sky130_fd_sc_hd__buf_4
XFILLER_201_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32361_ _34792_/CLK _32361_/D VGND VGND VPWR VPWR _32361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17295_ _17154_/X _17293_/X _17294_/X _17159_/X VGND VGND VPWR VPWR _17295_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31312_ _35871_/Q input9/X _31316_/S VGND VGND VPWR VPWR _31313_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19034_ _19034_/A VGND VGND VPWR VPWR _32096_/D sky130_fd_sc_hd__clkbuf_1
X_34100_ _34228_/CLK _34100_/D VGND VGND VPWR VPWR _34100_/Q sky130_fd_sc_hd__dfxtp_1
X_35080_ _35080_/CLK _35080_/D VGND VGND VPWR VPWR _35080_/Q sky130_fd_sc_hd__dfxtp_1
X_16246_ _16242_/X _16245_/X _16011_/X VGND VGND VPWR VPWR _16270_/A sky130_fd_sc_hd__o21ba_1
XFILLER_9_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32292_ _36003_/CLK _32292_/D VGND VGND VPWR VPWR _32292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34031_ _34032_/CLK _34031_/D VGND VGND VPWR VPWR _34031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31243_ _31243_/A VGND VGND VPWR VPWR _35838_/D sky130_fd_sc_hd__clkbuf_1
X_16177_ _33489_/Q _33425_/Q _33361_/Q _33297_/Q _15998_/X _15999_/X VGND VGND VPWR
+ VPWR _16177_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_343_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _34295_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_217_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput105 _31973_/Q VGND VGND VPWR VPWR D1[23] sky130_fd_sc_hd__buf_2
XFILLER_126_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput116 _31983_/Q VGND VGND VPWR VPWR D1[33] sky130_fd_sc_hd__buf_2
XFILLER_86_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput127 _31993_/Q VGND VGND VPWR VPWR D1[43] sky130_fd_sc_hd__buf_2
XFILLER_99_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput138 _32003_/Q VGND VGND VPWR VPWR D1[53] sky130_fd_sc_hd__buf_2
XFILLER_217_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31174_ _31174_/A VGND VGND VPWR VPWR _35805_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput149 _32013_/Q VGND VGND VPWR VPWR D1[63] sky130_fd_sc_hd__buf_2
XFILLER_88_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30125_ _30125_/A VGND VGND VPWR VPWR _35308_/D sky130_fd_sc_hd__clkbuf_1
X_19936_ _19647_/X _19934_/X _19935_/X _19650_/X VGND VGND VPWR VPWR _19936_/X sky130_fd_sc_hd__a22o_1
X_35982_ _35982_/CLK _35982_/D VGND VGND VPWR VPWR _35982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_991 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30056_ _30056_/A VGND VGND VPWR VPWR _35276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34933_ _35061_/CLK _34933_/D VGND VGND VPWR VPWR _34933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19867_ _19863_/X _19866_/X _19789_/X _19790_/X VGND VGND VPWR VPWR _19884_/B sky130_fd_sc_hd__o211a_1
XFILLER_233_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18818_ _18743_/X _18816_/X _18817_/X _18746_/X VGND VGND VPWR VPWR _18818_/X sky130_fd_sc_hd__a22o_1
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34864_ _35760_/CLK _34864_/D VGND VGND VPWR VPWR _34864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19798_ _33206_/Q _32566_/Q _35958_/Q _35894_/Q _19727_/X _19728_/X VGND VGND VPWR
+ VPWR _19798_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33815_ _35667_/CLK _33815_/D VGND VGND VPWR VPWR _33815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18749_ _34520_/Q _32408_/Q _34392_/Q _34328_/Q _18466_/X _18467_/X VGND VGND VPWR
+ VPWR _18749_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34795_ _36011_/CLK _34795_/D VGND VGND VPWR VPWR _34795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33746_ _34194_/CLK _33746_/D VGND VGND VPWR VPWR _33746_/Q sky130_fd_sc_hd__dfxtp_1
X_21760_ _21754_/X _21755_/X _21758_/X _21759_/X VGND VGND VPWR VPWR _21760_/X sky130_fd_sc_hd__a22o_1
X_30958_ _35703_/Q _29179_/X _30974_/S VGND VGND VPWR VPWR _30959_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20711_ _20597_/X _20707_/X _20710_/X _20603_/X VGND VGND VPWR VPWR _20711_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33677_ _36112_/CLK _33677_/D VGND VGND VPWR VPWR _33677_/Q sky130_fd_sc_hd__dfxtp_1
X_21691_ _34283_/Q _34219_/Q _34155_/Q _34091_/Q _21689_/X _21690_/X VGND VGND VPWR
+ VPWR _21691_/X sky130_fd_sc_hd__mux4_1
X_30889_ _30889_/A VGND VGND VPWR VPWR _35670_/D sky130_fd_sc_hd__clkbuf_1
X_23430_ _22883_/X _32271_/Q _23446_/S VGND VGND VPWR VPWR _23431_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35416_ _35864_/CLK _35416_/D VGND VGND VPWR VPWR _35416_/Q sky130_fd_sc_hd__dfxtp_1
X_20642_ _22443_/A VGND VGND VPWR VPWR _20642_/X sky130_fd_sc_hd__buf_2
X_32628_ _36085_/CLK _32628_/D VGND VGND VPWR VPWR _32628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20573_ _20573_/A _20573_/B _20573_/C _20573_/D VGND VGND VPWR VPWR _20574_/A sky130_fd_sc_hd__or4_1
X_35347_ _35925_/CLK _35347_/D VGND VGND VPWR VPWR _35347_/Q sky130_fd_sc_hd__dfxtp_1
X_23361_ _32240_/Q _23250_/X _23371_/S VGND VGND VPWR VPWR _23362_/A sky130_fd_sc_hd__mux2_1
X_32559_ _35952_/CLK _32559_/D VGND VGND VPWR VPWR _32559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25100_ input29/X VGND VGND VPWR VPWR _25100_/X sky130_fd_sc_hd__buf_2
X_22312_ _22312_/A VGND VGND VPWR VPWR _22312_/X sky130_fd_sc_hd__buf_6
XFILLER_191_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26080_ _25094_/X _33455_/Q _26092_/S VGND VGND VPWR VPWR _26081_/A sky130_fd_sc_hd__mux2_1
X_35278_ _36216_/CLK _35278_/D VGND VGND VPWR VPWR _35278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23292_ _32215_/Q _23223_/X _23350_/S VGND VGND VPWR VPWR _23293_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25031_ _25031_/A VGND VGND VPWR VPWR _32986_/D sky130_fd_sc_hd__clkbuf_1
X_22243_ _34810_/Q _34746_/Q _34682_/Q _34618_/Q _22241_/X _22242_/X VGND VGND VPWR
+ VPWR _22243_/X sky130_fd_sc_hd__mux4_1
X_34229_ _34229_/CLK _34229_/D VGND VGND VPWR VPWR _34229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_334_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _36089_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_192_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22174_ _22170_/X _22173_/X _22100_/X VGND VGND VPWR VPWR _22184_/C sky130_fd_sc_hd__o21ba_1
XFILLER_117_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21125_ _21125_/A _21125_/B _21125_/C _21125_/D VGND VGND VPWR VPWR _21126_/A sky130_fd_sc_hd__or4_2
X_29770_ _29770_/A VGND VGND VPWR VPWR _35140_/D sky130_fd_sc_hd__clkbuf_1
X_26982_ _26981_/X _33857_/Q _27006_/S VGND VGND VPWR VPWR _26983_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25933_ _25933_/A VGND VGND VPWR VPWR _33385_/D sky130_fd_sc_hd__clkbuf_1
X_28721_ _28721_/A VGND VGND VPWR VPWR _34674_/D sky130_fd_sc_hd__clkbuf_1
X_21056_ _21047_/X _21054_/X _21055_/X VGND VGND VPWR VPWR _21057_/D sky130_fd_sc_hd__o21ba_1
XFILLER_86_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20007_ _33212_/Q _32572_/Q _35964_/Q _35900_/Q _19727_/X _19728_/X VGND VGND VPWR
+ VPWR _20007_/X sky130_fd_sc_hd__mux4_1
X_28652_ _28652_/A VGND VGND VPWR VPWR _34641_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25864_ _25174_/X _33353_/Q _25864_/S VGND VGND VPWR VPWR _25865_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24815_ _23019_/X _32891_/Q _24823_/S VGND VGND VPWR VPWR _24816_/A sky130_fd_sc_hd__mux2_1
X_27603_ _27603_/A VGND VGND VPWR VPWR _34144_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28583_ _26931_/X _34609_/Q _28591_/S VGND VGND VPWR VPWR _28584_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25795_ _25072_/X _33320_/Q _25801_/S VGND VGND VPWR VPWR _25796_/A sky130_fd_sc_hd__mux2_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27534_ _27534_/A VGND VGND VPWR VPWR _34112_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24746_ _22917_/X _32858_/Q _24760_/S VGND VGND VPWR VPWR _24747_/A sky130_fd_sc_hd__mux2_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21958_ _34802_/Q _34738_/Q _34674_/Q _34610_/Q _21888_/X _21889_/X VGND VGND VPWR
+ VPWR _21958_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20909_ _20909_/A VGND VGND VPWR VPWR _36180_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27465_ _26878_/X _34080_/Q _27467_/S VGND VGND VPWR VPWR _27466_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24677_ _24677_/A VGND VGND VPWR VPWR _32826_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21889_ _22595_/A VGND VGND VPWR VPWR _21889_/X sky130_fd_sc_hd__buf_4
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26416_ _24989_/X _33614_/Q _26434_/S VGND VGND VPWR VPWR _26417_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29204_ _34879_/Q _29203_/X _29204_/S VGND VGND VPWR VPWR _29205_/A sky130_fd_sc_hd__mux2_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23628_ _32364_/Q _23237_/X _23646_/S VGND VGND VPWR VPWR _23629_/A sky130_fd_sc_hd__mux2_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27396_ _27396_/A VGND VGND VPWR VPWR _34047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29135_ input20/X VGND VGND VPWR VPWR _29135_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_167_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26347_ _26347_/A VGND VGND VPWR VPWR _33581_/D sky130_fd_sc_hd__clkbuf_1
X_23559_ _23074_/X _32333_/Q _23559_/S VGND VGND VPWR VPWR _23560_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16100_ _17867_/A VGND VGND VPWR VPWR _16100_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_156_836 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput18 DW[25] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__buf_4
X_29066_ _29066_/A VGND VGND VPWR VPWR _34834_/D sky130_fd_sc_hd__clkbuf_1
Xinput29 DW[35] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__buf_4
X_17080_ _35306_/Q _35242_/Q _35178_/Q _32298_/Q _17006_/X _17007_/X VGND VGND VPWR
+ VPWR _17080_/X sky130_fd_sc_hd__mux4_1
X_26278_ _26278_/A VGND VGND VPWR VPWR _33549_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16031_ _32462_/Q _32334_/Q _32014_/Q _35982_/Q _16028_/X _17863_/A VGND VGND VPWR
+ VPWR _16031_/X sky130_fd_sc_hd__mux4_1
X_28017_ _28017_/A VGND VGND VPWR VPWR _34340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25229_ _25229_/A VGND VGND VPWR VPWR _33056_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_325_CLK clkbuf_6_44__f_CLK/X VGND VGND VPWR VPWR _35828_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17982_ _17982_/A VGND VGND VPWR VPWR _17982_/X sky130_fd_sc_hd__buf_6
X_29968_ _35234_/Q _29113_/X _29986_/S VGND VGND VPWR VPWR _29969_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19721_ _19716_/X _19718_/X _19719_/X _19720_/X VGND VGND VPWR VPWR _19721_/X sky130_fd_sc_hd__a22o_1
X_28919_ _34768_/Q _24252_/X _28933_/S VGND VGND VPWR VPWR _28920_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16933_ _16646_/X _16931_/X _16932_/X _16649_/X VGND VGND VPWR VPWR _16933_/X sky130_fd_sc_hd__a22o_1
X_29899_ _29899_/A VGND VGND VPWR VPWR _35201_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31930_ _23316_/X _36164_/Q _31940_/S VGND VGND VPWR VPWR _31931_/A sky130_fd_sc_hd__mux2_1
X_19652_ _20160_/A VGND VGND VPWR VPWR _19652_/X sky130_fd_sc_hd__clkbuf_8
X_16864_ _16641_/X _16862_/X _16863_/X _16644_/X VGND VGND VPWR VPWR _16864_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18603_ _18374_/X _18599_/X _18602_/X _18384_/X VGND VGND VPWR VPWR _18603_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16795_ _16790_/X _16793_/X _16794_/X VGND VGND VPWR VPWR _16810_/C sky130_fd_sc_hd__o21ba_1
XFILLER_24_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19583_ _19294_/X _19581_/X _19582_/X _19297_/X VGND VGND VPWR VPWR _19583_/X sky130_fd_sc_hd__a22o_1
X_31861_ _23152_/X _36131_/Q _31877_/S VGND VGND VPWR VPWR _31862_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33600_ _34305_/CLK _33600_/D VGND VGND VPWR VPWR _33600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18534_ _34514_/Q _32402_/Q _34386_/Q _34322_/Q _18466_/X _18467_/X VGND VGND VPWR
+ VPWR _18534_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30812_ _23256_/X _35634_/Q _30818_/S VGND VGND VPWR VPWR _30813_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31792_ _31792_/A VGND VGND VPWR VPWR _36098_/D sky130_fd_sc_hd__clkbuf_1
X_34580_ _34775_/CLK _34580_/D VGND VGND VPWR VPWR _34580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33531_ _33723_/CLK _33531_/D VGND VGND VPWR VPWR _33531_/Q sky130_fd_sc_hd__dfxtp_1
X_18465_ _18374_/X _18463_/X _18464_/X _18384_/X VGND VGND VPWR VPWR _18465_/X sky130_fd_sc_hd__a22o_1
X_30743_ _23096_/X _35601_/Q _30755_/S VGND VGND VPWR VPWR _30744_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_270 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_281 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_292 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17416_ _17908_/A VGND VGND VPWR VPWR _17416_/X sky130_fd_sc_hd__clkbuf_4
X_18396_ _20073_/A VGND VGND VPWR VPWR _19459_/A sky130_fd_sc_hd__buf_12
X_33462_ _34297_/CLK _33462_/D VGND VGND VPWR VPWR _33462_/Q sky130_fd_sc_hd__dfxtp_1
X_30674_ _30674_/A VGND VGND VPWR VPWR _35568_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35201_ _35330_/CLK _35201_/D VGND VGND VPWR VPWR _35201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32413_ _35036_/CLK _32413_/D VGND VGND VPWR VPWR _32413_/Q sky130_fd_sc_hd__dfxtp_1
X_17347_ _17855_/A VGND VGND VPWR VPWR _17347_/X sky130_fd_sc_hd__buf_4
XFILLER_202_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36181_ _36202_/CLK _36181_/D VGND VGND VPWR VPWR _36181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33393_ _34033_/CLK _33393_/D VGND VGND VPWR VPWR _33393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35132_ _35772_/CLK _35132_/D VGND VGND VPWR VPWR _35132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32344_ _36121_/CLK _32344_/D VGND VGND VPWR VPWR _32344_/Q sky130_fd_sc_hd__dfxtp_1
X_17278_ _33008_/Q _32944_/Q _32880_/Q _32816_/Q _16989_/X _16990_/X VGND VGND VPWR
+ VPWR _17278_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16229_ _17994_/A VGND VGND VPWR VPWR _16229_/X sky130_fd_sc_hd__buf_6
X_19017_ _35808_/Q _32184_/Q _35680_/Q _35616_/Q _18907_/X _18908_/X VGND VGND VPWR
+ VPWR _19017_/X sky130_fd_sc_hd__mux4_1
X_32275_ _36211_/CLK _32275_/D VGND VGND VPWR VPWR _32275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_316_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _35766_/CLK sky130_fd_sc_hd__clkbuf_16
X_35063_ _35257_/CLK _35063_/D VGND VGND VPWR VPWR _35063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34014_ _34205_/CLK _34014_/D VGND VGND VPWR VPWR _34014_/Q sky130_fd_sc_hd__dfxtp_1
X_31226_ _35830_/Q input35/X _31244_/S VGND VGND VPWR VPWR _31227_/A sky130_fd_sc_hd__mux2_1
X_31157_ _31157_/A VGND VGND VPWR VPWR _35797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30108_ _30108_/A VGND VGND VPWR VPWR _35300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19919_ _34298_/Q _34234_/Q _34170_/Q _34106_/Q _19742_/X _19743_/X VGND VGND VPWR
+ VPWR _19919_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35965_ _35965_/CLK _35965_/D VGND VGND VPWR VPWR _35965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31088_ _35765_/Q _29172_/X _31088_/S VGND VGND VPWR VPWR _31089_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30039_ _35268_/Q _29219_/X _30049_/S VGND VGND VPWR VPWR _30040_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34916_ _35300_/CLK _34916_/D VGND VGND VPWR VPWR _34916_/Q sky130_fd_sc_hd__dfxtp_1
X_22930_ _22929_/X _32030_/Q _22939_/S VGND VGND VPWR VPWR _22931_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35896_ _36024_/CLK _35896_/D VGND VGND VPWR VPWR _35896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22861_ _20577_/X _22859_/X _22860_/X _20587_/X VGND VGND VPWR VPWR _22861_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34847_ _35039_/CLK _34847_/D VGND VGND VPWR VPWR _34847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24600_ _22904_/X _32790_/Q _24602_/S VGND VGND VPWR VPWR _24601_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21812_ _33006_/Q _32942_/Q _32878_/Q _32814_/Q _21589_/X _21590_/X VGND VGND VPWR
+ VPWR _21812_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25580_ _25580_/A VGND VGND VPWR VPWR _33220_/D sky130_fd_sc_hd__clkbuf_1
X_22792_ _32779_/Q _32715_/Q _32651_/Q _36107_/Q _22578_/X _21473_/A VGND VGND VPWR
+ VPWR _22792_/X sky130_fd_sc_hd__mux4_1
X_34778_ _35226_/CLK _34778_/D VGND VGND VPWR VPWR _34778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24531_ _24531_/A VGND VGND VPWR VPWR _32758_/D sky130_fd_sc_hd__clkbuf_1
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33729_ _33729_/CLK _33729_/D VGND VGND VPWR VPWR _33729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21743_ _21594_/X _21739_/X _21742_/X _21597_/X VGND VGND VPWR VPWR _21743_/X sky130_fd_sc_hd__a22o_1
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27250_ _26959_/X _33978_/Q _27260_/S VGND VGND VPWR VPWR _27251_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24462_ _22904_/X _32726_/Q _24464_/S VGND VGND VPWR VPWR _24463_/A sky130_fd_sc_hd__mux2_1
X_21674_ _22531_/A VGND VGND VPWR VPWR _21674_/X sky130_fd_sc_hd__buf_6
XFILLER_200_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26201_ _26201_/A VGND VGND VPWR VPWR _33512_/D sky130_fd_sc_hd__clkbuf_1
X_23413_ _32265_/Q _23333_/X _23413_/S VGND VGND VPWR VPWR _23414_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20625_ _22369_/A VGND VGND VPWR VPWR _22508_/A sky130_fd_sc_hd__buf_12
XFILLER_149_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27181_ _26857_/X _33945_/Q _27197_/S VGND VGND VPWR VPWR _27182_/A sky130_fd_sc_hd__mux2_1
X_24393_ _24393_/A VGND VGND VPWR VPWR _32701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26132_ _25171_/X _33480_/Q _26134_/S VGND VGND VPWR VPWR _26133_/A sky130_fd_sc_hd__mux2_1
X_23344_ _23344_/A VGND VGND VPWR VPWR _32232_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20556_ _33037_/Q _32973_/Q _32909_/Q _32845_/Q _18280_/X _18283_/X VGND VGND VPWR
+ VPWR _20556_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26063_ _25069_/X _33447_/Q _26071_/S VGND VGND VPWR VPWR _26064_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_307_CLK clkbuf_6_48__f_CLK/X VGND VGND VPWR VPWR _35577_/CLK sky130_fd_sc_hd__clkbuf_16
X_23275_ _32209_/Q _23274_/X _23301_/S VGND VGND VPWR VPWR _23276_/A sky130_fd_sc_hd__mux2_1
X_20487_ _20201_/X _20485_/X _20486_/X _20206_/X VGND VGND VPWR VPWR _20487_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25014_ _25013_/X _32981_/Q _25020_/S VGND VGND VPWR VPWR _25015_/A sky130_fd_sc_hd__mux2_1
X_22226_ _32762_/Q _32698_/Q _32634_/Q _36090_/Q _22225_/X _22009_/X VGND VGND VPWR
+ VPWR _22226_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29822_ _35165_/Q _29098_/X _29830_/S VGND VGND VPWR VPWR _29823_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22157_ _34040_/Q _33976_/Q _33912_/Q _32248_/Q _21973_/X _21974_/X VGND VGND VPWR
+ VPWR _22157_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21108_ _21104_/X _21107_/X _21030_/X _21031_/X VGND VGND VPWR VPWR _21125_/B sky130_fd_sc_hd__o211a_1
XTAP_6868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29753_ _29753_/A VGND VGND VPWR VPWR _35132_/D sky130_fd_sc_hd__clkbuf_1
X_26965_ input41/X VGND VGND VPWR VPWR _26965_/X sky130_fd_sc_hd__clkbuf_4
X_22088_ _22016_/X _22086_/X _22087_/X _22020_/X VGND VGND VPWR VPWR _22088_/X sky130_fd_sc_hd__a22o_1
XFILLER_247_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28704_ _28704_/A VGND VGND VPWR VPWR _34666_/D sky130_fd_sc_hd__clkbuf_1
X_25916_ _25916_/A VGND VGND VPWR VPWR _33377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21039_ _33176_/Q _32536_/Q _35928_/Q _35864_/Q _20968_/X _20969_/X VGND VGND VPWR
+ VPWR _21039_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26896_ _26896_/A VGND VGND VPWR VPWR _33829_/D sky130_fd_sc_hd__clkbuf_1
X_29684_ _29684_/A VGND VGND VPWR VPWR _35099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28635_ _27008_/X _34634_/Q _28641_/S VGND VGND VPWR VPWR _28636_/A sky130_fd_sc_hd__mux2_1
X_25847_ _25847_/A VGND VGND VPWR VPWR _33344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16580_ _16293_/X _16578_/X _16579_/X _16296_/X VGND VGND VPWR VPWR _16580_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28566_ _26906_/X _34601_/Q _28570_/S VGND VGND VPWR VPWR _28567_/A sky130_fd_sc_hd__mux2_1
X_25778_ _25047_/X _33312_/Q _25780_/S VGND VGND VPWR VPWR _25779_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_810 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24729_ _22892_/X _32850_/Q _24739_/S VGND VGND VPWR VPWR _24730_/A sky130_fd_sc_hd__mux2_1
X_27517_ _27517_/A VGND VGND VPWR VPWR _34104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28497_ _28497_/A VGND VGND VPWR VPWR _34568_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18250_ _16026_/X _18248_/X _18249_/X _16037_/X VGND VGND VPWR VPWR _18250_/X sky130_fd_sc_hd__a22o_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27448_ _27559_/S VGND VGND VPWR VPWR _27467_/S sky130_fd_sc_hd__clkbuf_8
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17195_/X _17198_/X _17199_/X _17200_/X VGND VGND VPWR VPWR _17201_/X sky130_fd_sc_hd__a22o_1
XFILLER_141_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18181_ _16056_/X _18179_/X _18180_/X _16068_/X VGND VGND VPWR VPWR _18181_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27379_ _34039_/Q _24373_/X _27395_/S VGND VGND VPWR VPWR _27380_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17132_ _17055_/X _17130_/X _17131_/X _17061_/X VGND VGND VPWR VPWR _17132_/X sky130_fd_sc_hd__a22o_1
XFILLER_156_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29118_ _34851_/Q _29117_/X _29142_/S VGND VGND VPWR VPWR _29119_/A sky130_fd_sc_hd__mux2_1
X_30390_ _23231_/X _35434_/Q _30392_/S VGND VGND VPWR VPWR _30391_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29049_ _30329_/A _29049_/B _30329_/B VGND VGND VPWR VPWR _29050_/A sky130_fd_sc_hd__or3b_1
X_17063_ _17908_/A VGND VGND VPWR VPWR _17063_/X sky130_fd_sc_hd__buf_4
XFILLER_195_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16014_ _17901_/A VGND VGND VPWR VPWR _16014_/X sky130_fd_sc_hd__buf_2
XFILLER_6_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32060_ _36028_/CLK _32060_/D VGND VGND VPWR VPWR _32060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31011_ _35728_/Q _29058_/X _31025_/S VGND VGND VPWR VPWR _31012_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_1243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17965_ _34563_/Q _32451_/Q _34435_/Q _34371_/Q _17931_/X _17932_/X VGND VGND VPWR
+ VPWR _17965_/X sky130_fd_sc_hd__mux4_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19704_ _33524_/Q _33460_/Q _33396_/Q _33332_/Q _19423_/X _19424_/X VGND VGND VPWR
+ VPWR _19704_/X sky130_fd_sc_hd__mux4_1
X_35750_ _35750_/CLK _35750_/D VGND VGND VPWR VPWR _35750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16916_ _34022_/Q _33958_/Q _33894_/Q _32193_/Q _16667_/X _16668_/X VGND VGND VPWR
+ VPWR _16916_/X sky130_fd_sc_hd__mux4_1
X_32962_ _32962_/CLK _32962_/D VGND VGND VPWR VPWR _32962_/Q sky130_fd_sc_hd__dfxtp_1
X_17896_ _35073_/Q _35009_/Q _34945_/Q _34881_/Q _17862_/X _17863_/X VGND VGND VPWR
+ VPWR _17896_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34701_ _35341_/CLK _34701_/D VGND VGND VPWR VPWR _34701_/Q sky130_fd_sc_hd__dfxtp_1
X_31913_ _23289_/X _36156_/Q _31919_/S VGND VGND VPWR VPWR _31914_/A sky130_fd_sc_hd__mux2_1
X_19635_ _34034_/Q _33970_/Q _33906_/Q _32242_/Q _19320_/X _19321_/X VGND VGND VPWR
+ VPWR _19635_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35681_ _35807_/CLK _35681_/D VGND VGND VPWR VPWR _35681_/Q sky130_fd_sc_hd__dfxtp_1
X_16847_ _17906_/A VGND VGND VPWR VPWR _16847_/X sky130_fd_sc_hd__clkbuf_4
X_32893_ _36031_/CLK _32893_/D VGND VGND VPWR VPWR _32893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34632_ _35337_/CLK _34632_/D VGND VGND VPWR VPWR _34632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31844_ _23127_/X _36123_/Q _31856_/S VGND VGND VPWR VPWR _31845_/A sky130_fd_sc_hd__mux2_1
X_19566_ _34288_/Q _34224_/Q _34160_/Q _34096_/Q _19389_/X _19390_/X VGND VGND VPWR
+ VPWR _19566_/X sky130_fd_sc_hd__mux4_1
XFILLER_213_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16778_ _33250_/Q _36130_/Q _33122_/Q _33058_/Q _16705_/X _16706_/X VGND VGND VPWR
+ VPWR _16778_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18517_ _20282_/A VGND VGND VPWR VPWR _18517_/X sky130_fd_sc_hd__buf_6
XFILLER_0_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34563_ _35331_/CLK _34563_/D VGND VGND VPWR VPWR _34563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31775_ _31775_/A VGND VGND VPWR VPWR _36090_/D sky130_fd_sc_hd__clkbuf_1
X_19497_ _20203_/A VGND VGND VPWR VPWR _19497_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33514_ _35386_/CLK _33514_/D VGND VGND VPWR VPWR _33514_/Q sky130_fd_sc_hd__dfxtp_1
X_18448_ _18442_/X _18447_/X _18311_/X VGND VGND VPWR VPWR _18472_/A sky130_fd_sc_hd__o21ba_1
X_30726_ _30726_/A VGND VGND VPWR VPWR _35593_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34494_ _35837_/CLK _34494_/D VGND VGND VPWR VPWR _34494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36233_ _36237_/CLK _36233_/D VGND VGND VPWR VPWR _36233_/Q sky130_fd_sc_hd__dfxtp_1
X_33445_ _35991_/CLK _33445_/D VGND VGND VPWR VPWR _33445_/Q sky130_fd_sc_hd__dfxtp_1
X_18379_ _20012_/A VGND VGND VPWR VPWR _18379_/X sky130_fd_sc_hd__buf_6
XFILLER_147_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30657_ _30657_/A VGND VGND VPWR VPWR _35560_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_93_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _36202_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_239_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20410_ _35784_/Q _35144_/Q _34504_/Q _33864_/Q _20146_/X _20147_/X VGND VGND VPWR
+ VPWR _20410_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36164_ _36166_/CLK _36164_/D VGND VGND VPWR VPWR _36164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21390_ _21241_/X _21386_/X _21389_/X _21244_/X VGND VGND VPWR VPWR _21390_/X sky130_fd_sc_hd__a22o_1
X_30588_ _23330_/X _35528_/Q _30590_/S VGND VGND VPWR VPWR _30589_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33376_ _34017_/CLK _33376_/D VGND VGND VPWR VPWR _33376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35115_ _35945_/CLK _35115_/D VGND VGND VPWR VPWR _35115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32327_ _35339_/CLK _32327_/D VGND VGND VPWR VPWR _32327_/Q sky130_fd_sc_hd__dfxtp_1
X_20341_ _20337_/X _20340_/X _20134_/X VGND VGND VPWR VPWR _20363_/A sky130_fd_sc_hd__o21ba_2
XFILLER_88_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36095_ _36095_/CLK _36095_/D VGND VGND VPWR VPWR _36095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20272_ _34308_/Q _34244_/Q _34180_/Q _34116_/Q _20095_/X _20096_/X VGND VGND VPWR
+ VPWR _20272_/X sky130_fd_sc_hd__mux4_1
X_23060_ _23059_/X _32072_/Q _23063_/S VGND VGND VPWR VPWR _23061_/A sky130_fd_sc_hd__mux2_1
X_35046_ _35942_/CLK _35046_/D VGND VGND VPWR VPWR _35046_/Q sky130_fd_sc_hd__dfxtp_1
X_32258_ _33922_/CLK _32258_/D VGND VGND VPWR VPWR _32258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22011_ _22582_/A VGND VGND VPWR VPWR _22011_/X sky130_fd_sc_hd__buf_4
XTAP_6109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31209_ _35822_/Q input26/X _31223_/S VGND VGND VPWR VPWR _31210_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32189_ _35749_/CLK _32189_/D VGND VGND VPWR VPWR _32189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26750_ _26819_/S VGND VGND VPWR VPWR _26769_/S sky130_fd_sc_hd__buf_6
XFILLER_233_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23962_ _23062_/X _32521_/Q _23962_/S VGND VGND VPWR VPWR _23963_/A sky130_fd_sc_hd__mux2_1
XTAP_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35948_ _35949_/CLK _35948_/D VGND VGND VPWR VPWR _35948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25701_ _25701_/A VGND VGND VPWR VPWR _33276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22913_ _22913_/A VGND VGND VPWR VPWR _32024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26681_ _25183_/X _33740_/Q _26683_/S VGND VGND VPWR VPWR _26682_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_867 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35879_ _35879_/CLK _35879_/D VGND VGND VPWR VPWR _35879_/Q sky130_fd_sc_hd__dfxtp_1
X_23893_ _22960_/X _32488_/Q _23899_/S VGND VGND VPWR VPWR _23894_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25632_ _25632_/A VGND VGND VPWR VPWR _33243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28420_ _28420_/A VGND VGND VPWR VPWR _34531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22844_ _22844_/A VGND VGND VPWR VPWR _36236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28351_ _34499_/Q _24410_/X _28363_/S VGND VGND VPWR VPWR _28352_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25563_ _25563_/A VGND VGND VPWR VPWR _33212_/D sky130_fd_sc_hd__clkbuf_1
X_22775_ _22771_/X _22774_/X _22453_/A VGND VGND VPWR VPWR _22783_/C sky130_fd_sc_hd__o21ba_1
XFILLER_52_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27302_ _27302_/A VGND VGND VPWR VPWR _34002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24514_ _24514_/A VGND VGND VPWR VPWR _32750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28282_ _34466_/Q _24307_/X _28300_/S VGND VGND VPWR VPWR _28283_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21726_ _34028_/Q _33964_/Q _33900_/Q _32236_/Q _21620_/X _21621_/X VGND VGND VPWR
+ VPWR _21726_/X sky130_fd_sc_hd__mux4_1
XFILLER_227_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25494_ _25494_/A VGND VGND VPWR VPWR _33179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27233_ _26934_/X _33970_/Q _27239_/S VGND VGND VPWR VPWR _27234_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24445_ _24577_/S VGND VGND VPWR VPWR _24464_/S sky130_fd_sc_hd__clkbuf_4
X_21657_ _32746_/Q _32682_/Q _32618_/Q _36074_/Q _21519_/X _21656_/X VGND VGND VPWR
+ VPWR _21657_/X sky130_fd_sc_hd__mux4_1
XFILLER_240_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_84_CLK clkbuf_leaf_87_CLK/A VGND VGND VPWR VPWR _35863_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27164_ _26832_/X _33937_/Q _27176_/S VGND VGND VPWR VPWR _27165_/A sky130_fd_sc_hd__mux2_1
X_20608_ _33998_/Q _33934_/Q _33870_/Q _32142_/Q _20605_/X _20607_/X VGND VGND VPWR
+ VPWR _20608_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24376_ input37/X VGND VGND VPWR VPWR _24376_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_149_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21588_ _32488_/Q _32360_/Q _32040_/Q _36008_/Q _21523_/X _21311_/X VGND VGND VPWR
+ VPWR _21588_/X sky130_fd_sc_hd__mux4_1
X_26115_ _26142_/S VGND VGND VPWR VPWR _26134_/S sky130_fd_sc_hd__buf_4
X_23327_ input53/X VGND VGND VPWR VPWR _23327_/X sky130_fd_sc_hd__buf_4
XFILLER_10_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20539_ _34572_/Q _32460_/Q _34444_/Q _34380_/Q _18363_/X _18365_/X VGND VGND VPWR
+ VPWR _20539_/X sky130_fd_sc_hd__mux4_1
XFILLER_193_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27095_ _27095_/A VGND VGND VPWR VPWR _33904_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26046_ _25044_/X _33439_/Q _26050_/S VGND VGND VPWR VPWR _26047_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23258_ _23258_/A VGND VGND VPWR VPWR _32203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22209_ _34809_/Q _34745_/Q _34681_/Q _34617_/Q _21888_/X _21889_/X VGND VGND VPWR
+ VPWR _22209_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23189_ _32177_/Q _23124_/X _23206_/S VGND VGND VPWR VPWR _23190_/A sky130_fd_sc_hd__mux2_1
XFILLER_234_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29805_ _35157_/Q _29073_/X _29809_/S VGND VGND VPWR VPWR _29806_/A sky130_fd_sc_hd__mux2_1
XTAP_6654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27997_ _26863_/X _34331_/Q _28009_/S VGND VGND VPWR VPWR _27998_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17750_ _17507_/X _17748_/X _17749_/X _17512_/X VGND VGND VPWR VPWR _17750_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29736_ _29736_/A VGND VGND VPWR VPWR _35124_/D sky130_fd_sc_hd__clkbuf_1
X_26948_ _26946_/X _33846_/Q _26975_/S VGND VGND VPWR VPWR _26949_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16701_ _16697_/X _16700_/X _16422_/X VGND VGND VPWR VPWR _16733_/A sky130_fd_sc_hd__o21ba_1
XFILLER_247_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29667_ _29667_/A VGND VGND VPWR VPWR _35091_/D sky130_fd_sc_hd__clkbuf_1
X_17681_ _17677_/X _17680_/X _17514_/X VGND VGND VPWR VPWR _17682_/D sky130_fd_sc_hd__o21ba_1
XFILLER_43_1198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26879_ _26878_/X _33824_/Q _26882_/S VGND VGND VPWR VPWR _26880_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19420_ _33772_/Q _33708_/Q _33644_/Q _33580_/Q _19143_/X _19144_/X VGND VGND VPWR
+ VPWR _19420_/X sky130_fd_sc_hd__mux4_1
X_28618_ _28618_/A VGND VGND VPWR VPWR _34625_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16632_ _32734_/Q _32670_/Q _32606_/Q _36062_/Q _16566_/X _16350_/X VGND VGND VPWR
+ VPWR _16632_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29598_ _35059_/Q _29166_/X _29602_/S VGND VGND VPWR VPWR _29599_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19351_ _33514_/Q _33450_/Q _33386_/Q _33322_/Q _19070_/X _19071_/X VGND VGND VPWR
+ VPWR _19351_/X sky130_fd_sc_hd__mux4_1
X_28549_ _26881_/X _34593_/Q _28549_/S VGND VGND VPWR VPWR _28550_/A sky130_fd_sc_hd__mux2_1
X_16563_ _34012_/Q _33948_/Q _33884_/Q _32156_/Q _16314_/X _16315_/X VGND VGND VPWR
+ VPWR _16563_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18302_ _20073_/A VGND VGND VPWR VPWR _20211_/A sky130_fd_sc_hd__buf_12
XFILLER_245_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31560_ _31560_/A VGND VGND VPWR VPWR _35988_/D sky130_fd_sc_hd__clkbuf_1
X_19282_ _34024_/Q _33960_/Q _33896_/Q _32215_/Q _18967_/X _18968_/X VGND VGND VPWR
+ VPWR _19282_/X sky130_fd_sc_hd__mux4_1
X_16494_ _17858_/A VGND VGND VPWR VPWR _16494_/X sky130_fd_sc_hd__buf_4
XFILLER_241_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18233_ _33228_/Q _32588_/Q _35980_/Q _35916_/Q _16075_/X _16076_/X VGND VGND VPWR
+ VPWR _18233_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30511_ _23152_/X _35491_/Q _30527_/S VGND VGND VPWR VPWR _30512_/A sky130_fd_sc_hd__mux2_1
X_31491_ _23264_/X _35956_/Q _31493_/S VGND VGND VPWR VPWR _31492_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_75_CLK clkbuf_leaf_76_CLK/A VGND VGND VPWR VPWR _36114_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30442_ _30442_/A VGND VGND VPWR VPWR _35458_/D sky130_fd_sc_hd__clkbuf_1
X_33230_ _33234_/CLK _33230_/D VGND VGND VPWR VPWR _33230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18164_ _17149_/A _18162_/X _18163_/X _17152_/A VGND VGND VPWR VPWR _18164_/X sky130_fd_sc_hd__a22o_1
XFILLER_184_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17115_ _35051_/Q _34987_/Q _34923_/Q _34859_/Q _16803_/X _16804_/X VGND VGND VPWR
+ VPWR _17115_/X sky130_fd_sc_hd__mux4_1
XFILLER_102_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18095_ _33800_/Q _33736_/Q _33672_/Q _33608_/Q _17902_/X _17903_/X VGND VGND VPWR
+ VPWR _18095_/X sky130_fd_sc_hd__mux4_1
XFILLER_183_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33161_ _35585_/CLK _33161_/D VGND VGND VPWR VPWR _33161_/Q sky130_fd_sc_hd__dfxtp_1
X_30373_ _30463_/S VGND VGND VPWR VPWR _30392_/S sky130_fd_sc_hd__buf_4
XFILLER_102_1248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32112_ _35552_/CLK _32112_/D VGND VGND VPWR VPWR _32112_/Q sky130_fd_sc_hd__dfxtp_1
X_17046_ _17046_/A _17046_/B _17046_/C _17046_/D VGND VGND VPWR VPWR _17047_/A sky130_fd_sc_hd__or4_4
X_33092_ _36166_/CLK _33092_/D VGND VGND VPWR VPWR _33092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32043_ _34794_/CLK _32043_/D VGND VGND VPWR VPWR _32043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _18789_/X _18995_/X _18996_/X _18794_/X VGND VGND VPWR VPWR _18997_/X sky130_fd_sc_hd__a22o_1
XFILLER_26_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35802_ _36063_/CLK _35802_/D VGND VGND VPWR VPWR _35802_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17948_ _17761_/X _17946_/X _17947_/X _17767_/X VGND VGND VPWR VPWR _17948_/X sky130_fd_sc_hd__a22o_1
XFILLER_152_1360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33994_ _35273_/CLK _33994_/D VGND VGND VPWR VPWR _33994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35733_ _35733_/CLK _35733_/D VGND VGND VPWR VPWR _35733_/Q sky130_fd_sc_hd__dfxtp_1
X_32945_ _36081_/CLK _32945_/D VGND VGND VPWR VPWR _32945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17879_ _33281_/Q _36161_/Q _33153_/Q _33089_/Q _17764_/X _17765_/X VGND VGND VPWR
+ VPWR _17879_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_26__f_CLK clkbuf_5_13_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_66_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_93_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19618_ _35569_/Q _35505_/Q _35441_/Q _35377_/Q _19550_/X _19551_/X VGND VGND VPWR
+ VPWR _19618_/X sky130_fd_sc_hd__mux4_1
XFILLER_214_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35664_ _35664_/CLK _35664_/D VGND VGND VPWR VPWR _35664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20890_ _35732_/Q _35092_/Q _34452_/Q _33812_/Q _20649_/X _20651_/X VGND VGND VPWR
+ VPWR _20890_/X sky130_fd_sc_hd__mux4_1
X_32876_ _36080_/CLK _32876_/D VGND VGND VPWR VPWR _32876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34615_ _34745_/CLK _34615_/D VGND VGND VPWR VPWR _34615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31827_ _23102_/X _36115_/Q _31835_/S VGND VGND VPWR VPWR _31828_/A sky130_fd_sc_hd__mux2_1
X_19549_ _19294_/X _19547_/X _19548_/X _19297_/X VGND VGND VPWR VPWR _19549_/X sky130_fd_sc_hd__a22o_1
X_35595_ _35851_/CLK _35595_/D VGND VGND VPWR VPWR _35595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22560_ _22305_/X _22558_/X _22559_/X _22308_/X VGND VGND VPWR VPWR _22560_/X sky130_fd_sc_hd__a22o_1
X_34546_ _34997_/CLK _34546_/D VGND VGND VPWR VPWR _34546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31758_ _31758_/A VGND VGND VPWR VPWR _36082_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21511_ _21511_/A VGND VGND VPWR VPWR _36197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30709_ _35585_/Q _29210_/X _30725_/S VGND VGND VPWR VPWR _30710_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22491_ _22487_/X _22490_/X _22453_/X VGND VGND VPWR VPWR _22499_/C sky130_fd_sc_hd__o21ba_1
X_34477_ _35564_/CLK _34477_/D VGND VGND VPWR VPWR _34477_/Q sky130_fd_sc_hd__dfxtp_1
X_31689_ _31689_/A VGND VGND VPWR VPWR _36049_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_66_CLK clkbuf_leaf_66_CLK/A VGND VGND VPWR VPWR _36052_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24230_ _23056_/X _32647_/Q _24234_/S VGND VGND VPWR VPWR _24231_/A sky130_fd_sc_hd__mux2_1
X_36216_ _36216_/CLK _36216_/D VGND VGND VPWR VPWR _36216_/Q sky130_fd_sc_hd__dfxtp_1
X_33428_ _36237_/CLK _33428_/D VGND VGND VPWR VPWR _33428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21442_ _22501_/A VGND VGND VPWR VPWR _21442_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_222_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36147_ _36147_/CLK _36147_/D VGND VGND VPWR VPWR _36147_/Q sky130_fd_sc_hd__dfxtp_1
X_24161_ _22954_/X _32614_/Q _24171_/S VGND VGND VPWR VPWR _24162_/A sky130_fd_sc_hd__mux2_1
X_33359_ _33490_/CLK _33359_/D VGND VGND VPWR VPWR _33359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21373_ _34018_/Q _33954_/Q _33890_/Q _32162_/Q _21267_/X _21268_/X VGND VGND VPWR
+ VPWR _21373_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23112_ _32150_/Q _23111_/X _23115_/S VGND VGND VPWR VPWR _23113_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20324_ _20005_/X _20322_/X _20323_/X _20008_/X VGND VGND VPWR VPWR _20324_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24092_ _23053_/X _32582_/Q _24098_/S VGND VGND VPWR VPWR _24093_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36078_ _36078_/CLK _36078_/D VGND VGND VPWR VPWR _36078_/Q sky130_fd_sc_hd__dfxtp_1
X_23043_ _23043_/A VGND VGND VPWR VPWR _32066_/D sky130_fd_sc_hd__clkbuf_1
X_35029_ _36196_/CLK _35029_/D VGND VGND VPWR VPWR _35029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27920_ _27920_/A VGND VGND VPWR VPWR _34294_/D sky130_fd_sc_hd__clkbuf_1
X_20255_ _20000_/X _20253_/X _20254_/X _20003_/X VGND VGND VPWR VPWR _20255_/X sky130_fd_sc_hd__a22o_1
XFILLER_235_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27851_ _34262_/Q _24270_/X _27853_/S VGND VGND VPWR VPWR _27852_/A sky130_fd_sc_hd__mux2_1
X_20186_ _35777_/Q _35137_/Q _34497_/Q _33857_/Q _20146_/X _20147_/X VGND VGND VPWR
+ VPWR _20186_/X sky130_fd_sc_hd__mux4_1
XTAP_5205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26802_ _26802_/A VGND VGND VPWR VPWR _33796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24994_ _24994_/A VGND VGND VPWR VPWR _32974_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27782_ _27782_/A VGND VGND VPWR VPWR _34229_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29521_ _35022_/Q _29048_/X _29539_/S VGND VGND VPWR VPWR _29522_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23945_ _23945_/A VGND VGND VPWR VPWR _32512_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26733_ _26733_/A VGND VGND VPWR VPWR _33763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26664_ _26664_/A VGND VGND VPWR VPWR _33731_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29452_ _29452_/A VGND VGND VPWR VPWR _34989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_803 _22892_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23876_ _22935_/X _32480_/Q _23878_/S VGND VGND VPWR VPWR _23877_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_814 _22920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_825 _23105_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25615_ _25615_/A VGND VGND VPWR VPWR _33235_/D sky130_fd_sc_hd__clkbuf_1
X_28403_ _28403_/A VGND VGND VPWR VPWR _34523_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_836 _23270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22827_ _21754_/A _22825_/X _22826_/X _21759_/A VGND VGND VPWR VPWR _22827_/X sky130_fd_sc_hd__a22o_1
X_29383_ _29383_/A VGND VGND VPWR VPWR _34957_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_847 _23970_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26595_ _26595_/A VGND VGND VPWR VPWR _33698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_858 _24348_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_869 _24577_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28334_ _34491_/Q _24385_/X _28342_/S VGND VGND VPWR VPWR _28335_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25546_ _25546_/A VGND VGND VPWR VPWR _33204_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22758_ _33546_/Q _33482_/Q _33418_/Q _33354_/Q _20633_/X _20635_/X VGND VGND VPWR
+ VPWR _22758_/X sky130_fd_sc_hd__mux4_2
XFILLER_71_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21709_ _21599_/X _21707_/X _21708_/X _21602_/X VGND VGND VPWR VPWR _21709_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28265_ _34458_/Q _24283_/X _28279_/S VGND VGND VPWR VPWR _28266_/A sky130_fd_sc_hd__mux2_1
X_25477_ _25477_/A VGND VGND VPWR VPWR _33171_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22689_ _34567_/Q _32455_/Q _34439_/Q _34375_/Q _22531_/X _22532_/X VGND VGND VPWR
+ VPWR _22689_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_57_CLK clkbuf_leaf_57_CLK/A VGND VGND VPWR VPWR _35992_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_240_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24428_ input55/X VGND VGND VPWR VPWR _24428_/X sky130_fd_sc_hd__buf_6
X_27216_ _26909_/X _33962_/Q _27218_/S VGND VGND VPWR VPWR _27217_/A sky130_fd_sc_hd__mux2_1
X_28196_ _28196_/A VGND VGND VPWR VPWR _34425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27147_ _27147_/A VGND VGND VPWR VPWR _33929_/D sky130_fd_sc_hd__clkbuf_1
X_24359_ _24359_/A VGND VGND VPWR VPWR _32690_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27078_ _27078_/A VGND VGND VPWR VPWR _33896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26029_ _25019_/X _33431_/Q _26029_/S VGND VGND VPWR VPWR _26030_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18920_ _35037_/Q _34973_/Q _34909_/Q _34845_/Q _18750_/X _18751_/X VGND VGND VPWR
+ VPWR _18920_/X sky130_fd_sc_hd__mux4_1
XTAP_7130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1202 _23102_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1213 _23327_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18851_ _35291_/Q _35227_/Q _35163_/Q _32283_/Q _18600_/X _18601_/X VGND VGND VPWR
+ VPWR _18851_/X sky130_fd_sc_hd__mux4_1
XTAP_6440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1224 _24342_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1235 _24852_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1246 _26412_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17802_ _17798_/X _17801_/X _17481_/X VGND VGND VPWR VPWR _17824_/A sky130_fd_sc_hd__o21ba_1
XFILLER_132_1219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1257 _27509_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1268 _30192_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18782_ _18743_/X _18780_/X _18781_/X _18746_/X VGND VGND VPWR VPWR _18782_/X sky130_fd_sc_hd__a22o_1
XFILLER_227_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15994_ input67/X input68/X VGND VGND VPWR VPWR _15995_/A sky130_fd_sc_hd__and2_1
XANTENNA_1279 _17911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17733_ _17408_/X _17731_/X _17732_/X _17414_/X VGND VGND VPWR VPWR _17733_/X sky130_fd_sc_hd__a22o_1
X_29719_ _35116_/Q _29144_/X _29737_/S VGND VGND VPWR VPWR _29720_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30991_ _35719_/Q _29228_/X _30995_/S VGND VGND VPWR VPWR _30992_/A sky130_fd_sc_hd__mux2_1
XTAP_5794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32730_ _36121_/CLK _32730_/D VGND VGND VPWR VPWR _32730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17664_ _17416_/X _17662_/X _17663_/X _17420_/X VGND VGND VPWR VPWR _17664_/X sky130_fd_sc_hd__a22o_1
XFILLER_247_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19403_ _19399_/X _19402_/X _19083_/X _19084_/X VGND VGND VPWR VPWR _19418_/B sky130_fd_sc_hd__o211a_1
XFILLER_223_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16615_ _16611_/X _16614_/X _16441_/X VGND VGND VPWR VPWR _16623_/C sky130_fd_sc_hd__o21ba_1
X_32661_ _36116_/CLK _32661_/D VGND VGND VPWR VPWR _32661_/Q sky130_fd_sc_hd__dfxtp_1
X_17595_ _17408_/X _17593_/X _17594_/X _17414_/X VGND VGND VPWR VPWR _17595_/X sky130_fd_sc_hd__a22o_1
X_34400_ _35039_/CLK _34400_/D VGND VGND VPWR VPWR _34400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19334_ _19294_/X _19332_/X _19333_/X _19297_/X VGND VGND VPWR VPWR _19334_/X sky130_fd_sc_hd__a22o_1
X_31612_ _36013_/Q input25/X _31628_/S VGND VGND VPWR VPWR _31613_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16546_ _35547_/Q _35483_/Q _35419_/Q _35355_/Q _16544_/X _16545_/X VGND VGND VPWR
+ VPWR _16546_/X sky130_fd_sc_hd__mux4_1
X_35380_ _35700_/CLK _35380_/D VGND VGND VPWR VPWR _35380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32592_ _36048_/CLK _32592_/D VGND VGND VPWR VPWR _32592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34331_ _34970_/CLK _34331_/D VGND VGND VPWR VPWR _34331_/Q sky130_fd_sc_hd__dfxtp_1
X_31543_ _23345_/X _35981_/Q _31543_/S VGND VGND VPWR VPWR _31544_/A sky130_fd_sc_hd__mux2_1
X_19265_ _35559_/Q _35495_/Q _35431_/Q _35367_/Q _19197_/X _19198_/X VGND VGND VPWR
+ VPWR _19265_/X sky130_fd_sc_hd__mux4_1
X_16477_ _33177_/Q _32537_/Q _35929_/Q _35865_/Q _16368_/X _16369_/X VGND VGND VPWR
+ VPWR _16477_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_48_CLK clkbuf_leaf_50_CLK/A VGND VGND VPWR VPWR _36129_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_176_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18216_ _34316_/Q _34252_/Q _34188_/Q _34124_/Q _16045_/X _16046_/X VGND VGND VPWR
+ VPWR _18216_/X sky130_fd_sc_hd__mux4_1
X_34262_ _34262_/CLK _34262_/D VGND VGND VPWR VPWR _34262_/Q sky130_fd_sc_hd__dfxtp_1
X_19196_ _18941_/X _19194_/X _19195_/X _18944_/X VGND VGND VPWR VPWR _19196_/X sky130_fd_sc_hd__a22o_1
X_31474_ _31543_/S VGND VGND VPWR VPWR _31493_/S sky130_fd_sc_hd__buf_6
X_36001_ _36001_/CLK _36001_/D VGND VGND VPWR VPWR _36001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33213_ _35965_/CLK _33213_/D VGND VGND VPWR VPWR _33213_/Q sky130_fd_sc_hd__dfxtp_1
X_18147_ _35337_/Q _35273_/Q _35209_/Q _32329_/Q _16088_/X _16090_/X VGND VGND VPWR
+ VPWR _18147_/X sky130_fd_sc_hd__mux4_1
X_30425_ _30425_/A VGND VGND VPWR VPWR _35450_/D sky130_fd_sc_hd__clkbuf_1
X_34193_ _34262_/CLK _34193_/D VGND VGND VPWR VPWR _34193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33144_ _36088_/CLK _33144_/D VGND VGND VPWR VPWR _33144_/Q sky130_fd_sc_hd__dfxtp_1
X_18078_ _18074_/X _18077_/X _17842_/X _17843_/X VGND VGND VPWR VPWR _18093_/B sky130_fd_sc_hd__o211a_1
XFILLER_172_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30356_ _30356_/A VGND VGND VPWR VPWR _35417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17029_ _33001_/Q _32937_/Q _32873_/Q _32809_/Q _16989_/X _16990_/X VGND VGND VPWR
+ VPWR _17029_/X sky130_fd_sc_hd__mux4_1
X_30287_ _30287_/A VGND VGND VPWR VPWR _35385_/D sky130_fd_sc_hd__clkbuf_1
X_33075_ _34033_/CLK _33075_/D VGND VGND VPWR VPWR _33075_/Q sky130_fd_sc_hd__dfxtp_1
X_20040_ _20000_/X _20038_/X _20039_/X _20003_/X VGND VGND VPWR VPWR _20040_/X sky130_fd_sc_hd__a22o_1
XFILLER_217_1154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32026_ _35994_/CLK _32026_/D VGND VGND VPWR VPWR _32026_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33977_ _36154_/CLK _33977_/D VGND VGND VPWR VPWR _33977_/Q sky130_fd_sc_hd__dfxtp_1
X_21991_ _21987_/X _21990_/X _21747_/X VGND VGND VPWR VPWR _21999_/C sky130_fd_sc_hd__o21ba_1
XFILLER_66_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35716_ _35843_/CLK _35716_/D VGND VGND VPWR VPWR _35716_/Q sky130_fd_sc_hd__dfxtp_1
X_23730_ _22920_/X _32411_/Q _23742_/S VGND VGND VPWR VPWR _23731_/A sky130_fd_sc_hd__mux2_1
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20942_ _33750_/Q _33686_/Q _33622_/Q _33558_/Q _20737_/X _20738_/X VGND VGND VPWR
+ VPWR _20942_/X sky130_fd_sc_hd__mux4_1
X_32928_ _36001_/CLK _32928_/D VGND VGND VPWR VPWR _32928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35647_ _35710_/CLK _35647_/D VGND VGND VPWR VPWR _35647_/Q sky130_fd_sc_hd__dfxtp_1
X_23661_ _32380_/Q _23289_/X _23667_/S VGND VGND VPWR VPWR _23662_/A sky130_fd_sc_hd__mux2_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20873_ _34260_/Q _34196_/Q _34132_/Q _34068_/Q _20605_/X _20607_/X VGND VGND VPWR
+ VPWR _20873_/X sky130_fd_sc_hd__mux4_1
X_32859_ _35995_/CLK _32859_/D VGND VGND VPWR VPWR _32859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25400_ _25100_/X _33137_/Q _25408_/S VGND VGND VPWR VPWR _25401_/A sky130_fd_sc_hd__mux2_1
X_22612_ _32773_/Q _32709_/Q _32645_/Q _36101_/Q _22578_/X _22362_/X VGND VGND VPWR
+ VPWR _22612_/X sky130_fd_sc_hd__mux4_1
X_26380_ _26380_/A VGND VGND VPWR VPWR _33597_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35578_ _35578_/CLK _35578_/D VGND VGND VPWR VPWR _35578_/Q sky130_fd_sc_hd__dfxtp_1
X_23592_ _32347_/Q _23127_/X _23604_/S VGND VGND VPWR VPWR _23593_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25331_ _24998_/X _33104_/Q _25345_/S VGND VGND VPWR VPWR _25332_/A sky130_fd_sc_hd__mux2_1
X_22543_ _34051_/Q _33987_/Q _33923_/Q _32259_/Q _22326_/X _22327_/X VGND VGND VPWR
+ VPWR _22543_/X sky130_fd_sc_hd__mux4_1
X_34529_ _35807_/CLK _34529_/D VGND VGND VPWR VPWR _34529_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_39_CLK clkbuf_6_7__f_CLK/X VGND VGND VPWR VPWR _32666_/CLK sky130_fd_sc_hd__clkbuf_16
X_28050_ _28050_/A VGND VGND VPWR VPWR _34356_/D sky130_fd_sc_hd__clkbuf_1
X_25262_ _25097_/X _33072_/Q _25272_/S VGND VGND VPWR VPWR _25263_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22474_ _33537_/Q _33473_/Q _33409_/Q _33345_/Q _22429_/X _22430_/X VGND VGND VPWR
+ VPWR _22474_/X sky130_fd_sc_hd__mux4_1
X_27001_ _27001_/A VGND VGND VPWR VPWR _33863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24213_ _23031_/X _32639_/Q _24213_/S VGND VGND VPWR VPWR _24214_/A sky130_fd_sc_hd__mux2_1
X_21425_ _21421_/X _21424_/X _21383_/X _21384_/X VGND VGND VPWR VPWR _21440_/B sky130_fd_sc_hd__o211a_1
XFILLER_194_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25193_ _24995_/X _33039_/Q _25209_/S VGND VGND VPWR VPWR _25194_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24144_ _22929_/X _32606_/Q _24150_/S VGND VGND VPWR VPWR _24145_/A sky130_fd_sc_hd__mux2_1
X_21356_ _21246_/X _21354_/X _21355_/X _21249_/X VGND VGND VPWR VPWR _21356_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20307_ _20201_/X _20305_/X _20306_/X _20206_/X VGND VGND VPWR VPWR _20307_/X sky130_fd_sc_hd__a22o_1
XFILLER_150_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24075_ _23028_/X _32574_/Q _24077_/S VGND VGND VPWR VPWR _24076_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28952_ _34784_/Q _24301_/X _28954_/S VGND VGND VPWR VPWR _28953_/A sky130_fd_sc_hd__mux2_1
X_21287_ _35295_/Q _35231_/Q _35167_/Q _32287_/Q _21253_/X _21254_/X VGND VGND VPWR
+ VPWR _21287_/X sky130_fd_sc_hd__mux4_1
X_23026_ _23025_/X _32061_/Q _23032_/S VGND VGND VPWR VPWR _23027_/A sky130_fd_sc_hd__mux2_1
X_27903_ _27903_/A VGND VGND VPWR VPWR _34286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20238_ _20238_/A VGND VGND VPWR VPWR _32130_/D sky130_fd_sc_hd__clkbuf_4
XTAP_5002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28883_ _28883_/A VGND VGND VPWR VPWR _34751_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27834_ _27966_/S VGND VGND VPWR VPWR _27853_/S sky130_fd_sc_hd__buf_4
XTAP_5035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20169_ _20169_/A _20169_/B _20169_/C _20169_/D VGND VGND VPWR VPWR _20170_/A sky130_fd_sc_hd__or4_2
XTAP_5046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27765_ _34221_/Q _24342_/X _27781_/S VGND VGND VPWR VPWR _27766_/A sky130_fd_sc_hd__mux2_1
X_24977_ _23059_/X _32968_/Q _24979_/S VGND VGND VPWR VPWR _24978_/A sky130_fd_sc_hd__mux2_1
XTAP_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29504_ _29504_/A VGND VGND VPWR VPWR _35014_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26716_ _26716_/A VGND VGND VPWR VPWR _33755_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23928_ _23928_/A VGND VGND VPWR VPWR _32504_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27696_ _34189_/Q _24440_/X _27696_/S VGND VGND VPWR VPWR _27697_/A sky130_fd_sc_hd__mux2_1
XTAP_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_600 _20167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_611 _18505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_622 _18609_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29435_ _29435_/A VGND VGND VPWR VPWR _34981_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26647_ _26647_/A VGND VGND VPWR VPWR _33723_/D sky130_fd_sc_hd__clkbuf_1
X_23859_ _23970_/S VGND VGND VPWR VPWR _23878_/S sky130_fd_sc_hd__buf_4
XANTENNA_633 _18993_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_644 _19390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_655 _20333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_919 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_666 _22396_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16400_ _16288_/X _16398_/X _16399_/X _16291_/X VGND VGND VPWR VPWR _16400_/X sky130_fd_sc_hd__a22o_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29366_ _23319_/X _34949_/Q _29374_/S VGND VGND VPWR VPWR _29367_/A sky130_fd_sc_hd__mux2_1
XANTENNA_677 _22556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17380_ _17055_/X _17378_/X _17379_/X _17061_/X VGND VGND VPWR VPWR _17380_/X sky130_fd_sc_hd__a22o_1
XFILLER_60_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_688 _22442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26578_ _26578_/A VGND VGND VPWR VPWR _33690_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_699 _22458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16331_ _16293_/X _16329_/X _16330_/X _16296_/X VGND VGND VPWR VPWR _16331_/X sky130_fd_sc_hd__a22o_1
X_28317_ _34483_/Q _24360_/X _28321_/S VGND VGND VPWR VPWR _28318_/A sky130_fd_sc_hd__mux2_1
X_25529_ _33196_/Q _24338_/X _25547_/S VGND VGND VPWR VPWR _25530_/A sky130_fd_sc_hd__mux2_1
X_29297_ _23175_/X _34916_/Q _29311_/S VGND VGND VPWR VPWR _29298_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16262_ _16258_/X _16261_/X _16071_/X VGND VGND VPWR VPWR _16270_/C sky130_fd_sc_hd__o21ba_1
X_19050_ _19046_/X _19049_/X _18730_/X _18731_/X VGND VGND VPWR VPWR _19065_/B sky130_fd_sc_hd__o211a_2
XFILLER_200_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28248_ _34450_/Q _24258_/X _28258_/S VGND VGND VPWR VPWR _28249_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18001_ _17860_/X _17999_/X _18000_/X _17865_/X VGND VGND VPWR VPWR _18001_/X sky130_fd_sc_hd__a22o_1
XFILLER_51_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16193_ _35537_/Q _35473_/Q _35409_/Q _35345_/Q _16191_/X _16192_/X VGND VGND VPWR
+ VPWR _16193_/X sky130_fd_sc_hd__mux4_1
X_28179_ _28179_/A VGND VGND VPWR VPWR _34417_/D sky130_fd_sc_hd__clkbuf_1
X_30210_ _35349_/Q _29073_/X _30214_/S VGND VGND VPWR VPWR _30211_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31190_ _35813_/Q input16/X _31202_/S VGND VGND VPWR VPWR _31191_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30141_ _30141_/A VGND VGND VPWR VPWR _35316_/D sky130_fd_sc_hd__clkbuf_1
X_19952_ _33787_/Q _33723_/Q _33659_/Q _33595_/Q _19849_/X _19850_/X VGND VGND VPWR
+ VPWR _19952_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18903_ _32477_/Q _32349_/Q _32029_/Q _35997_/Q _18870_/X _18658_/X VGND VGND VPWR
+ VPWR _18903_/X sky130_fd_sc_hd__mux4_1
X_30072_ _30072_/A VGND VGND VPWR VPWR _35283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19883_ _19877_/X _19882_/X _19814_/X VGND VGND VPWR VPWR _19884_/D sky130_fd_sc_hd__o21ba_1
XFILLER_49_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1010 _17908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1021 _17847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1032 _17865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33900_ _35574_/CLK _33900_/D VGND VGND VPWR VPWR _33900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18834_ _32731_/Q _32667_/Q _32603_/Q _36059_/Q _18513_/X _18650_/X VGND VGND VPWR
+ VPWR _18834_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1043 _17154_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_34880_ _35075_/CLK _34880_/D VGND VGND VPWR VPWR _34880_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1054 _16173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1065 _17056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1076 _17164_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33831_ _35943_/CLK _33831_/D VGND VGND VPWR VPWR _33831_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1087 _17232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18765_ _18761_/X _18764_/X _18722_/X VGND VGND VPWR VPWR _18787_/A sky130_fd_sc_hd__o21ba_1
XFILLER_3_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1098 _17330_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15977_ _17855_/A VGND VGND VPWR VPWR _15977_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17716_ _34556_/Q _32444_/Q _34428_/Q _34364_/Q _17578_/X _17579_/X VGND VGND VPWR
+ VPWR _17716_/X sky130_fd_sc_hd__mux4_1
XFILLER_208_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33762_ _34276_/CLK _33762_/D VGND VGND VPWR VPWR _33762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30974_ _35711_/Q _29203_/X _30974_/S VGND VGND VPWR VPWR _30975_/A sky130_fd_sc_hd__mux2_1
X_18696_ _18657_/X _18694_/X _18695_/X _18661_/X VGND VGND VPWR VPWR _18696_/X sky130_fd_sc_hd__a22o_1
XFILLER_36_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35501_ _35562_/CLK _35501_/D VGND VGND VPWR VPWR _35501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32713_ _36105_/CLK _32713_/D VGND VGND VPWR VPWR _32713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17647_ _35066_/Q _35002_/Q _34938_/Q _34874_/Q _17509_/X _17510_/X VGND VGND VPWR
+ VPWR _17647_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33693_ _34010_/CLK _33693_/D VGND VGND VPWR VPWR _33693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35432_ _35945_/CLK _35432_/D VGND VGND VPWR VPWR _35432_/Q sky130_fd_sc_hd__dfxtp_1
X_32644_ _36103_/CLK _32644_/D VGND VGND VPWR VPWR _32644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17578_ _17931_/A VGND VGND VPWR VPWR _17578_/X sky130_fd_sc_hd__buf_6
XFILLER_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19317_ _34281_/Q _34217_/Q _34153_/Q _34089_/Q _19036_/X _19037_/X VGND VGND VPWR
+ VPWR _19317_/X sky130_fd_sc_hd__mux4_1
XFILLER_188_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16529_ _16489_/X _16527_/X _16528_/X _16494_/X VGND VGND VPWR VPWR _16529_/X sky130_fd_sc_hd__a22o_1
X_35363_ _35552_/CLK _35363_/D VGND VGND VPWR VPWR _35363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32575_ _35906_/CLK _32575_/D VGND VGND VPWR VPWR _32575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34314_ _35851_/CLK _34314_/D VGND VGND VPWR VPWR _34314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31526_ _31526_/A VGND VGND VPWR VPWR _35972_/D sky130_fd_sc_hd__clkbuf_1
X_19248_ _19142_/X _19246_/X _19247_/X _19147_/X VGND VGND VPWR VPWR _19248_/X sky130_fd_sc_hd__a22o_1
X_35294_ _35294_/CLK _35294_/D VGND VGND VPWR VPWR _35294_/Q sky130_fd_sc_hd__dfxtp_1
X_34245_ _34308_/CLK _34245_/D VGND VGND VPWR VPWR _34245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31457_ _31457_/A VGND VGND VPWR VPWR _35939_/D sky130_fd_sc_hd__clkbuf_1
X_19179_ _19179_/A VGND VGND VPWR VPWR _32100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21210_ _35741_/Q _35101_/Q _34461_/Q _33821_/Q _21034_/X _21035_/X VGND VGND VPWR
+ VPWR _21210_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30408_ _30408_/A VGND VGND VPWR VPWR _35442_/D sky130_fd_sc_hd__clkbuf_1
X_34176_ _36160_/CLK _34176_/D VGND VGND VPWR VPWR _34176_/Q sky130_fd_sc_hd__dfxtp_1
X_22190_ _34041_/Q _33977_/Q _33913_/Q _32249_/Q _21973_/X _21974_/X VGND VGND VPWR
+ VPWR _22190_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_1216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31388_ _35907_/Q input49/X _31400_/S VGND VGND VPWR VPWR _31389_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_5_5_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_5_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_117_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21141_ _35803_/Q _32178_/Q _35675_/Q _35611_/Q _20854_/X _20855_/X VGND VGND VPWR
+ VPWR _21141_/X sky130_fd_sc_hd__mux4_1
X_33127_ _36135_/CLK _33127_/D VGND VGND VPWR VPWR _33127_/Q sky130_fd_sc_hd__dfxtp_1
X_30339_ _30339_/A VGND VGND VPWR VPWR _35409_/D sky130_fd_sc_hd__clkbuf_1
X_21072_ _21068_/X _21071_/X _21030_/X _21031_/X VGND VGND VPWR VPWR _21087_/B sky130_fd_sc_hd__o211a_1
X_33058_ _36130_/CLK _33058_/D VGND VGND VPWR VPWR _33058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20023_ _34301_/Q _34237_/Q _34173_/Q _34109_/Q _19742_/X _19743_/X VGND VGND VPWR
+ VPWR _20023_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32009_ _36194_/CLK _32009_/D VGND VGND VPWR VPWR _32009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24900_ _22945_/X _32931_/Q _24916_/S VGND VGND VPWR VPWR _24901_/A sky130_fd_sc_hd__mux2_1
X_25880_ _24998_/X _33360_/Q _25894_/S VGND VGND VPWR VPWR _25881_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24831_ _24831_/A VGND VGND VPWR VPWR _32898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27550_ _27550_/A VGND VGND VPWR VPWR _34120_/D sky130_fd_sc_hd__clkbuf_1
X_24762_ _24852_/S VGND VGND VPWR VPWR _24781_/S sky130_fd_sc_hd__buf_4
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21974_ _22447_/A VGND VGND VPWR VPWR _21974_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_227_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1001 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23713_ _22895_/X _32403_/Q _23721_/S VGND VGND VPWR VPWR _23714_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26501_ _26501_/A VGND VGND VPWR VPWR _33654_/D sky130_fd_sc_hd__clkbuf_1
X_20925_ _20921_/X _20924_/X _20640_/X _20642_/X VGND VGND VPWR VPWR _20940_/B sky130_fd_sc_hd__o211a_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27481_ _27481_/A VGND VGND VPWR VPWR _34087_/D sky130_fd_sc_hd__clkbuf_1
X_24693_ _23041_/X _32834_/Q _24707_/S VGND VGND VPWR VPWR _24694_/A sky130_fd_sc_hd__mux2_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29220_ _34884_/Q _29219_/X _29235_/S VGND VGND VPWR VPWR _29221_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26432_ _25016_/X _33622_/Q _26434_/S VGND VGND VPWR VPWR _26433_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23644_ _32372_/Q _23264_/X _23646_/S VGND VGND VPWR VPWR _23645_/A sky130_fd_sc_hd__mux2_1
X_20856_ _35795_/Q _32169_/Q _35667_/Q _35603_/Q _20854_/X _20855_/X VGND VGND VPWR
+ VPWR _20856_/X sky130_fd_sc_hd__mux4_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_968 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29151_ input26/X VGND VGND VPWR VPWR _29151_/X sky130_fd_sc_hd__clkbuf_4
X_26363_ _26363_/A VGND VGND VPWR VPWR _33589_/D sky130_fd_sc_hd__clkbuf_1
X_23575_ _32339_/Q _23102_/X _23583_/S VGND VGND VPWR VPWR _23576_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20787_ _20783_/X _20786_/X _20640_/X _20642_/X VGND VGND VPWR VPWR _20804_/B sky130_fd_sc_hd__o211a_1
XFILLER_211_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28102_ _28102_/A VGND VGND VPWR VPWR _34381_/D sky130_fd_sc_hd__clkbuf_1
X_25314_ _25174_/X _33097_/Q _25314_/S VGND VGND VPWR VPWR _25315_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22526_ _22305_/X _22524_/X _22525_/X _22308_/X VGND VGND VPWR VPWR _22526_/X sky130_fd_sc_hd__a22o_1
XFILLER_168_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26294_ _26294_/A VGND VGND VPWR VPWR _33556_/D sky130_fd_sc_hd__clkbuf_1
X_29082_ input2/X VGND VGND VPWR VPWR _29082_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_210_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28033_ _26915_/X _34348_/Q _28051_/S VGND VGND VPWR VPWR _28034_/A sky130_fd_sc_hd__mux2_1
X_25245_ _25072_/X _33064_/Q _25251_/S VGND VGND VPWR VPWR _25246_/A sky130_fd_sc_hd__mux2_1
X_22457_ _35328_/Q _35264_/Q _35200_/Q _32320_/Q _22312_/X _22313_/X VGND VGND VPWR
+ VPWR _22457_/X sky130_fd_sc_hd__mux4_1
X_21408_ _22467_/A VGND VGND VPWR VPWR _21408_/X sky130_fd_sc_hd__buf_2
XFILLER_202_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25176_ _25176_/A VGND VGND VPWR VPWR _33033_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22388_ _34558_/Q _32446_/Q _34430_/Q _34366_/Q _22178_/X _22179_/X VGND VGND VPWR
+ VPWR _22388_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24127_ _22904_/X _32598_/Q _24129_/S VGND VGND VPWR VPWR _24128_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21339_ _21089_/X _21335_/X _21338_/X _21094_/X VGND VGND VPWR VPWR _21339_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29984_ _35242_/Q _29138_/X _29986_/S VGND VGND VPWR VPWR _29985_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24058_ _24106_/S VGND VGND VPWR VPWR _24077_/S sky130_fd_sc_hd__buf_4
XFILLER_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28935_ _28998_/A VGND VGND VPWR VPWR _28954_/S sky130_fd_sc_hd__buf_4
XFILLER_137_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23009_ _23009_/A VGND VGND VPWR VPWR _32055_/D sky130_fd_sc_hd__clkbuf_1
X_16880_ _33765_/Q _33701_/Q _33637_/Q _33573_/Q _16843_/X _16844_/X VGND VGND VPWR
+ VPWR _16880_/X sky130_fd_sc_hd__mux4_1
X_28866_ _26950_/X _34743_/Q _28882_/S VGND VGND VPWR VPWR _28867_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27817_ _34246_/Q _24419_/X _27823_/S VGND VGND VPWR VPWR _27818_/A sky130_fd_sc_hd__mux2_1
XTAP_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28797_ _28797_/A VGND VGND VPWR VPWR _34710_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18550_ _32467_/Q _32339_/Q _32019_/Q _35987_/Q _18517_/X _20163_/A VGND VGND VPWR
+ VPWR _18550_/X sky130_fd_sc_hd__mux4_1
XTAP_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27748_ _34213_/Q _24317_/X _27760_/S VGND VGND VPWR VPWR _27749_/A sky130_fd_sc_hd__mux2_1
XTAP_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ _17496_/X _17499_/X _17500_/X VGND VGND VPWR VPWR _17516_/C sky130_fd_sc_hd__o21ba_1
XTAP_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18481_ _32721_/Q _32657_/Q _32593_/Q _36049_/Q _20162_/A _20013_/A VGND VGND VPWR
+ VPWR _18481_/X sky130_fd_sc_hd__mux4_1
XTAP_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27679_ _27679_/A VGND VGND VPWR VPWR _34180_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_430 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_441 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29418_ _29418_/A VGND VGND VPWR VPWR _34973_/D sky130_fd_sc_hd__clkbuf_1
X_17432_ _34804_/Q _34740_/Q _34676_/Q _34612_/Q _17288_/X _17289_/X VGND VGND VPWR
+ VPWR _17432_/X sky130_fd_sc_hd__mux4_1
XFILLER_75_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_452 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_463 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_474 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30690_ _35576_/Q _29182_/X _30704_/S VGND VGND VPWR VPWR _30691_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_485 _31994_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_496 _32005_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29349_ _23294_/X _34941_/Q _29353_/S VGND VGND VPWR VPWR _29350_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17363_ _34546_/Q _32434_/Q _34418_/Q _34354_/Q _17225_/X _17226_/X VGND VGND VPWR
+ VPWR _17363_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19102_ _34530_/Q _32418_/Q _34402_/Q _34338_/Q _18819_/X _18820_/X VGND VGND VPWR
+ VPWR _19102_/X sky130_fd_sc_hd__mux4_1
XFILLER_207_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16314_ _17846_/A VGND VGND VPWR VPWR _16314_/X sky130_fd_sc_hd__buf_6
X_32360_ _36072_/CLK _32360_/D VGND VGND VPWR VPWR _32360_/Q sky130_fd_sc_hd__dfxtp_1
X_17294_ _35056_/Q _34992_/Q _34928_/Q _34864_/Q _17156_/X _17157_/X VGND VGND VPWR
+ VPWR _17294_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31311_ _31311_/A VGND VGND VPWR VPWR _35870_/D sky130_fd_sc_hd__clkbuf_1
X_19033_ _19033_/A _19033_/B _19033_/C _19033_/D VGND VGND VPWR VPWR _19034_/A sky130_fd_sc_hd__or4_1
X_16245_ _16143_/X _16243_/X _16244_/X _16146_/X VGND VGND VPWR VPWR _16245_/X sky130_fd_sc_hd__a22o_1
XFILLER_220_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32291_ _35298_/CLK _32291_/D VGND VGND VPWR VPWR _32291_/Q sky130_fd_sc_hd__dfxtp_1
X_34030_ _34032_/CLK _34030_/D VGND VGND VPWR VPWR _34030_/Q sky130_fd_sc_hd__dfxtp_1
X_31242_ _35838_/Q input43/X _31244_/S VGND VGND VPWR VPWR _31243_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16176_ _16136_/X _16174_/X _16175_/X _16141_/X VGND VGND VPWR VPWR _16176_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput106 _31974_/Q VGND VGND VPWR VPWR D1[24] sky130_fd_sc_hd__buf_2
XFILLER_217_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput117 _31984_/Q VGND VGND VPWR VPWR D1[34] sky130_fd_sc_hd__buf_2
XFILLER_173_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput128 _31994_/Q VGND VGND VPWR VPWR D1[44] sky130_fd_sc_hd__buf_2
X_31173_ _35805_/Q input7/X _31181_/S VGND VGND VPWR VPWR _31174_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput139 _32004_/Q VGND VGND VPWR VPWR D1[54] sky130_fd_sc_hd__buf_2
XFILLER_142_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19935_ _35770_/Q _35130_/Q _34490_/Q _33850_/Q _19793_/X _19794_/X VGND VGND VPWR
+ VPWR _19935_/X sky130_fd_sc_hd__mux4_1
X_30124_ _35308_/Q _29144_/X _30142_/S VGND VGND VPWR VPWR _30125_/A sky130_fd_sc_hd__mux2_1
X_35981_ _35981_/CLK _35981_/D VGND VGND VPWR VPWR _35981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30055_ _35276_/Q _29243_/X _30057_/S VGND VGND VPWR VPWR _30056_/A sky130_fd_sc_hd__mux2_1
X_34932_ _34932_/CLK _34932_/D VGND VGND VPWR VPWR _34932_/Q sky130_fd_sc_hd__dfxtp_1
X_19866_ _19716_/X _19864_/X _19865_/X _19720_/X VGND VGND VPWR VPWR _19866_/X sky130_fd_sc_hd__a22o_1
XFILLER_96_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18817_ _35290_/Q _35226_/Q _35162_/Q _32282_/Q _18600_/X _18601_/X VGND VGND VPWR
+ VPWR _18817_/X sky130_fd_sc_hd__mux4_1
X_34863_ _35758_/CLK _34863_/D VGND VGND VPWR VPWR _34863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19797_ _35574_/Q _35510_/Q _35446_/Q _35382_/Q _19550_/X _19551_/X VGND VGND VPWR
+ VPWR _19797_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33814_ _35733_/CLK _33814_/D VGND VGND VPWR VPWR _33814_/Q sky130_fd_sc_hd__dfxtp_1
X_18748_ _19454_/A VGND VGND VPWR VPWR _18748_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34794_ _34794_/CLK _34794_/D VGND VGND VPWR VPWR _34794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33745_ _34259_/CLK _33745_/D VGND VGND VPWR VPWR _33745_/Q sky130_fd_sc_hd__dfxtp_1
X_18679_ _18675_/X _18678_/X _18400_/X VGND VGND VPWR VPWR _18680_/D sky130_fd_sc_hd__o21ba_1
X_30957_ _30957_/A VGND VGND VPWR VPWR _35702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20710_ _33999_/Q _33935_/Q _33871_/Q _32143_/Q _20708_/X _20709_/X VGND VGND VPWR
+ VPWR _20710_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33676_ _34317_/CLK _33676_/D VGND VGND VPWR VPWR _33676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21690_ _22557_/A VGND VGND VPWR VPWR _21690_/X sky130_fd_sc_hd__buf_4
X_30888_ _35670_/Q _29076_/X _30890_/S VGND VGND VPWR VPWR _30889_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35415_ _35863_/CLK _35415_/D VGND VGND VPWR VPWR _35415_/Q sky130_fd_sc_hd__dfxtp_1
X_20641_ input76/X VGND VGND VPWR VPWR _22443_/A sky130_fd_sc_hd__buf_12
XFILLER_11_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32627_ _36018_/CLK _32627_/D VGND VGND VPWR VPWR _32627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35346_ _35922_/CLK _35346_/D VGND VGND VPWR VPWR _35346_/Q sky130_fd_sc_hd__dfxtp_1
X_23360_ _23360_/A VGND VGND VPWR VPWR _32239_/D sky130_fd_sc_hd__clkbuf_1
X_20572_ _20568_/X _20571_/X _20167_/A VGND VGND VPWR VPWR _20573_/D sky130_fd_sc_hd__o21ba_1
XFILLER_149_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32558_ _35950_/CLK _32558_/D VGND VGND VPWR VPWR _32558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22311_ _34812_/Q _34748_/Q _34684_/Q _34620_/Q _22241_/X _22242_/X VGND VGND VPWR
+ VPWR _22311_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31509_ _31509_/A VGND VGND VPWR VPWR _35964_/D sky130_fd_sc_hd__clkbuf_1
X_35277_ _35277_/CLK _35277_/D VGND VGND VPWR VPWR _35277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23291_ _23291_/A VGND VGND VPWR VPWR _32214_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32489_ _36009_/CLK _32489_/D VGND VGND VPWR VPWR _32489_/Q sky130_fd_sc_hd__dfxtp_1
X_25030_ _25029_/X _32986_/Q _25051_/S VGND VGND VPWR VPWR _25031_/A sky130_fd_sc_hd__mux2_1
X_22242_ _22595_/A VGND VGND VPWR VPWR _22242_/X sky130_fd_sc_hd__buf_6
X_34228_ _34228_/CLK _34228_/D VGND VGND VPWR VPWR _34228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22173_ _21952_/X _22171_/X _22172_/X _21955_/X VGND VGND VPWR VPWR _22173_/X sky130_fd_sc_hd__a22o_1
X_34159_ _34286_/CLK _34159_/D VGND VGND VPWR VPWR _34159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21124_ _21118_/X _21123_/X _21055_/X VGND VGND VPWR VPWR _21125_/D sky130_fd_sc_hd__o21ba_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26981_ input47/X VGND VGND VPWR VPWR _26981_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_120_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28720_ _26934_/X _34674_/Q _28726_/S VGND VGND VPWR VPWR _28721_/A sky130_fd_sc_hd__mux2_1
X_25932_ _25075_/X _33385_/Q _25936_/S VGND VGND VPWR VPWR _25933_/A sky130_fd_sc_hd__mux2_1
X_21055_ _22467_/A VGND VGND VPWR VPWR _21055_/X sky130_fd_sc_hd__buf_2
XFILLER_154_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20006_ _35580_/Q _35516_/Q _35452_/Q _35388_/Q _19903_/X _19904_/X VGND VGND VPWR
+ VPWR _20006_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28651_ _26832_/X _34641_/Q _28663_/S VGND VGND VPWR VPWR _28652_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25863_ _25863_/A VGND VGND VPWR VPWR _33352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27602_ _34144_/Q _24301_/X _27604_/S VGND VGND VPWR VPWR _27603_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24814_ _24814_/A VGND VGND VPWR VPWR _32890_/D sky130_fd_sc_hd__clkbuf_1
X_28582_ _28582_/A VGND VGND VPWR VPWR _34608_/D sky130_fd_sc_hd__clkbuf_1
X_25794_ _25794_/A VGND VGND VPWR VPWR _33319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_228_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27533_ _26977_/X _34112_/Q _27551_/S VGND VGND VPWR VPWR _27534_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24745_ _24745_/A VGND VGND VPWR VPWR _32857_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21957_ _21951_/X _21956_/X _21747_/X VGND VGND VPWR VPWR _21967_/C sky130_fd_sc_hd__o21ba_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_270_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _34303_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ _20908_/A _20908_/B _20908_/C _20908_/D VGND VGND VPWR VPWR _20909_/A sky130_fd_sc_hd__or4_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24676_ _23016_/X _32826_/Q _24686_/S VGND VGND VPWR VPWR _24677_/A sky130_fd_sc_hd__mux2_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27464_ _27464_/A VGND VGND VPWR VPWR _34079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21888_ _22594_/A VGND VGND VPWR VPWR _21888_/X sky130_fd_sc_hd__buf_6
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29203_ input44/X VGND VGND VPWR VPWR _29203_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26415_ _26547_/S VGND VGND VPWR VPWR _26434_/S sky130_fd_sc_hd__buf_4
XFILLER_39_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23627_ _23696_/S VGND VGND VPWR VPWR _23646_/S sky130_fd_sc_hd__buf_6
X_20839_ _20839_/A VGND VGND VPWR VPWR _36178_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27395_ _34047_/Q _24397_/X _27395_/S VGND VGND VPWR VPWR _27396_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29134_ _29134_/A VGND VGND VPWR VPWR _34856_/D sky130_fd_sc_hd__clkbuf_1
X_23558_ _23558_/A VGND VGND VPWR VPWR _32332_/D sky130_fd_sc_hd__clkbuf_1
X_26346_ _25088_/X _33581_/Q _26362_/S VGND VGND VPWR VPWR _26347_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22509_ _33538_/Q _33474_/Q _33410_/Q _33346_/Q _22429_/X _22430_/X VGND VGND VPWR
+ VPWR _22509_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput19 DW[26] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__buf_4
XFILLER_195_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26277_ _25186_/X _33549_/Q _26277_/S VGND VGND VPWR VPWR _26278_/A sky130_fd_sc_hd__mux2_1
X_29065_ _34834_/Q _29064_/X _29080_/S VGND VGND VPWR VPWR _29066_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23489_ _23489_/A VGND VGND VPWR VPWR _32299_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16030_ _17770_/A VGND VGND VPWR VPWR _17863_/A sky130_fd_sc_hd__buf_4
X_28016_ _26891_/X _34340_/Q _28030_/S VGND VGND VPWR VPWR _28017_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25228_ _25047_/X _33056_/Q _25230_/S VGND VGND VPWR VPWR _25229_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25159_ input50/X VGND VGND VPWR VPWR _25159_/X sky130_fd_sc_hd__buf_2
X_17981_ _17761_/X _17979_/X _17980_/X _17767_/X VGND VGND VPWR VPWR _17981_/X sky130_fd_sc_hd__a22o_1
X_29967_ _30057_/S VGND VGND VPWR VPWR _29986_/S sky130_fd_sc_hd__buf_6
XFILLER_97_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19720_ _20211_/A VGND VGND VPWR VPWR _19720_/X sky130_fd_sc_hd__clkbuf_4
X_28918_ _28918_/A VGND VGND VPWR VPWR _34767_/D sky130_fd_sc_hd__clkbuf_1
X_16932_ _33190_/Q _32550_/Q _35942_/Q _35878_/Q _16721_/X _16722_/X VGND VGND VPWR
+ VPWR _16932_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29898_ _35201_/Q _29210_/X _29914_/S VGND VGND VPWR VPWR _29899_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19651_ _19647_/X _19648_/X _19649_/X _19650_/X VGND VGND VPWR VPWR _19651_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16863_ _35748_/Q _35108_/Q _34468_/Q _33828_/Q _16787_/X _16788_/X VGND VGND VPWR
+ VPWR _16863_/X sky130_fd_sc_hd__mux4_1
X_28849_ _26925_/X _34735_/Q _28861_/S VGND VGND VPWR VPWR _28850_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18602_ _35284_/Q _35220_/Q _35156_/Q _32276_/Q _18600_/X _18601_/X VGND VGND VPWR
+ VPWR _18602_/X sky130_fd_sc_hd__mux4_1
X_19582_ _35760_/Q _35120_/Q _34480_/Q _33840_/Q _19440_/X _19441_/X VGND VGND VPWR
+ VPWR _19582_/X sky130_fd_sc_hd__mux4_1
X_31860_ _31860_/A VGND VGND VPWR VPWR _36130_/D sky130_fd_sc_hd__clkbuf_1
X_16794_ _17853_/A VGND VGND VPWR VPWR _16794_/X sky130_fd_sc_hd__buf_2
XFILLER_206_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18533_ _18374_/X _18531_/X _18532_/X _18384_/X VGND VGND VPWR VPWR _18533_/X sky130_fd_sc_hd__a22o_1
X_30811_ _30811_/A VGND VGND VPWR VPWR _35633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31791_ _36098_/Q input48/X _31805_/S VGND VGND VPWR VPWR _31792_/A sky130_fd_sc_hd__mux2_1
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_261_CLK clkbuf_6_60__f_CLK/X VGND VGND VPWR VPWR _32962_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33530_ _33787_/CLK _33530_/D VGND VGND VPWR VPWR _33530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30742_ _30742_/A VGND VGND VPWR VPWR _35600_/D sky130_fd_sc_hd__clkbuf_1
X_18464_ _35280_/Q _35216_/Q _35152_/Q _32272_/Q _18379_/X _18381_/X VGND VGND VPWR
+ VPWR _18464_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_260 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_271 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_282 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17415_ _17408_/X _17410_/X _17413_/X _17414_/X VGND VGND VPWR VPWR _17415_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_293 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33461_ _33780_/CLK _33461_/D VGND VGND VPWR VPWR _33461_/Q sky130_fd_sc_hd__dfxtp_1
X_18395_ _35022_/Q _34958_/Q _34894_/Q _34830_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _18395_/X sky130_fd_sc_hd__mux4_1
X_30673_ _35568_/Q _29157_/X _30683_/S VGND VGND VPWR VPWR _30674_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35200_ _35328_/CLK _35200_/D VGND VGND VPWR VPWR _35200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32412_ _35166_/CLK _32412_/D VGND VGND VPWR VPWR _32412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36180_ _36202_/CLK _36180_/D VGND VGND VPWR VPWR _36180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17346_ _17340_/X _17345_/X _17136_/X _17137_/X VGND VGND VPWR VPWR _17367_/B sky130_fd_sc_hd__o211a_1
XFILLER_105_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33392_ _33520_/CLK _33392_/D VGND VGND VPWR VPWR _33392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35131_ _35963_/CLK _35131_/D VGND VGND VPWR VPWR _35131_/Q sky130_fd_sc_hd__dfxtp_1
X_32343_ _36116_/CLK _32343_/D VGND VGND VPWR VPWR _32343_/Q sky130_fd_sc_hd__dfxtp_1
X_17277_ _32496_/Q _32368_/Q _32048_/Q _36016_/Q _17276_/X _17064_/X VGND VGND VPWR
+ VPWR _17277_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19016_ _19009_/X _19015_/X _18730_/X _18731_/X VGND VGND VPWR VPWR _19033_/B sky130_fd_sc_hd__o211a_2
X_16228_ _16224_/X _16227_/X _16071_/X VGND VGND VPWR VPWR _16238_/C sky130_fd_sc_hd__o21ba_1
X_35062_ _35257_/CLK _35062_/D VGND VGND VPWR VPWR _35062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32274_ _35026_/CLK _32274_/D VGND VGND VPWR VPWR _32274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34013_ _34142_/CLK _34013_/D VGND VGND VPWR VPWR _34013_/Q sky130_fd_sc_hd__dfxtp_1
X_31225_ _31273_/S VGND VGND VPWR VPWR _31244_/S sky130_fd_sc_hd__buf_4
X_16159_ _35536_/Q _35472_/Q _35408_/Q _35344_/Q _16058_/X _16060_/X VGND VGND VPWR
+ VPWR _16159_/X sky130_fd_sc_hd__mux4_1
XFILLER_115_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31156_ _35797_/Q input62/X _31160_/S VGND VGND VPWR VPWR _31157_/A sky130_fd_sc_hd__mux2_1
X_30107_ _35300_/Q _29120_/X _30121_/S VGND VGND VPWR VPWR _30108_/A sky130_fd_sc_hd__mux2_1
X_19918_ _33786_/Q _33722_/Q _33658_/Q _33594_/Q _19849_/X _19850_/X VGND VGND VPWR
+ VPWR _19918_/X sky130_fd_sc_hd__mux4_1
X_35964_ _35965_/CLK _35964_/D VGND VGND VPWR VPWR _35964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31087_ _31087_/A VGND VGND VPWR VPWR _35764_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30038_ _30038_/A VGND VGND VPWR VPWR _35267_/D sky130_fd_sc_hd__clkbuf_1
X_19849_ _20202_/A VGND VGND VPWR VPWR _19849_/X sky130_fd_sc_hd__buf_4
X_34915_ _35299_/CLK _34915_/D VGND VGND VPWR VPWR _34915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35895_ _36023_/CLK _35895_/D VGND VGND VPWR VPWR _35895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22860_ _35789_/Q _35149_/Q _34509_/Q _33869_/Q _20708_/X _20709_/X VGND VGND VPWR
+ VPWR _22860_/X sky130_fd_sc_hd__mux4_1
XFILLER_216_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34846_ _35038_/CLK _34846_/D VGND VGND VPWR VPWR _34846_/Q sky130_fd_sc_hd__dfxtp_1
X_21811_ _32494_/Q _32366_/Q _32046_/Q _36014_/Q _21523_/X _21664_/X VGND VGND VPWR
+ VPWR _21811_/X sky130_fd_sc_hd__mux4_1
X_22791_ _22787_/X _22790_/X _22434_/A VGND VGND VPWR VPWR _22813_/A sky130_fd_sc_hd__o21ba_1
X_34777_ _34777_/CLK _34777_/D VGND VGND VPWR VPWR _34777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31989_ _36201_/CLK _31989_/D VGND VGND VPWR VPWR _31989_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_252_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _34050_/CLK sky130_fd_sc_hd__clkbuf_16
X_24530_ _23003_/X _32758_/Q _24548_/S VGND VGND VPWR VPWR _24531_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33728_ _33793_/CLK _33728_/D VGND VGND VPWR VPWR _33728_/Q sky130_fd_sc_hd__dfxtp_1
X_21742_ _35756_/Q _35116_/Q _34476_/Q _33836_/Q _21740_/X _21741_/X VGND VGND VPWR
+ VPWR _21742_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_1053 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24461_ _24461_/A VGND VGND VPWR VPWR _32725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_212_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33659_ _34044_/CLK _33659_/D VGND VGND VPWR VPWR _33659_/Q sky130_fd_sc_hd__dfxtp_1
X_21673_ _35562_/Q _35498_/Q _35434_/Q _35370_/Q _21497_/X _21498_/X VGND VGND VPWR
+ VPWR _21673_/X sky130_fd_sc_hd__mux4_1
XFILLER_212_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23412_ _23412_/A VGND VGND VPWR VPWR _32264_/D sky130_fd_sc_hd__clkbuf_1
X_26200_ _25072_/X _33512_/Q _26206_/S VGND VGND VPWR VPWR _26201_/A sky130_fd_sc_hd__mux2_1
X_20624_ _20614_/X _20619_/X _20622_/X _20623_/X VGND VGND VPWR VPWR _20624_/X sky130_fd_sc_hd__a22o_1
X_27180_ _27180_/A VGND VGND VPWR VPWR _33944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24392_ _32701_/Q _24391_/X _24398_/S VGND VGND VPWR VPWR _24393_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26131_ _26131_/A VGND VGND VPWR VPWR _33479_/D sky130_fd_sc_hd__clkbuf_1
X_35329_ _35330_/CLK _35329_/D VGND VGND VPWR VPWR _35329_/Q sky130_fd_sc_hd__dfxtp_1
X_23343_ _32232_/Q _23342_/X _23346_/S VGND VGND VPWR VPWR _23344_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20555_ _32525_/Q _32397_/Q _32077_/Q _36045_/Q _20282_/X _19307_/A VGND VGND VPWR
+ VPWR _20555_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26062_ _26062_/A VGND VGND VPWR VPWR _33446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23274_ input36/X VGND VGND VPWR VPWR _23274_/X sky130_fd_sc_hd__buf_4
X_20486_ _34315_/Q _34251_/Q _34187_/Q _34123_/Q _18345_/X _18346_/X VGND VGND VPWR
+ VPWR _20486_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25013_ input62/X VGND VGND VPWR VPWR _25013_/X sky130_fd_sc_hd__clkbuf_8
X_22225_ _22578_/A VGND VGND VPWR VPWR _22225_/X sky130_fd_sc_hd__buf_6
XFILLER_106_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29821_ _29821_/A VGND VGND VPWR VPWR _35164_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22156_ _33528_/Q _33464_/Q _33400_/Q _33336_/Q _22076_/X _22077_/X VGND VGND VPWR
+ VPWR _22156_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21107_ _20957_/X _21105_/X _21106_/X _20961_/X VGND VGND VPWR VPWR _21107_/X sky130_fd_sc_hd__a22o_1
XFILLER_154_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29752_ _35132_/Q _29194_/X _29758_/S VGND VGND VPWR VPWR _29753_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26964_ _26964_/A VGND VGND VPWR VPWR _33851_/D sky130_fd_sc_hd__clkbuf_1
X_22087_ _33014_/Q _32950_/Q _32886_/Q _32822_/Q _21942_/X _21943_/X VGND VGND VPWR
+ VPWR _22087_/X sky130_fd_sc_hd__mux4_1
XTAP_6869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28703_ _26909_/X _34666_/Q _28705_/S VGND VGND VPWR VPWR _28704_/A sky130_fd_sc_hd__mux2_1
X_25915_ _25050_/X _33377_/Q _25915_/S VGND VGND VPWR VPWR _25916_/A sky130_fd_sc_hd__mux2_1
X_21038_ _35544_/Q _35480_/Q _35416_/Q _35352_/Q _20791_/X _20792_/X VGND VGND VPWR
+ VPWR _21038_/X sky130_fd_sc_hd__mux4_1
XFILLER_102_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29683_ _35099_/Q _29092_/X _29695_/S VGND VGND VPWR VPWR _29684_/A sky130_fd_sc_hd__mux2_1
X_26895_ _26894_/X _33829_/Q _26913_/S VGND VGND VPWR VPWR _26896_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_491_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _35745_/CLK sky130_fd_sc_hd__clkbuf_16
X_28634_ _28634_/A VGND VGND VPWR VPWR _34633_/D sky130_fd_sc_hd__clkbuf_1
X_25846_ _25146_/X _33344_/Q _25864_/S VGND VGND VPWR VPWR _25847_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28565_ _28565_/A VGND VGND VPWR VPWR _34600_/D sky130_fd_sc_hd__clkbuf_1
X_22989_ _22988_/X _32049_/Q _23001_/S VGND VGND VPWR VPWR _22990_/A sky130_fd_sc_hd__mux2_1
X_25777_ _25777_/A VGND VGND VPWR VPWR _33311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_243_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _34310_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27516_ _26953_/X _34104_/Q _27530_/S VGND VGND VPWR VPWR _27517_/A sky130_fd_sc_hd__mux2_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24728_ _24728_/A VGND VGND VPWR VPWR _32849_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28496_ _27002_/X _34568_/Q _28498_/S VGND VGND VPWR VPWR _28497_/A sky130_fd_sc_hd__mux2_1
XFILLER_231_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27447_ _27447_/A VGND VGND VPWR VPWR _34071_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24659_ _22991_/X _32818_/Q _24665_/S VGND VGND VPWR VPWR _24660_/A sky130_fd_sc_hd__mux2_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17200_ _17906_/A VGND VGND VPWR VPWR _17200_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_208_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18180_ _35082_/Q _35018_/Q _34954_/Q _34890_/Q _16079_/X _16081_/X VGND VGND VPWR
+ VPWR _18180_/X sky130_fd_sc_hd__mux4_1
XFILLER_187_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27378_ _27378_/A VGND VGND VPWR VPWR _34038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29117_ input14/X VGND VGND VPWR VPWR _29117_/X sky130_fd_sc_hd__buf_2
X_17131_ _33260_/Q _36140_/Q _33132_/Q _33068_/Q _17058_/X _17059_/X VGND VGND VPWR
+ VPWR _17131_/X sky130_fd_sc_hd__mux4_1
X_26329_ _25063_/X _33573_/Q _26341_/S VGND VGND VPWR VPWR _26330_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_954 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29048_ input1/X VGND VGND VPWR VPWR _29048_/X sky130_fd_sc_hd__clkbuf_4
X_17062_ _17055_/X _17057_/X _17060_/X _17061_/X VGND VGND VPWR VPWR _17062_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16013_ _17761_/A VGND VGND VPWR VPWR _17901_/A sky130_fd_sc_hd__buf_12
XFILLER_87_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31010_ _31010_/A VGND VGND VPWR VPWR _35727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ _17855_/X _17962_/X _17963_/X _17858_/X VGND VGND VPWR VPWR _17964_/X sky130_fd_sc_hd__a22o_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19703_ _19495_/X _19701_/X _19702_/X _19500_/X VGND VGND VPWR VPWR _19703_/X sky130_fd_sc_hd__a22o_1
XFILLER_211_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16915_ _33510_/Q _33446_/Q _33382_/Q _33318_/Q _16770_/X _16771_/X VGND VGND VPWR
+ VPWR _16915_/X sky130_fd_sc_hd__mux4_1
X_32961_ _36098_/CLK _32961_/D VGND VGND VPWR VPWR _32961_/Q sky130_fd_sc_hd__dfxtp_1
X_17895_ _34561_/Q _32449_/Q _34433_/Q _34369_/Q _17578_/X _17579_/X VGND VGND VPWR
+ VPWR _17895_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_482_CLK clkbuf_6_3__f_CLK/X VGND VGND VPWR VPWR _35869_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_93_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34700_ _35341_/CLK _34700_/D VGND VGND VPWR VPWR _34700_/Q sky130_fd_sc_hd__dfxtp_1
X_31912_ _31912_/A VGND VGND VPWR VPWR _36155_/D sky130_fd_sc_hd__clkbuf_1
X_19634_ _33522_/Q _33458_/Q _33394_/Q _33330_/Q _19423_/X _19424_/X VGND VGND VPWR
+ VPWR _19634_/X sky130_fd_sc_hd__mux4_1
X_35680_ _35809_/CLK _35680_/D VGND VGND VPWR VPWR _35680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16846_ _34276_/Q _34212_/Q _34148_/Q _34084_/Q _16736_/X _16737_/X VGND VGND VPWR
+ VPWR _16846_/X sky130_fd_sc_hd__mux4_1
X_32892_ _36029_/CLK _32892_/D VGND VGND VPWR VPWR _32892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34631_ _34822_/CLK _34631_/D VGND VGND VPWR VPWR _34631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19565_ _33776_/Q _33712_/Q _33648_/Q _33584_/Q _19496_/X _19497_/X VGND VGND VPWR
+ VPWR _19565_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31843_ _31843_/A VGND VGND VPWR VPWR _36122_/D sky130_fd_sc_hd__clkbuf_1
X_16777_ _32738_/Q _32674_/Q _32610_/Q _36066_/Q _16566_/X _16703_/X VGND VGND VPWR
+ VPWR _16777_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_234_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _34752_/CLK sky130_fd_sc_hd__clkbuf_16
X_18516_ _18314_/X _18514_/X _18515_/X _18323_/X VGND VGND VPWR VPWR _18516_/X sky130_fd_sc_hd__a22o_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34562_ _34562_/CLK _34562_/D VGND VGND VPWR VPWR _34562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31774_ _36090_/Q input39/X _31784_/S VGND VGND VPWR VPWR _31775_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19496_ _20202_/A VGND VGND VPWR VPWR _19496_/X sky130_fd_sc_hd__buf_4
XFILLER_55_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33513_ _35386_/CLK _33513_/D VGND VGND VPWR VPWR _33513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18447_ _18443_/X _18444_/X _18445_/X _18446_/X VGND VGND VPWR VPWR _18447_/X sky130_fd_sc_hd__a22o_1
X_30725_ _35593_/Q _29234_/X _30725_/S VGND VGND VPWR VPWR _30726_/A sky130_fd_sc_hd__mux2_1
X_34493_ _35837_/CLK _34493_/D VGND VGND VPWR VPWR _34493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36232_ _36232_/CLK _36232_/D VGND VGND VPWR VPWR _36232_/Q sky130_fd_sc_hd__dfxtp_1
X_33444_ _33507_/CLK _33444_/D VGND VGND VPWR VPWR _33444_/Q sky130_fd_sc_hd__dfxtp_1
X_18378_ _20278_/A VGND VGND VPWR VPWR _20012_/A sky130_fd_sc_hd__buf_12
XFILLER_18_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30656_ _35560_/Q _29132_/X _30662_/S VGND VGND VPWR VPWR _30657_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_1032 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36163_ _36165_/CLK _36163_/D VGND VGND VPWR VPWR _36163_/Q sky130_fd_sc_hd__dfxtp_1
X_17329_ _17329_/A _17329_/B _17329_/C _17329_/D VGND VGND VPWR VPWR _17330_/A sky130_fd_sc_hd__or4_4
XFILLER_146_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33375_ _33692_/CLK _33375_/D VGND VGND VPWR VPWR _33375_/Q sky130_fd_sc_hd__dfxtp_1
X_30587_ _30587_/A VGND VGND VPWR VPWR _35527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35114_ _35945_/CLK _35114_/D VGND VGND VPWR VPWR _35114_/Q sky130_fd_sc_hd__dfxtp_1
X_32326_ _35334_/CLK _32326_/D VGND VGND VPWR VPWR _32326_/Q sky130_fd_sc_hd__dfxtp_1
X_20340_ _20208_/X _20338_/X _20339_/X _20211_/X VGND VGND VPWR VPWR _20340_/X sky130_fd_sc_hd__a22o_1
X_36094_ _36095_/CLK _36094_/D VGND VGND VPWR VPWR _36094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_49__f_CLK clkbuf_5_24_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_49__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_35045_ _35941_/CLK _35045_/D VGND VGND VPWR VPWR _35045_/Q sky130_fd_sc_hd__dfxtp_1
X_20271_ _33796_/Q _33732_/Q _33668_/Q _33604_/Q _20202_/X _20203_/X VGND VGND VPWR
+ VPWR _20271_/X sky130_fd_sc_hd__mux4_1
X_32257_ _36165_/CLK _32257_/D VGND VGND VPWR VPWR _32257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22010_ _32756_/Q _32692_/Q _32628_/Q _36084_/Q _21872_/X _22009_/X VGND VGND VPWR
+ VPWR _22010_/X sky130_fd_sc_hd__mux4_1
X_31208_ _31208_/A VGND VGND VPWR VPWR _35821_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32188_ _35811_/CLK _32188_/D VGND VGND VPWR VPWR _32188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31139_ _31139_/A VGND VGND VPWR VPWR _35789_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23961_ _23961_/A VGND VGND VPWR VPWR _32520_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35947_ _35947_/CLK _35947_/D VGND VGND VPWR VPWR _35947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25700_ _33276_/Q _24388_/X _25706_/S VGND VGND VPWR VPWR _25701_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_473_CLK clkbuf_6_8__f_CLK/X VGND VGND VPWR VPWR _35940_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22912_ _22910_/X _32024_/Q _22939_/S VGND VGND VPWR VPWR _22913_/A sky130_fd_sc_hd__mux2_1
X_26680_ _26680_/A VGND VGND VPWR VPWR _33739_/D sky130_fd_sc_hd__clkbuf_1
X_23892_ _23892_/A VGND VGND VPWR VPWR _32487_/D sky130_fd_sc_hd__clkbuf_1
X_35878_ _35942_/CLK _35878_/D VGND VGND VPWR VPWR _35878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22843_ _22843_/A _22843_/B _22843_/C _22843_/D VGND VGND VPWR VPWR _22844_/A sky130_fd_sc_hd__or4_4
X_25631_ _33243_/Q _24286_/X _25643_/S VGND VGND VPWR VPWR _25632_/A sky130_fd_sc_hd__mux2_1
X_34829_ _35277_/CLK _34829_/D VGND VGND VPWR VPWR _34829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_225_CLK clkbuf_6_55__f_CLK/X VGND VGND VPWR VPWR _35778_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28350_ _28350_/A VGND VGND VPWR VPWR _34498_/D sky130_fd_sc_hd__clkbuf_1
X_22774_ _20597_/X _22772_/X _22773_/X _20603_/X VGND VGND VPWR VPWR _22774_/X sky130_fd_sc_hd__a22o_1
X_25562_ _33212_/Q _24388_/X _25568_/S VGND VGND VPWR VPWR _25563_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27301_ _34002_/Q _24258_/X _27311_/S VGND VGND VPWR VPWR _27302_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24513_ _22979_/X _32750_/Q _24527_/S VGND VGND VPWR VPWR _24514_/A sky130_fd_sc_hd__mux2_1
X_21725_ _33516_/Q _33452_/Q _33388_/Q _33324_/Q _21723_/X _21724_/X VGND VGND VPWR
+ VPWR _21725_/X sky130_fd_sc_hd__mux4_2
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28281_ _28371_/S VGND VGND VPWR VPWR _28300_/S sky130_fd_sc_hd__buf_4
X_25493_ _33179_/Q _24286_/X _25505_/S VGND VGND VPWR VPWR _25494_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27232_ _27232_/A VGND VGND VPWR VPWR _33969_/D sky130_fd_sc_hd__clkbuf_1
X_24444_ _24444_/A VGND VGND VPWR VPWR _24577_/S sky130_fd_sc_hd__buf_12
XFILLER_200_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21656_ _22362_/A VGND VGND VPWR VPWR _21656_/X sky130_fd_sc_hd__buf_6
XFILLER_240_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20607_ _22557_/A VGND VGND VPWR VPWR _20607_/X sky130_fd_sc_hd__buf_4
XFILLER_205_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27163_ _27163_/A VGND VGND VPWR VPWR _33936_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24375_ _24375_/A VGND VGND VPWR VPWR _32695_/D sky130_fd_sc_hd__clkbuf_1
X_21587_ _21302_/X _21585_/X _21586_/X _21308_/X VGND VGND VPWR VPWR _21587_/X sky130_fd_sc_hd__a22o_1
XFILLER_71_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26114_ _26114_/A VGND VGND VPWR VPWR _33471_/D sky130_fd_sc_hd__clkbuf_1
X_23326_ _23326_/A VGND VGND VPWR VPWR _32226_/D sky130_fd_sc_hd__clkbuf_1
X_20538_ _18344_/X _20536_/X _20537_/X _18354_/X VGND VGND VPWR VPWR _20538_/X sky130_fd_sc_hd__a22o_1
XFILLER_181_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27094_ _26928_/X _33904_/Q _27104_/S VGND VGND VPWR VPWR _27095_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23257_ _32203_/Q _23256_/X _23268_/S VGND VGND VPWR VPWR _23258_/A sky130_fd_sc_hd__mux2_1
X_26045_ _26045_/A VGND VGND VPWR VPWR _33438_/D sky130_fd_sc_hd__clkbuf_1
X_20469_ _35850_/Q _32230_/Q _35722_/Q _35658_/Q _18289_/X _18291_/X VGND VGND VPWR
+ VPWR _20469_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22208_ _22202_/X _22207_/X _22100_/X VGND VGND VPWR VPWR _22216_/C sky130_fd_sc_hd__o21ba_1
XTAP_6600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23188_ _23188_/A VGND VGND VPWR VPWR _32176_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29804_ _29804_/A VGND VGND VPWR VPWR _35156_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22139_ _34807_/Q _34743_/Q _34679_/Q _34615_/Q _21888_/X _21889_/X VGND VGND VPWR
+ VPWR _22139_/X sky130_fd_sc_hd__mux4_1
XTAP_6644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27996_ _27996_/A VGND VGND VPWR VPWR _34330_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29735_ _35124_/Q _29169_/X _29737_/S VGND VGND VPWR VPWR _29736_/A sky130_fd_sc_hd__mux2_1
XTAP_6688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26947_ _27018_/S VGND VGND VPWR VPWR _26975_/S sky130_fd_sc_hd__buf_4
XTAP_6699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_464_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _35815_/CLK sky130_fd_sc_hd__clkbuf_16
X_16700_ _16496_/X _16698_/X _16699_/X _16499_/X VGND VGND VPWR VPWR _16700_/X sky130_fd_sc_hd__a22o_1
XFILLER_236_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29666_ _35091_/Q _29067_/X _29674_/S VGND VGND VPWR VPWR _29667_/A sky130_fd_sc_hd__mux2_1
X_17680_ _17507_/X _17678_/X _17679_/X _17512_/X VGND VGND VPWR VPWR _17680_/X sky130_fd_sc_hd__a22o_1
XTAP_5998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26878_ input10/X VGND VGND VPWR VPWR _26878_/X sky130_fd_sc_hd__buf_4
XFILLER_75_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28617_ _26981_/X _34625_/Q _28633_/S VGND VGND VPWR VPWR _28618_/A sky130_fd_sc_hd__mux2_1
XFILLER_235_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16631_ _16627_/X _16630_/X _16422_/X VGND VGND VPWR VPWR _16661_/A sky130_fd_sc_hd__o21ba_1
X_25829_ _25122_/X _33336_/Q _25843_/S VGND VGND VPWR VPWR _25830_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29597_ _29597_/A VGND VGND VPWR VPWR _35058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_216_CLK clkbuf_6_53__f_CLK/X VGND VGND VPWR VPWR _35333_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19350_ _19142_/X _19348_/X _19349_/X _19147_/X VGND VGND VPWR VPWR _19350_/X sky130_fd_sc_hd__a22o_1
X_28548_ _28548_/A VGND VGND VPWR VPWR _34592_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16562_ _33500_/Q _33436_/Q _33372_/Q _33308_/Q _16417_/X _16418_/X VGND VGND VPWR
+ VPWR _16562_/X sky130_fd_sc_hd__mux4_1
X_18301_ input80/X input79/X VGND VGND VPWR VPWR _20073_/A sky130_fd_sc_hd__nor2b_4
XFILLER_43_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19281_ _33512_/Q _33448_/Q _33384_/Q _33320_/Q _19070_/X _19071_/X VGND VGND VPWR
+ VPWR _19281_/X sky130_fd_sc_hd__mux4_1
X_28479_ _28506_/S VGND VGND VPWR VPWR _28498_/S sky130_fd_sc_hd__buf_6
X_16493_ _34266_/Q _34202_/Q _34138_/Q _34074_/Q _16383_/X _16384_/X VGND VGND VPWR
+ VPWR _16493_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18232_ _35596_/Q _35532_/Q _35468_/Q _35404_/Q _17956_/X _17957_/X VGND VGND VPWR
+ VPWR _18232_/X sky130_fd_sc_hd__mux4_1
X_30510_ _30510_/A VGND VGND VPWR VPWR _35490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31490_ _31490_/A VGND VGND VPWR VPWR _35955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18163_ _33290_/Q _36170_/Q _33162_/Q _33098_/Q _16028_/X _17157_/A VGND VGND VPWR
+ VPWR _18163_/X sky130_fd_sc_hd__mux4_1
X_30441_ _23310_/X _35458_/Q _30455_/S VGND VGND VPWR VPWR _30442_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17114_ _34539_/Q _32427_/Q _34411_/Q _34347_/Q _16872_/X _16873_/X VGND VGND VPWR
+ VPWR _17114_/X sky130_fd_sc_hd__mux4_1
X_33160_ _35909_/CLK _33160_/D VGND VGND VPWR VPWR _33160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18094_ _18094_/A VGND VGND VPWR VPWR _32007_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_141_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30372_ _30372_/A VGND VGND VPWR VPWR _35425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_209_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32111_ _35552_/CLK _32111_/D VGND VGND VPWR VPWR _32111_/Q sky130_fd_sc_hd__dfxtp_1
X_17045_ _17041_/X _17044_/X _16808_/X VGND VGND VPWR VPWR _17046_/D sky130_fd_sc_hd__o21ba_1
X_33091_ _33922_/CLK _33091_/D VGND VGND VPWR VPWR _33091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32042_ _36075_/CLK _32042_/D VGND VGND VPWR VPWR _32042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ _34272_/Q _34208_/Q _34144_/Q _34080_/Q _18683_/X _18684_/X VGND VGND VPWR
+ VPWR _18996_/X sky130_fd_sc_hd__mux4_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35801_ _35801_/CLK _35801_/D VGND VGND VPWR VPWR _35801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17947_ _33283_/Q _36163_/Q _33155_/Q _33091_/Q _17764_/X _17765_/X VGND VGND VPWR
+ VPWR _17947_/X sky130_fd_sc_hd__mux4_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33993_ _34817_/CLK _33993_/D VGND VGND VPWR VPWR _33993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_455_CLK clkbuf_6_11__f_CLK/X VGND VGND VPWR VPWR _35303_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_239_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35732_ _35733_/CLK _35732_/D VGND VGND VPWR VPWR _35732_/Q sky130_fd_sc_hd__dfxtp_1
X_32944_ _33009_/CLK _32944_/D VGND VGND VPWR VPWR _32944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17878_ _32769_/Q _32705_/Q _32641_/Q _36097_/Q _17625_/X _17762_/X VGND VGND VPWR
+ VPWR _17878_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19617_ _19294_/X _19615_/X _19616_/X _19297_/X VGND VGND VPWR VPWR _19617_/X sky130_fd_sc_hd__a22o_1
X_16829_ _35555_/Q _35491_/Q _35427_/Q _35363_/Q _16544_/X _16545_/X VGND VGND VPWR
+ VPWR _16829_/X sky130_fd_sc_hd__mux4_1
X_35663_ _35792_/CLK _35663_/D VGND VGND VPWR VPWR _35663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32875_ _36075_/CLK _32875_/D VGND VGND VPWR VPWR _32875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_207_CLK clkbuf_6_52__f_CLK/X VGND VGND VPWR VPWR _35975_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31826_ _31826_/A VGND VGND VPWR VPWR _36114_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19548_ _35759_/Q _35119_/Q _34479_/Q _33839_/Q _19440_/X _19441_/X VGND VGND VPWR
+ VPWR _19548_/X sky130_fd_sc_hd__mux4_1
X_34614_ _34745_/CLK _34614_/D VGND VGND VPWR VPWR _34614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35594_ _35852_/CLK _35594_/D VGND VGND VPWR VPWR _35594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34545_ _34866_/CLK _34545_/D VGND VGND VPWR VPWR _34545_/Q sky130_fd_sc_hd__dfxtp_1
X_19479_ _35821_/Q _32198_/Q _35693_/Q _35629_/Q _19260_/X _19261_/X VGND VGND VPWR
+ VPWR _19479_/X sky130_fd_sc_hd__mux4_1
X_31757_ _36082_/Q input30/X _31763_/S VGND VGND VPWR VPWR _31758_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21510_ _21510_/A _21510_/B _21510_/C _21510_/D VGND VGND VPWR VPWR _21511_/A sky130_fd_sc_hd__or4_4
X_30708_ _30708_/A VGND VGND VPWR VPWR _35584_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22490_ _22305_/X _22488_/X _22489_/X _22308_/X VGND VGND VPWR VPWR _22490_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34476_ _35885_/CLK _34476_/D VGND VGND VPWR VPWR _34476_/Q sky130_fd_sc_hd__dfxtp_1
X_31688_ _36049_/Q input34/X _31700_/S VGND VGND VPWR VPWR _31689_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33427_ _36237_/CLK _33427_/D VGND VGND VPWR VPWR _33427_/Q sky130_fd_sc_hd__dfxtp_1
X_36215_ _36220_/CLK _36215_/D VGND VGND VPWR VPWR _36215_/Q sky130_fd_sc_hd__dfxtp_1
X_21441_ _21441_/A VGND VGND VPWR VPWR _36195_/D sky130_fd_sc_hd__clkbuf_1
X_30639_ _35552_/Q _29107_/X _30641_/S VGND VGND VPWR VPWR _30640_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_954 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36146_ _36146_/CLK _36146_/D VGND VGND VPWR VPWR _36146_/Q sky130_fd_sc_hd__dfxtp_1
X_24160_ _24160_/A VGND VGND VPWR VPWR _32613_/D sky130_fd_sc_hd__clkbuf_1
X_33358_ _33490_/CLK _33358_/D VGND VGND VPWR VPWR _33358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21372_ _33506_/Q _33442_/Q _33378_/Q _33314_/Q _21370_/X _21371_/X VGND VGND VPWR
+ VPWR _21372_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23111_ input63/X VGND VGND VPWR VPWR _23111_/X sky130_fd_sc_hd__buf_4
X_20323_ _33221_/Q _32581_/Q _35973_/Q _35909_/Q _20080_/X _20081_/X VGND VGND VPWR
+ VPWR _20323_/X sky130_fd_sc_hd__mux4_1
X_32309_ _35956_/CLK _32309_/D VGND VGND VPWR VPWR _32309_/Q sky130_fd_sc_hd__dfxtp_1
X_24091_ _24091_/A VGND VGND VPWR VPWR _32581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36077_ _36077_/CLK _36077_/D VGND VGND VPWR VPWR _36077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33289_ _36169_/CLK _33289_/D VGND VGND VPWR VPWR _33289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23042_ _23041_/X _32066_/Q _23063_/S VGND VGND VPWR VPWR _23043_/A sky130_fd_sc_hd__mux2_1
X_35028_ _35028_/CLK _35028_/D VGND VGND VPWR VPWR _35028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20254_ _35779_/Q _35139_/Q _34499_/Q _33859_/Q _20146_/X _20147_/X VGND VGND VPWR
+ VPWR _20254_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27850_ _27850_/A VGND VGND VPWR VPWR _34261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20185_ _35841_/Q _32220_/Q _35713_/Q _35649_/Q _19966_/X _19967_/X VGND VGND VPWR
+ VPWR _20185_/X sky130_fd_sc_hd__mux4_1
XTAP_5206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26801_ _33796_/Q _24413_/X _26811_/S VGND VGND VPWR VPWR _26802_/A sky130_fd_sc_hd__mux2_1
XTAP_5228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27781_ _34229_/Q _24366_/X _27781_/S VGND VGND VPWR VPWR _27782_/A sky130_fd_sc_hd__mux2_1
X_24993_ _24989_/X _32974_/Q _25020_/S VGND VGND VPWR VPWR _24994_/A sky130_fd_sc_hd__mux2_1
XTAP_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29520_ _29652_/S VGND VGND VPWR VPWR _29539_/S sky130_fd_sc_hd__buf_4
XTAP_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_446_CLK clkbuf_leaf_50_CLK/A VGND VGND VPWR VPWR _36067_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_218_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26732_ _33763_/Q _24311_/X _26748_/S VGND VGND VPWR VPWR _26733_/A sky130_fd_sc_hd__mux2_1
X_23944_ _23034_/X _32512_/Q _23962_/S VGND VGND VPWR VPWR _23945_/A sky130_fd_sc_hd__mux2_1
XTAP_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29451_ _23241_/X _34989_/Q _29467_/S VGND VGND VPWR VPWR _29452_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26663_ _25156_/X _33731_/Q _26675_/S VGND VGND VPWR VPWR _26664_/A sky130_fd_sc_hd__mux2_1
XTAP_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_804 _22892_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23875_ _23875_/A VGND VGND VPWR VPWR _32479_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_815 _22923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28402_ _26863_/X _34523_/Q _28414_/S VGND VGND VPWR VPWR _28403_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25614_ _33235_/Q _24261_/X _25622_/S VGND VGND VPWR VPWR _25615_/A sky130_fd_sc_hd__mux2_1
XANTENNA_826 _23121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29382_ _23345_/X _34957_/Q _29382_/S VGND VGND VPWR VPWR _29383_/A sky130_fd_sc_hd__mux2_1
X_22826_ _33036_/Q _32972_/Q _32908_/Q _32844_/Q _20580_/X _20583_/X VGND VGND VPWR
+ VPWR _22826_/X sky130_fd_sc_hd__mux4_1
XANTENNA_837 _23280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26594_ _25053_/X _33698_/Q _26612_/S VGND VGND VPWR VPWR _26595_/A sky130_fd_sc_hd__mux2_1
XANTENNA_848 _23970_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_859 _24354_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28333_ _28333_/A VGND VGND VPWR VPWR _34490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_871 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25545_ _33204_/Q _24363_/X _25547_/S VGND VGND VPWR VPWR _25546_/A sky130_fd_sc_hd__mux2_1
X_22757_ _22501_/X _22755_/X _22756_/X _22506_/X VGND VGND VPWR VPWR _22757_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_1243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21708_ _33195_/Q _32555_/Q _35947_/Q _35883_/Q _21674_/X _21675_/X VGND VGND VPWR
+ VPWR _21708_/X sky130_fd_sc_hd__mux4_1
X_28264_ _28264_/A VGND VGND VPWR VPWR _34457_/D sky130_fd_sc_hd__clkbuf_1
X_22688_ _22455_/X _22686_/X _22687_/X _22458_/X VGND VGND VPWR VPWR _22688_/X sky130_fd_sc_hd__a22o_1
XFILLER_200_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25476_ _33171_/Q _24261_/X _25484_/S VGND VGND VPWR VPWR _25477_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27215_ _27215_/A VGND VGND VPWR VPWR _33961_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24427_ _24427_/A VGND VGND VPWR VPWR _32712_/D sky130_fd_sc_hd__clkbuf_1
X_21639_ _34793_/Q _34729_/Q _34665_/Q _34601_/Q _21535_/X _21536_/X VGND VGND VPWR
+ VPWR _21639_/X sky130_fd_sc_hd__mux4_1
X_28195_ _26956_/X _34425_/Q _28207_/S VGND VGND VPWR VPWR _28196_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27146_ _27005_/X _33929_/Q _27146_/S VGND VGND VPWR VPWR _27147_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24358_ _32690_/Q _24357_/X _24367_/S VGND VGND VPWR VPWR _24359_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23309_ _23309_/A VGND VGND VPWR VPWR _32220_/D sky130_fd_sc_hd__clkbuf_1
X_24289_ input6/X VGND VGND VPWR VPWR _24289_/X sky130_fd_sc_hd__buf_4
X_27077_ _26903_/X _33896_/Q _27083_/S VGND VGND VPWR VPWR _27078_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26028_ _26028_/A VGND VGND VPWR VPWR _33430_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_32__f_CLK clkbuf_5_16_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_32__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_153_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1203 _23105_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18850_ _34779_/Q _34715_/Q _34651_/Q _34587_/Q _18529_/X _18530_/X VGND VGND VPWR
+ VPWR _18850_/X sky130_fd_sc_hd__mux4_1
XTAP_6430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1214 _23327_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1225 _24345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17801_ _17555_/X _17799_/X _17800_/X _17558_/X VGND VGND VPWR VPWR _17801_/X sky130_fd_sc_hd__a22o_1
XANTENNA_1236 _25013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1247 _26547_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18781_ _35289_/Q _35225_/Q _35161_/Q _32281_/Q _18600_/X _18601_/X VGND VGND VPWR
+ VPWR _18781_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1258 _27646_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15993_ _15977_/X _15984_/X _15987_/X _15992_/X VGND VGND VPWR VPWR _15993_/X sky130_fd_sc_hd__a22o_1
XFILLER_212_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1269 _30327_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27979_ _27979_/A VGND VGND VPWR VPWR _34322_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_437_CLK clkbuf_leaf_61_CLK/A VGND VGND VPWR VPWR _34087_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_5762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17732_ _33277_/Q _36157_/Q _33149_/Q _33085_/Q _17411_/X _17412_/X VGND VGND VPWR
+ VPWR _17732_/X sky130_fd_sc_hd__mux4_1
X_29718_ _29787_/S VGND VGND VPWR VPWR _29737_/S sky130_fd_sc_hd__buf_4
XTAP_5773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30990_ _30990_/A VGND VGND VPWR VPWR _35718_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29649_ _29649_/A VGND VGND VPWR VPWR _35083_/D sky130_fd_sc_hd__clkbuf_1
X_17663_ _33019_/Q _32955_/Q _32891_/Q _32827_/Q _17342_/X _17343_/X VGND VGND VPWR
+ VPWR _17663_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19402_ _19363_/X _19400_/X _19401_/X _19367_/X VGND VGND VPWR VPWR _19402_/X sky130_fd_sc_hd__a22o_1
XFILLER_236_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16614_ _16293_/X _16612_/X _16613_/X _16296_/X VGND VGND VPWR VPWR _16614_/X sky130_fd_sc_hd__a22o_1
X_32660_ _36116_/CLK _32660_/D VGND VGND VPWR VPWR _32660_/Q sky130_fd_sc_hd__dfxtp_1
X_17594_ _33273_/Q _36153_/Q _33145_/Q _33081_/Q _17411_/X _17412_/X VGND VGND VPWR
+ VPWR _17594_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19333_ _35753_/Q _35113_/Q _34473_/Q _33833_/Q _19087_/X _19088_/X VGND VGND VPWR
+ VPWR _19333_/X sky130_fd_sc_hd__mux4_1
X_31611_ _31611_/A VGND VGND VPWR VPWR _36012_/D sky130_fd_sc_hd__clkbuf_1
X_16545_ _17957_/A VGND VGND VPWR VPWR _16545_/X sky130_fd_sc_hd__clkbuf_4
X_32591_ _36048_/CLK _32591_/D VGND VGND VPWR VPWR _32591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34330_ _34970_/CLK _34330_/D VGND VGND VPWR VPWR _34330_/Q sky130_fd_sc_hd__dfxtp_1
X_31542_ _31542_/A VGND VGND VPWR VPWR _35980_/D sky130_fd_sc_hd__clkbuf_1
X_19264_ _18941_/X _19262_/X _19263_/X _18944_/X VGND VGND VPWR VPWR _19264_/X sky130_fd_sc_hd__a22o_1
XFILLER_204_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16476_ _35545_/Q _35481_/Q _35417_/Q _35353_/Q _16191_/X _16192_/X VGND VGND VPWR
+ VPWR _16476_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18215_ _33804_/Q _33740_/Q _33676_/Q _33612_/Q _16020_/X _16021_/X VGND VGND VPWR
+ VPWR _18215_/X sky130_fd_sc_hd__mux4_1
X_34261_ _34262_/CLK _34261_/D VGND VGND VPWR VPWR _34261_/Q sky130_fd_sc_hd__dfxtp_1
X_31473_ _31473_/A VGND VGND VPWR VPWR _35947_/D sky130_fd_sc_hd__clkbuf_1
X_19195_ _35749_/Q _35109_/Q _34469_/Q _33829_/Q _19087_/X _19088_/X VGND VGND VPWR
+ VPWR _19195_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36000_ _36001_/CLK _36000_/D VGND VGND VPWR VPWR _36000_/Q sky130_fd_sc_hd__dfxtp_1
X_33212_ _36028_/CLK _33212_/D VGND VGND VPWR VPWR _33212_/Q sky130_fd_sc_hd__dfxtp_1
X_18146_ _34825_/Q _34761_/Q _34697_/Q _34633_/Q _17994_/X _17995_/X VGND VGND VPWR
+ VPWR _18146_/X sky130_fd_sc_hd__mux4_1
X_30424_ _23283_/X _35450_/Q _30434_/S VGND VGND VPWR VPWR _30425_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34192_ _34259_/CLK _34192_/D VGND VGND VPWR VPWR _34192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33143_ _36087_/CLK _33143_/D VGND VGND VPWR VPWR _33143_/Q sky130_fd_sc_hd__dfxtp_1
X_18077_ _17769_/X _18075_/X _18076_/X _17773_/X VGND VGND VPWR VPWR _18077_/X sky130_fd_sc_hd__a22o_1
X_30355_ _23121_/X _35417_/Q _30371_/S VGND VGND VPWR VPWR _30356_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17028_ _32489_/Q _32361_/Q _32041_/Q _36009_/Q _16923_/X _16711_/X VGND VGND VPWR
+ VPWR _17028_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33074_ _33520_/CLK _33074_/D VGND VGND VPWR VPWR _33074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30286_ _35385_/Q _29185_/X _30298_/S VGND VGND VPWR VPWR _30287_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32025_ _35995_/CLK _32025_/D VGND VGND VPWR VPWR _32025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ _35807_/Q _32183_/Q _35679_/Q _35615_/Q _18907_/X _18908_/X VGND VGND VPWR
+ VPWR _18979_/X sky130_fd_sc_hd__mux4_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_428_CLK clkbuf_6_36__f_CLK/X VGND VGND VPWR VPWR _36136_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21990_ _21952_/X _21988_/X _21989_/X _21955_/X VGND VGND VPWR VPWR _21990_/X sky130_fd_sc_hd__a22o_1
XFILLER_230_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33976_ _36152_/CLK _33976_/D VGND VGND VPWR VPWR _33976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35715_ _35715_/CLK _35715_/D VGND VGND VPWR VPWR _35715_/Q sky130_fd_sc_hd__dfxtp_1
X_20941_ _20941_/A VGND VGND VPWR VPWR _36181_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32927_ _36065_/CLK _32927_/D VGND VGND VPWR VPWR _32927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20872_ _33748_/Q _33684_/Q _33620_/Q _33556_/Q _20737_/X _20738_/X VGND VGND VPWR
+ VPWR _20872_/X sky130_fd_sc_hd__mux4_1
X_35646_ _35710_/CLK _35646_/D VGND VGND VPWR VPWR _35646_/Q sky130_fd_sc_hd__dfxtp_1
X_23660_ _23660_/A VGND VGND VPWR VPWR _32379_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32858_ _32860_/CLK _32858_/D VGND VGND VPWR VPWR _32858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22611_ _22607_/X _22610_/X _22434_/X VGND VGND VPWR VPWR _22633_/A sky130_fd_sc_hd__o21ba_2
XFILLER_41_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31809_ _36107_/Q input58/X _31813_/S VGND VGND VPWR VPWR _31810_/A sky130_fd_sc_hd__mux2_1
X_23591_ _23591_/A VGND VGND VPWR VPWR _32346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32789_ _32983_/CLK _32789_/D VGND VGND VPWR VPWR _32789_/Q sky130_fd_sc_hd__dfxtp_1
X_35577_ _35577_/CLK _35577_/D VGND VGND VPWR VPWR _35577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22542_ _33539_/Q _33475_/Q _33411_/Q _33347_/Q _22429_/X _22430_/X VGND VGND VPWR
+ VPWR _22542_/X sky130_fd_sc_hd__mux4_1
X_25330_ _25330_/A VGND VGND VPWR VPWR _33103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34528_ _35039_/CLK _34528_/D VGND VGND VPWR VPWR _34528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22473_ _22148_/X _22471_/X _22472_/X _22153_/X VGND VGND VPWR VPWR _22473_/X sky130_fd_sc_hd__a22o_1
X_25261_ _25261_/A VGND VGND VPWR VPWR _33071_/D sky130_fd_sc_hd__clkbuf_1
X_34459_ _35098_/CLK _34459_/D VGND VGND VPWR VPWR _34459_/Q sky130_fd_sc_hd__dfxtp_1
X_27000_ _26999_/X _33863_/Q _27006_/S VGND VGND VPWR VPWR _27001_/A sky130_fd_sc_hd__mux2_1
X_24212_ _24212_/A VGND VGND VPWR VPWR _32638_/D sky130_fd_sc_hd__clkbuf_1
X_21424_ _21310_/X _21422_/X _21423_/X _21314_/X VGND VGND VPWR VPWR _21424_/X sky130_fd_sc_hd__a22o_1
X_25192_ _25192_/A VGND VGND VPWR VPWR _33038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24143_ _24143_/A VGND VGND VPWR VPWR _32605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21355_ _33185_/Q _32545_/Q _35937_/Q _35873_/Q _21321_/X _21322_/X VGND VGND VPWR
+ VPWR _21355_/X sky130_fd_sc_hd__mux4_1
X_36129_ _36129_/CLK _36129_/D VGND VGND VPWR VPWR _36129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20306_ _34309_/Q _34245_/Q _34181_/Q _34117_/Q _20095_/X _20096_/X VGND VGND VPWR
+ VPWR _20306_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24074_ _24074_/A VGND VGND VPWR VPWR _32573_/D sky130_fd_sc_hd__clkbuf_1
X_28951_ _28951_/A VGND VGND VPWR VPWR _34783_/D sky130_fd_sc_hd__clkbuf_1
X_21286_ _34783_/Q _34719_/Q _34655_/Q _34591_/Q _21182_/X _21183_/X VGND VGND VPWR
+ VPWR _21286_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_1211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23025_ input42/X VGND VGND VPWR VPWR _23025_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27902_ _34286_/Q _24345_/X _27916_/S VGND VGND VPWR VPWR _27903_/A sky130_fd_sc_hd__mux2_1
X_20237_ _20237_/A _20237_/B _20237_/C _20237_/D VGND VGND VPWR VPWR _20238_/A sky130_fd_sc_hd__or4_4
X_28882_ _26974_/X _34751_/Q _28882_/S VGND VGND VPWR VPWR _28883_/A sky130_fd_sc_hd__mux2_1
XTAP_5003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27833_ _27833_/A _31140_/B VGND VGND VPWR VPWR _27966_/S sky130_fd_sc_hd__nor2_8
XTAP_5025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20168_ _20159_/X _20166_/X _20167_/X VGND VGND VPWR VPWR _20169_/D sky130_fd_sc_hd__o21ba_1
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_419_CLK clkbuf_6_38__f_CLK/X VGND VGND VPWR VPWR _34805_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_5069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27764_ _27764_/A VGND VGND VPWR VPWR _34220_/D sky130_fd_sc_hd__clkbuf_1
X_24976_ _24976_/A VGND VGND VPWR VPWR _32967_/D sky130_fd_sc_hd__clkbuf_1
X_20099_ _33535_/Q _33471_/Q _33407_/Q _33343_/Q _19776_/X _19777_/X VGND VGND VPWR
+ VPWR _20099_/X sky130_fd_sc_hd__mux4_1
XTAP_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29503_ _23322_/X _35014_/Q _29509_/S VGND VGND VPWR VPWR _29504_/A sky130_fd_sc_hd__mux2_1
XTAP_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26715_ _33755_/Q _24286_/X _26727_/S VGND VGND VPWR VPWR _26716_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23927_ _23010_/X _32504_/Q _23941_/S VGND VGND VPWR VPWR _23928_/A sky130_fd_sc_hd__mux2_1
X_27695_ _27695_/A VGND VGND VPWR VPWR _34188_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_601 _20167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_612 _18505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29434_ _23199_/X _34981_/Q _29446_/S VGND VGND VPWR VPWR _29435_/A sky130_fd_sc_hd__mux2_1
XFILLER_233_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26646_ _25131_/X _33723_/Q _26654_/S VGND VGND VPWR VPWR _26647_/A sky130_fd_sc_hd__mux2_1
XTAP_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_623 _18609_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23858_ _23858_/A VGND VGND VPWR VPWR _32471_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_634 _19065_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_645 _19428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_656 _20334_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22809_ _34571_/Q _32459_/Q _34443_/Q _34379_/Q _22531_/X _22532_/X VGND VGND VPWR
+ VPWR _22809_/X sky130_fd_sc_hd__mux4_1
X_29365_ _29365_/A VGND VGND VPWR VPWR _34948_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_667 _22460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_678 _22556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26577_ _25029_/X _33690_/Q _26591_/S VGND VGND VPWR VPWR _26578_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23789_ _23007_/X _32439_/Q _23805_/S VGND VGND VPWR VPWR _23790_/A sky130_fd_sc_hd__mux2_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_689 _22442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16330_ _33173_/Q _32533_/Q _35925_/Q _35861_/Q _16063_/X _16065_/X VGND VGND VPWR
+ VPWR _16330_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28316_ _28316_/A VGND VGND VPWR VPWR _34482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25528_ _25597_/S VGND VGND VPWR VPWR _25547_/S sky130_fd_sc_hd__buf_6
XFILLER_129_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29296_ _29296_/A VGND VGND VPWR VPWR _34915_/D sky130_fd_sc_hd__clkbuf_1
X_28247_ _28247_/A VGND VGND VPWR VPWR _34449_/D sky130_fd_sc_hd__clkbuf_1
X_16261_ _16056_/X _16259_/X _16260_/X _16068_/X VGND VGND VPWR VPWR _16261_/X sky130_fd_sc_hd__a22o_1
XFILLER_185_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25459_ _25459_/A VGND VGND VPWR VPWR _33165_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18000_ _35076_/Q _35012_/Q _34948_/Q _34884_/Q _17862_/X _17863_/X VGND VGND VPWR
+ VPWR _18000_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16192_ _17847_/A VGND VGND VPWR VPWR _16192_/X sky130_fd_sc_hd__buf_4
X_28178_ _26931_/X _34417_/Q _28186_/S VGND VGND VPWR VPWR _28179_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27129_ _27129_/A VGND VGND VPWR VPWR _33920_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30140_ _35316_/Q _29169_/X _30142_/S VGND VGND VPWR VPWR _30141_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19951_ _19951_/A VGND VGND VPWR VPWR _32122_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18902_ _18649_/X _18900_/X _18901_/X _18655_/X VGND VGND VPWR VPWR _18902_/X sky130_fd_sc_hd__a22o_1
X_30071_ _35283_/Q _29067_/X _30079_/S VGND VGND VPWR VPWR _30072_/A sky130_fd_sc_hd__mux2_1
XANTENNA_1000 _17957_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19882_ _19807_/X _19880_/X _19881_/X _19812_/X VGND VGND VPWR VPWR _19882_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1011 _17908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1022 _17865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1033 _17853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18833_ _18829_/X _18832_/X _18722_/X VGND VGND VPWR VPWR _18857_/A sky130_fd_sc_hd__o21ba_1
XANTENNA_1044 _17159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1055 _16205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1066 _17064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1077 _17164_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18764_ _18443_/X _18762_/X _18763_/X _18446_/X VGND VGND VPWR VPWR _18764_/X sky130_fd_sc_hd__a22o_1
X_33830_ _35942_/CLK _33830_/D VGND VGND VPWR VPWR _33830_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1088 _17232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15976_ _17761_/A VGND VGND VPWR VPWR _17855_/A sky130_fd_sc_hd__buf_12
XANTENNA_1099 _17368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17715_ _17502_/X _17711_/X _17714_/X _17505_/X VGND VGND VPWR VPWR _17715_/X sky130_fd_sc_hd__a22o_1
X_33761_ _36123_/CLK _33761_/D VGND VGND VPWR VPWR _33761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30973_ _30973_/A VGND VGND VPWR VPWR _35710_/D sky130_fd_sc_hd__clkbuf_1
X_18695_ _32983_/Q _32919_/Q _32855_/Q _32791_/Q _18583_/X _18584_/X VGND VGND VPWR
+ VPWR _18695_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_1378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35500_ _35500_/CLK _35500_/D VGND VGND VPWR VPWR _35500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32712_ _36168_/CLK _32712_/D VGND VGND VPWR VPWR _32712_/Q sky130_fd_sc_hd__dfxtp_1
X_17646_ _34554_/Q _32442_/Q _34426_/Q _34362_/Q _17578_/X _17579_/X VGND VGND VPWR
+ VPWR _17646_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33692_ _33692_/CLK _33692_/D VGND VGND VPWR VPWR _33692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32643_ _33026_/CLK _32643_/D VGND VGND VPWR VPWR _32643_/Q sky130_fd_sc_hd__dfxtp_1
X_35431_ _35750_/CLK _35431_/D VGND VGND VPWR VPWR _35431_/Q sky130_fd_sc_hd__dfxtp_1
X_17577_ _17502_/X _17575_/X _17576_/X _17505_/X VGND VGND VPWR VPWR _17577_/X sky130_fd_sc_hd__a22o_1
XFILLER_1_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19316_ _33769_/Q _33705_/Q _33641_/Q _33577_/Q _19143_/X _19144_/X VGND VGND VPWR
+ VPWR _19316_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16528_ _34267_/Q _34203_/Q _34139_/Q _34075_/Q _16383_/X _16384_/X VGND VGND VPWR
+ VPWR _16528_/X sky130_fd_sc_hd__mux4_1
X_35362_ _35940_/CLK _35362_/D VGND VGND VPWR VPWR _35362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32574_ _35968_/CLK _32574_/D VGND VGND VPWR VPWR _32574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34313_ _36103_/CLK _34313_/D VGND VGND VPWR VPWR _34313_/Q sky130_fd_sc_hd__dfxtp_1
X_31525_ _23316_/X _35972_/Q _31535_/S VGND VGND VPWR VPWR _31526_/A sky130_fd_sc_hd__mux2_1
X_19247_ _34279_/Q _34215_/Q _34151_/Q _34087_/Q _19036_/X _19037_/X VGND VGND VPWR
+ VPWR _19247_/X sky130_fd_sc_hd__mux4_1
X_16459_ _33753_/Q _33689_/Q _33625_/Q _33561_/Q _16137_/X _16138_/X VGND VGND VPWR
+ VPWR _16459_/X sky130_fd_sc_hd__mux4_1
X_35293_ _35293_/CLK _35293_/D VGND VGND VPWR VPWR _35293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34244_ _34310_/CLK _34244_/D VGND VGND VPWR VPWR _34244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31456_ _23152_/X _35939_/Q _31472_/S VGND VGND VPWR VPWR _31457_/A sky130_fd_sc_hd__mux2_1
X_19178_ _19178_/A _19178_/B _19178_/C _19178_/D VGND VGND VPWR VPWR _19179_/A sky130_fd_sc_hd__or4_4
XFILLER_191_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18129_ _34057_/Q _33993_/Q _33929_/Q _32265_/Q _16058_/X _16060_/X VGND VGND VPWR
+ VPWR _18129_/X sky130_fd_sc_hd__mux4_1
X_30407_ _23256_/X _35442_/Q _30413_/S VGND VGND VPWR VPWR _30408_/A sky130_fd_sc_hd__mux2_1
X_34175_ _36161_/CLK _34175_/D VGND VGND VPWR VPWR _34175_/Q sky130_fd_sc_hd__dfxtp_1
X_31387_ _31387_/A VGND VGND VPWR VPWR _35906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21140_ _21136_/X _21139_/X _21030_/X _21031_/X VGND VGND VPWR VPWR _21157_/B sky130_fd_sc_hd__o211a_1
X_33126_ _36135_/CLK _33126_/D VGND VGND VPWR VPWR _33126_/Q sky130_fd_sc_hd__dfxtp_1
X_30338_ _23096_/X _35409_/Q _30350_/S VGND VGND VPWR VPWR _30339_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21071_ _20957_/X _21069_/X _21070_/X _20961_/X VGND VGND VPWR VPWR _21071_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33057_ _36130_/CLK _33057_/D VGND VGND VPWR VPWR _33057_/Q sky130_fd_sc_hd__dfxtp_1
X_30269_ _35377_/Q _29160_/X _30277_/S VGND VGND VPWR VPWR _30270_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20022_ _33789_/Q _33725_/Q _33661_/Q _33597_/Q _19849_/X _19850_/X VGND VGND VPWR
+ VPWR _20022_/X sky130_fd_sc_hd__mux4_1
X_32008_ _36185_/CLK _32008_/D VGND VGND VPWR VPWR _32008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24830_ _23041_/X _32898_/Q _24844_/S VGND VGND VPWR VPWR _24831_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24761_ _24761_/A VGND VGND VPWR VPWR _32865_/D sky130_fd_sc_hd__clkbuf_1
X_33959_ _34087_/CLK _33959_/D VGND VGND VPWR VPWR _33959_/Q sky130_fd_sc_hd__dfxtp_1
X_21973_ _22446_/A VGND VGND VPWR VPWR _21973_/X sky130_fd_sc_hd__buf_4
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26500_ _25115_/X _33654_/Q _26518_/S VGND VGND VPWR VPWR _26501_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23712_ _23712_/A VGND VGND VPWR VPWR _32402_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20924_ _20626_/X _20922_/X _20923_/X _20637_/X VGND VGND VPWR VPWR _20924_/X sky130_fd_sc_hd__a22o_1
X_27480_ _26900_/X _34087_/Q _27488_/S VGND VGND VPWR VPWR _27481_/A sky130_fd_sc_hd__mux2_1
X_24692_ _24692_/A VGND VGND VPWR VPWR _32833_/D sky130_fd_sc_hd__clkbuf_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26431_ _26431_/A VGND VGND VPWR VPWR _33621_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20855_ _22396_/A VGND VGND VPWR VPWR _20855_/X sky130_fd_sc_hd__buf_4
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35629_ _35949_/CLK _35629_/D VGND VGND VPWR VPWR _35629_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23643_ _23643_/A VGND VGND VPWR VPWR _32371_/D sky130_fd_sc_hd__clkbuf_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29150_ _29150_/A VGND VGND VPWR VPWR _34861_/D sky130_fd_sc_hd__clkbuf_1
X_26362_ _25112_/X _33589_/Q _26362_/S VGND VGND VPWR VPWR _26363_/A sky130_fd_sc_hd__mux2_1
X_20786_ _20626_/X _20784_/X _20785_/X _20637_/X VGND VGND VPWR VPWR _20786_/X sky130_fd_sc_hd__a22o_1
X_23574_ _23574_/A VGND VGND VPWR VPWR _32338_/D sky130_fd_sc_hd__clkbuf_1
X_28101_ _27017_/X _34381_/Q _28101_/S VGND VGND VPWR VPWR _28102_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25313_ _25313_/A VGND VGND VPWR VPWR _33096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22525_ _33218_/Q _32578_/Q _35970_/Q _35906_/Q _22380_/X _22381_/X VGND VGND VPWR
+ VPWR _22525_/X sky130_fd_sc_hd__mux4_1
X_29081_ _29081_/A VGND VGND VPWR VPWR _34839_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26293_ _25010_/X _33556_/Q _26299_/S VGND VGND VPWR VPWR _26294_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28032_ _28101_/S VGND VGND VPWR VPWR _28051_/S sky130_fd_sc_hd__buf_6
XFILLER_183_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25244_ _25244_/A VGND VGND VPWR VPWR _33063_/D sky130_fd_sc_hd__clkbuf_1
X_22456_ _34816_/Q _34752_/Q _34688_/Q _34624_/Q _22241_/X _22242_/X VGND VGND VPWR
+ VPWR _22456_/X sky130_fd_sc_hd__mux4_1
XFILLER_183_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21407_ _21401_/X _21402_/X _21405_/X _21406_/X VGND VGND VPWR VPWR _21407_/X sky130_fd_sc_hd__a22o_1
X_25175_ _25174_/X _33033_/Q _25175_/S VGND VGND VPWR VPWR _25176_/A sky130_fd_sc_hd__mux2_1
X_22387_ _22102_/X _22385_/X _22386_/X _22105_/X VGND VGND VPWR VPWR _22387_/X sky130_fd_sc_hd__a22o_1
X_24126_ _24126_/A VGND VGND VPWR VPWR _32597_/D sky130_fd_sc_hd__clkbuf_1
X_21338_ _34273_/Q _34209_/Q _34145_/Q _34081_/Q _21336_/X _21337_/X VGND VGND VPWR
+ VPWR _21338_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29983_ _29983_/A VGND VGND VPWR VPWR _35241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28934_ _28934_/A VGND VGND VPWR VPWR _34775_/D sky130_fd_sc_hd__clkbuf_1
X_24057_ _24057_/A VGND VGND VPWR VPWR _32565_/D sky130_fd_sc_hd__clkbuf_1
X_21269_ _34015_/Q _33951_/Q _33887_/Q _32159_/Q _21267_/X _21268_/X VGND VGND VPWR
+ VPWR _21269_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23008_ _23007_/X _32055_/Q _23032_/S VGND VGND VPWR VPWR _23009_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28865_ _28865_/A VGND VGND VPWR VPWR _34742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27816_ _27816_/A VGND VGND VPWR VPWR _34245_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28796_ _26847_/X _34710_/Q _28798_/S VGND VGND VPWR VPWR _28797_/A sky130_fd_sc_hd__mux2_1
XTAP_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27747_ _27747_/A VGND VGND VPWR VPWR _34212_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24959_ _24959_/A VGND VGND VPWR VPWR _32959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _17853_/A VGND VGND VPWR VPWR _17500_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ _18476_/X _18479_/X _18311_/X VGND VGND VPWR VPWR _18504_/A sky130_fd_sc_hd__o21ba_1
XTAP_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27678_ _34180_/Q _24413_/X _27688_/S VGND VGND VPWR VPWR _27679_/A sky130_fd_sc_hd__mux2_1
XTAP_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_420 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_431 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29417_ _23133_/X _34973_/Q _29425_/S VGND VGND VPWR VPWR _29418_/A sky130_fd_sc_hd__mux2_1
X_17431_ _17425_/X _17430_/X _17147_/X VGND VGND VPWR VPWR _17439_/C sky130_fd_sc_hd__o21ba_1
XANTENNA_442 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26629_ _25106_/X _33715_/Q _26633_/S VGND VGND VPWR VPWR _26630_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_453 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_464 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_475 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_486 _31994_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29348_ _29348_/A VGND VGND VPWR VPWR _34940_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_497 _32005_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17362_ _17149_/X _17358_/X _17361_/X _17152_/X VGND VGND VPWR VPWR _17362_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19101_ _19454_/A VGND VGND VPWR VPWR _19101_/X sky130_fd_sc_hd__buf_4
X_16313_ _33493_/Q _33429_/Q _33365_/Q _33301_/Q _15998_/X _15999_/X VGND VGND VPWR
+ VPWR _16313_/X sky130_fd_sc_hd__mux4_1
XFILLER_198_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29279_ _29279_/A VGND VGND VPWR VPWR _34907_/D sky130_fd_sc_hd__clkbuf_1
X_17293_ _34544_/Q _32432_/Q _34416_/Q _34352_/Q _17225_/X _17226_/X VGND VGND VPWR
+ VPWR _17293_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31310_ _35870_/Q input8/X _31316_/S VGND VGND VPWR VPWR _31311_/A sky130_fd_sc_hd__mux2_1
X_19032_ _19028_/X _19031_/X _18755_/X VGND VGND VPWR VPWR _19033_/D sky130_fd_sc_hd__o21ba_1
X_16244_ _34003_/Q _33939_/Q _33875_/Q _32147_/Q _16108_/X _16109_/X VGND VGND VPWR
+ VPWR _16244_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32290_ _35298_/CLK _32290_/D VGND VGND VPWR VPWR _32290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31241_ _31241_/A VGND VGND VPWR VPWR _35837_/D sky130_fd_sc_hd__clkbuf_1
X_16175_ _34257_/Q _34193_/Q _34129_/Q _34065_/Q _16005_/X _16007_/X VGND VGND VPWR
+ VPWR _16175_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput107 _31975_/Q VGND VGND VPWR VPWR D1[25] sky130_fd_sc_hd__buf_2
Xoutput118 _31985_/Q VGND VGND VPWR VPWR D1[35] sky130_fd_sc_hd__buf_2
XFILLER_182_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31172_ _31172_/A VGND VGND VPWR VPWR _35804_/D sky130_fd_sc_hd__clkbuf_1
Xoutput129 _31995_/Q VGND VGND VPWR VPWR D1[45] sky130_fd_sc_hd__buf_2
XFILLER_115_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30123_ _30192_/S VGND VGND VPWR VPWR _30142_/S sky130_fd_sc_hd__buf_4
X_19934_ _35834_/Q _32212_/Q _35706_/Q _35642_/Q _19613_/X _19614_/X VGND VGND VPWR
+ VPWR _19934_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35980_ _35981_/CLK _35980_/D VGND VGND VPWR VPWR _35980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_218_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30054_ _30054_/A VGND VGND VPWR VPWR _35275_/D sky130_fd_sc_hd__clkbuf_1
X_34931_ _34997_/CLK _34931_/D VGND VGND VPWR VPWR _34931_/Q sky130_fd_sc_hd__dfxtp_1
X_19865_ _33016_/Q _32952_/Q _32888_/Q _32824_/Q _19642_/X _19643_/X VGND VGND VPWR
+ VPWR _19865_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18816_ _34778_/Q _34714_/Q _34650_/Q _34586_/Q _18529_/X _18530_/X VGND VGND VPWR
+ VPWR _18816_/X sky130_fd_sc_hd__mux4_1
XTAP_6090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34862_ _35054_/CLK _34862_/D VGND VGND VPWR VPWR _34862_/Q sky130_fd_sc_hd__dfxtp_1
X_19796_ _19647_/X _19792_/X _19795_/X _19650_/X VGND VGND VPWR VPWR _19796_/X sky130_fd_sc_hd__a22o_1
X_33813_ _35730_/CLK _33813_/D VGND VGND VPWR VPWR _33813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18747_ _18743_/X _18744_/X _18745_/X _18746_/X VGND VGND VPWR VPWR _18747_/X sky130_fd_sc_hd__a22o_1
X_34793_ _34794_/CLK _34793_/D VGND VGND VPWR VPWR _34793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33744_ _34194_/CLK _33744_/D VGND VGND VPWR VPWR _33744_/Q sky130_fd_sc_hd__dfxtp_1
X_18678_ _18387_/X _18676_/X _18677_/X _18397_/X VGND VGND VPWR VPWR _18678_/X sky130_fd_sc_hd__a22o_1
X_30956_ _35702_/Q _29175_/X _30974_/S VGND VGND VPWR VPWR _30957_/A sky130_fd_sc_hd__mux2_1
XFILLER_224_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17629_ _17982_/A VGND VGND VPWR VPWR _17629_/X sky130_fd_sc_hd__buf_6
X_33675_ _35977_/CLK _33675_/D VGND VGND VPWR VPWR _33675_/Q sky130_fd_sc_hd__dfxtp_1
X_30887_ _30887_/A VGND VGND VPWR VPWR _35669_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_225_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35414_ _35927_/CLK _35414_/D VGND VGND VPWR VPWR _35414_/Q sky130_fd_sc_hd__dfxtp_1
X_20640_ _22442_/A VGND VGND VPWR VPWR _20640_/X sky130_fd_sc_hd__buf_2
X_32626_ _36141_/CLK _32626_/D VGND VGND VPWR VPWR _32626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20571_ _18356_/X _20569_/X _20570_/X _18368_/X VGND VGND VPWR VPWR _20571_/X sky130_fd_sc_hd__a22o_1
X_35345_ _35793_/CLK _35345_/D VGND VGND VPWR VPWR _35345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32557_ _35949_/CLK _32557_/D VGND VGND VPWR VPWR _32557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22310_ _22304_/X _22309_/X _22100_/X VGND VGND VPWR VPWR _22320_/C sky130_fd_sc_hd__o21ba_1
X_31508_ _23289_/X _35964_/Q _31514_/S VGND VGND VPWR VPWR _31509_/A sky130_fd_sc_hd__mux2_1
X_23290_ _32214_/Q _23289_/X _23301_/S VGND VGND VPWR VPWR _23291_/A sky130_fd_sc_hd__mux2_1
X_35276_ _35341_/CLK _35276_/D VGND VGND VPWR VPWR _35276_/Q sky130_fd_sc_hd__dfxtp_1
X_32488_ _34792_/CLK _32488_/D VGND VGND VPWR VPWR _32488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22241_ _22594_/A VGND VGND VPWR VPWR _22241_/X sky130_fd_sc_hd__buf_6
XFILLER_180_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31439_ _23127_/X _35931_/Q _31451_/S VGND VGND VPWR VPWR _31440_/A sky130_fd_sc_hd__mux2_1
X_34227_ _34227_/CLK _34227_/D VGND VGND VPWR VPWR _34227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22172_ _33208_/Q _32568_/Q _35960_/Q _35896_/Q _22027_/X _22028_/X VGND VGND VPWR
+ VPWR _22172_/X sky130_fd_sc_hd__mux4_1
X_34158_ _34222_/CLK _34158_/D VGND VGND VPWR VPWR _34158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21123_ _21048_/X _21121_/X _21122_/X _21053_/X VGND VGND VPWR VPWR _21123_/X sky130_fd_sc_hd__a22o_1
X_33109_ _36115_/CLK _33109_/D VGND VGND VPWR VPWR _33109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26980_ _26980_/A VGND VGND VPWR VPWR _33856_/D sky130_fd_sc_hd__clkbuf_1
X_34089_ _34153_/CLK _34089_/D VGND VGND VPWR VPWR _34089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25931_ _25931_/A VGND VGND VPWR VPWR _33384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21054_ _21048_/X _21049_/X _21052_/X _21053_/X VGND VGND VPWR VPWR _21054_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_1012 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1075 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20005_ _20160_/A VGND VGND VPWR VPWR _20005_/X sky130_fd_sc_hd__clkbuf_4
X_28650_ _28650_/A VGND VGND VPWR VPWR _34640_/D sky130_fd_sc_hd__clkbuf_1
X_25862_ _25171_/X _33352_/Q _25864_/S VGND VGND VPWR VPWR _25863_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27601_ _27601_/A VGND VGND VPWR VPWR _34143_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24813_ _23016_/X _32890_/Q _24823_/S VGND VGND VPWR VPWR _24814_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28581_ _26928_/X _34608_/Q _28591_/S VGND VGND VPWR VPWR _28582_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25793_ _25069_/X _33319_/Q _25801_/S VGND VGND VPWR VPWR _25794_/A sky130_fd_sc_hd__mux2_1
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27532_ _27559_/S VGND VGND VPWR VPWR _27551_/S sky130_fd_sc_hd__clkbuf_8
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24744_ _22914_/X _32857_/Q _24760_/S VGND VGND VPWR VPWR _24745_/A sky130_fd_sc_hd__mux2_1
X_21956_ _21952_/X _21953_/X _21954_/X _21955_/X VGND VGND VPWR VPWR _21956_/X sky130_fd_sc_hd__a22o_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20907_ _20903_/X _20906_/X _20700_/X VGND VGND VPWR VPWR _20908_/D sky130_fd_sc_hd__o21ba_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27463_ _26875_/X _34079_/Q _27467_/S VGND VGND VPWR VPWR _27464_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24675_ _24675_/A VGND VGND VPWR VPWR _32825_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21887_ _21883_/X _21886_/X _21747_/X VGND VGND VPWR VPWR _21897_/C sky130_fd_sc_hd__o21ba_1
X_29202_ _29202_/A VGND VGND VPWR VPWR _34878_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26414_ _28643_/B _26685_/B VGND VGND VPWR VPWR _26547_/S sky130_fd_sc_hd__nand2_8
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23626_ _23626_/A VGND VGND VPWR VPWR _32363_/D sky130_fd_sc_hd__clkbuf_1
X_20838_ _20838_/A _20838_/B _20838_/C _20838_/D VGND VGND VPWR VPWR _20839_/A sky130_fd_sc_hd__or4_2
X_27394_ _27394_/A VGND VGND VPWR VPWR _34046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29133_ _34856_/Q _29132_/X _29142_/S VGND VGND VPWR VPWR _29134_/A sky130_fd_sc_hd__mux2_1
X_26345_ _26345_/A VGND VGND VPWR VPWR _33580_/D sky130_fd_sc_hd__clkbuf_1
X_23557_ _23071_/X _32332_/Q _23559_/S VGND VGND VPWR VPWR _23558_/A sky130_fd_sc_hd__mux2_1
X_20769_ _35024_/Q _34960_/Q _34896_/Q _34832_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _20769_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22508_ _22508_/A VGND VGND VPWR VPWR _22508_/X sky130_fd_sc_hd__buf_6
X_29064_ input45/X VGND VGND VPWR VPWR _29064_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26276_ _26276_/A VGND VGND VPWR VPWR _33548_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23488_ _22969_/X _32299_/Q _23488_/S VGND VGND VPWR VPWR _23489_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28015_ _28015_/A VGND VGND VPWR VPWR _34339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25227_ _25227_/A VGND VGND VPWR VPWR _33055_/D sky130_fd_sc_hd__clkbuf_1
X_22439_ _32512_/Q _32384_/Q _32064_/Q _36032_/Q _22229_/X _22370_/X VGND VGND VPWR
+ VPWR _22439_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_1366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25158_ _25158_/A VGND VGND VPWR VPWR _33027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24109_ _24109_/A VGND VGND VPWR VPWR _24242_/S sky130_fd_sc_hd__buf_12
X_17980_ _33284_/Q _36164_/Q _33156_/Q _33092_/Q _17764_/X _17765_/X VGND VGND VPWR
+ VPWR _17980_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29966_ _29966_/A VGND VGND VPWR VPWR _35233_/D sky130_fd_sc_hd__clkbuf_1
X_25089_ _25088_/X _33005_/Q _25113_/S VGND VGND VPWR VPWR _25090_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16931_ _35558_/Q _35494_/Q _35430_/Q _35366_/Q _16897_/X _16898_/X VGND VGND VPWR
+ VPWR _16931_/X sky130_fd_sc_hd__mux4_1
X_28917_ _34767_/Q _24249_/X _28933_/S VGND VGND VPWR VPWR _28918_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29897_ _29897_/A VGND VGND VPWR VPWR _35200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16862_ _35812_/Q _32188_/Q _35684_/Q _35620_/Q _16607_/X _16608_/X VGND VGND VPWR
+ VPWR _16862_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19650_ _20158_/A VGND VGND VPWR VPWR _19650_/X sky130_fd_sc_hd__buf_4
X_28848_ _28848_/A VGND VGND VPWR VPWR _34734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_899 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18601_ _19307_/A VGND VGND VPWR VPWR _18601_/X sky130_fd_sc_hd__buf_4
XFILLER_111_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19581_ _35824_/Q _32201_/Q _35696_/Q _35632_/Q _19260_/X _19261_/X VGND VGND VPWR
+ VPWR _19581_/X sky130_fd_sc_hd__mux4_1
X_28779_ _28911_/S VGND VGND VPWR VPWR _28798_/S sky130_fd_sc_hd__clkbuf_8
X_16793_ _16646_/X _16791_/X _16792_/X _16649_/X VGND VGND VPWR VPWR _16793_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18532_ _35282_/Q _35218_/Q _35154_/Q _32274_/Q _18379_/X _18381_/X VGND VGND VPWR
+ VPWR _18532_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30810_ _23253_/X _35633_/Q _30818_/S VGND VGND VPWR VPWR _30811_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31790_ _31790_/A VGND VGND VPWR VPWR _36097_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30741_ _23093_/X _35600_/Q _30755_/S VGND VGND VPWR VPWR _30742_/A sky130_fd_sc_hd__mux2_1
X_18463_ _34768_/Q _34704_/Q _34640_/Q _34576_/Q _18375_/X _18376_/X VGND VGND VPWR
+ VPWR _18463_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_5_4_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_4_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_250 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_261 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_272 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _17906_/A VGND VGND VPWR VPWR _17414_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33460_ _33780_/CLK _33460_/D VGND VGND VPWR VPWR _33460_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_283 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18394_ _19457_/A VGND VGND VPWR VPWR _18394_/X sky130_fd_sc_hd__buf_4
X_30672_ _30672_/A VGND VGND VPWR VPWR _35567_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_294 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32411_ _34781_/CLK _32411_/D VGND VGND VPWR VPWR _32411_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _17063_/X _17341_/X _17344_/X _17067_/X VGND VGND VPWR VPWR _17345_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33391_ _33520_/CLK _33391_/D VGND VGND VPWR VPWR _33391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35130_ _35771_/CLK _35130_/D VGND VGND VPWR VPWR _35130_/Q sky130_fd_sc_hd__dfxtp_1
X_32342_ _36116_/CLK _32342_/D VGND VGND VPWR VPWR _32342_/Q sky130_fd_sc_hd__dfxtp_1
X_17276_ _17982_/A VGND VGND VPWR VPWR _17276_/X sky130_fd_sc_hd__buf_6
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19015_ _19010_/X _19012_/X _19013_/X _19014_/X VGND VGND VPWR VPWR _19015_/X sky130_fd_sc_hd__a22o_1
X_16227_ _16056_/X _16225_/X _16226_/X _16068_/X VGND VGND VPWR VPWR _16227_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35061_ _35061_/CLK _35061_/D VGND VGND VPWR VPWR _35061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32273_ _36216_/CLK _32273_/D VGND VGND VPWR VPWR _32273_/Q sky130_fd_sc_hd__dfxtp_1
X_34012_ _34074_/CLK _34012_/D VGND VGND VPWR VPWR _34012_/Q sky130_fd_sc_hd__dfxtp_1
X_31224_ _31224_/A VGND VGND VPWR VPWR _35829_/D sky130_fd_sc_hd__clkbuf_1
X_16158_ _16044_/X _16156_/X _16157_/X _16054_/X VGND VGND VPWR VPWR _16158_/X sky130_fd_sc_hd__a22o_1
XFILLER_138_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31155_ _31155_/A VGND VGND VPWR VPWR _35796_/D sky130_fd_sc_hd__clkbuf_1
X_16089_ _17762_/A VGND VGND VPWR VPWR _16873_/A sky130_fd_sc_hd__buf_12
XFILLER_114_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30106_ _30106_/A VGND VGND VPWR VPWR _35299_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19917_ _19917_/A VGND VGND VPWR VPWR _32121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35963_ _35963_/CLK _35963_/D VGND VGND VPWR VPWR _35963_/Q sky130_fd_sc_hd__dfxtp_1
X_31086_ _35764_/Q _29169_/X _31088_/S VGND VGND VPWR VPWR _31087_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30037_ _35267_/Q _29216_/X _30049_/S VGND VGND VPWR VPWR _30038_/A sky130_fd_sc_hd__mux2_1
X_34914_ _35299_/CLK _34914_/D VGND VGND VPWR VPWR _34914_/Q sky130_fd_sc_hd__dfxtp_1
X_19848_ _20201_/A VGND VGND VPWR VPWR _19848_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35894_ _36023_/CLK _35894_/D VGND VGND VPWR VPWR _35894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34845_ _34973_/CLK _34845_/D VGND VGND VPWR VPWR _34845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19779_ _34038_/Q _33974_/Q _33910_/Q _32246_/Q _19673_/X _19674_/X VGND VGND VPWR
+ VPWR _19779_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21810_ _21655_/X _21808_/X _21809_/X _21661_/X VGND VGND VPWR VPWR _21810_/X sky130_fd_sc_hd__a22o_1
X_22790_ _22508_/X _22788_/X _22789_/X _22511_/X VGND VGND VPWR VPWR _22790_/X sky130_fd_sc_hd__a22o_1
X_34776_ _35675_/CLK _34776_/D VGND VGND VPWR VPWR _34776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31988_ _36201_/CLK _31988_/D VGND VGND VPWR VPWR _31988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33727_ _33729_/CLK _33727_/D VGND VGND VPWR VPWR _33727_/Q sky130_fd_sc_hd__dfxtp_1
X_21741_ _22595_/A VGND VGND VPWR VPWR _21741_/X sky130_fd_sc_hd__buf_4
XFILLER_24_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30939_ _35694_/Q _29151_/X _30953_/S VGND VGND VPWR VPWR _30940_/A sky130_fd_sc_hd__mux2_1
XFILLER_225_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_969 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24460_ _22901_/X _32725_/Q _24464_/S VGND VGND VPWR VPWR _24461_/A sky130_fd_sc_hd__mux2_1
X_33658_ _34298_/CLK _33658_/D VGND VGND VPWR VPWR _33658_/Q sky130_fd_sc_hd__dfxtp_1
X_21672_ _21594_/X _21670_/X _21671_/X _21597_/X VGND VGND VPWR VPWR _21672_/X sky130_fd_sc_hd__a22o_1
X_23411_ _32264_/Q _23330_/X _23413_/S VGND VGND VPWR VPWR _23412_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20623_ _22506_/A VGND VGND VPWR VPWR _20623_/X sky130_fd_sc_hd__clkbuf_4
X_32609_ _36065_/CLK _32609_/D VGND VGND VPWR VPWR _32609_/Q sky130_fd_sc_hd__dfxtp_1
X_24391_ input42/X VGND VGND VPWR VPWR _24391_/X sky130_fd_sc_hd__clkbuf_4
X_33589_ _34292_/CLK _33589_/D VGND VGND VPWR VPWR _33589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26130_ _25168_/X _33479_/Q _26134_/S VGND VGND VPWR VPWR _26131_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35328_ _35328_/CLK _35328_/D VGND VGND VPWR VPWR _35328_/Q sky130_fd_sc_hd__dfxtp_1
X_23342_ input59/X VGND VGND VPWR VPWR _23342_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_193_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20554_ _19449_/A _20552_/X _20553_/X _19452_/A VGND VGND VPWR VPWR _20554_/X sky130_fd_sc_hd__a22o_1
XFILLER_36_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26061_ _25066_/X _33446_/Q _26071_/S VGND VGND VPWR VPWR _26062_/A sky130_fd_sc_hd__mux2_1
X_20485_ _33803_/Q _33739_/Q _33675_/Q _33611_/Q _20202_/X _20203_/X VGND VGND VPWR
+ VPWR _20485_/X sky130_fd_sc_hd__mux4_1
XFILLER_193_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35259_ _35515_/CLK _35259_/D VGND VGND VPWR VPWR _35259_/Q sky130_fd_sc_hd__dfxtp_1
X_23273_ _23273_/A VGND VGND VPWR VPWR _32208_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25012_ _25012_/A VGND VGND VPWR VPWR _32980_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22224_ _22220_/X _22223_/X _22081_/X VGND VGND VPWR VPWR _22250_/A sky130_fd_sc_hd__o21ba_1
XFILLER_161_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22155_ _22508_/A VGND VGND VPWR VPWR _22155_/X sky130_fd_sc_hd__clkbuf_4
X_29820_ _35164_/Q _29095_/X _29830_/S VGND VGND VPWR VPWR _29821_/A sky130_fd_sc_hd__mux2_1
XTAP_6804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21106_ _32986_/Q _32922_/Q _32858_/Q _32794_/Q _20883_/X _20884_/X VGND VGND VPWR
+ VPWR _21106_/X sky130_fd_sc_hd__mux4_1
XFILLER_248_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29751_ _29751_/A VGND VGND VPWR VPWR _35131_/D sky130_fd_sc_hd__clkbuf_1
X_26963_ _26962_/X _33851_/Q _26975_/S VGND VGND VPWR VPWR _26964_/A sky130_fd_sc_hd__mux2_1
X_22086_ _32502_/Q _32374_/Q _32054_/Q _36022_/Q _21876_/X _22017_/X VGND VGND VPWR
+ VPWR _22086_/X sky130_fd_sc_hd__mux4_1
XTAP_6859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28702_ _28702_/A VGND VGND VPWR VPWR _34665_/D sky130_fd_sc_hd__clkbuf_1
X_21037_ _20888_/X _21033_/X _21036_/X _20891_/X VGND VGND VPWR VPWR _21037_/X sky130_fd_sc_hd__a22o_1
X_25914_ _25914_/A VGND VGND VPWR VPWR _33376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29682_ _29682_/A VGND VGND VPWR VPWR _35098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26894_ input16/X VGND VGND VPWR VPWR _26894_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_248_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28633_ _27005_/X _34633_/Q _28633_/S VGND VGND VPWR VPWR _28634_/A sky130_fd_sc_hd__mux2_1
X_25845_ _25872_/S VGND VGND VPWR VPWR _25864_/S sky130_fd_sc_hd__buf_4
X_28564_ _26903_/X _34600_/Q _28570_/S VGND VGND VPWR VPWR _28565_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_842 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25776_ _25044_/X _33311_/Q _25780_/S VGND VGND VPWR VPWR _25777_/A sky130_fd_sc_hd__mux2_1
XFILLER_234_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22988_ input29/X VGND VGND VPWR VPWR _22988_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_167_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27515_ _27515_/A VGND VGND VPWR VPWR _34103_/D sky130_fd_sc_hd__clkbuf_1
X_24727_ _22889_/X _32849_/Q _24739_/S VGND VGND VPWR VPWR _24728_/A sky130_fd_sc_hd__mux2_1
X_28495_ _28495_/A VGND VGND VPWR VPWR _34567_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21939_ _33266_/Q _36146_/Q _33138_/Q _33074_/Q _21658_/X _21659_/X VGND VGND VPWR
+ VPWR _21939_/X sky130_fd_sc_hd__mux4_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27446_ _26850_/X _34071_/Q _27446_/S VGND VGND VPWR VPWR _27447_/A sky130_fd_sc_hd__mux2_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24658_ _24658_/A VGND VGND VPWR VPWR _32817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_203_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23609_ _32355_/Q _23152_/X _23625_/S VGND VGND VPWR VPWR _23610_/A sky130_fd_sc_hd__mux2_1
X_27377_ _34038_/Q _24369_/X _27395_/S VGND VGND VPWR VPWR _27378_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24589_ _24589_/A VGND VGND VPWR VPWR _32784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17130_ _32748_/Q _32684_/Q _32620_/Q _36076_/Q _16919_/X _17056_/X VGND VGND VPWR
+ VPWR _17130_/X sky130_fd_sc_hd__mux4_1
X_29116_ _29116_/A VGND VGND VPWR VPWR _34850_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26328_ _26328_/A VGND VGND VPWR VPWR _33572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29047_ _29047_/A VGND VGND VPWR VPWR _34829_/D sky130_fd_sc_hd__clkbuf_1
X_17061_ _17906_/A VGND VGND VPWR VPWR _17061_/X sky130_fd_sc_hd__buf_6
X_26259_ _25159_/X _33540_/Q _26269_/S VGND VGND VPWR VPWR _26260_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16012_ _15993_/X _16009_/X _16011_/X VGND VGND VPWR VPWR _16102_/A sky130_fd_sc_hd__o21ba_1
XFILLER_171_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17963_ _35331_/Q _35267_/Q _35203_/Q _32323_/Q _17712_/X _17713_/X VGND VGND VPWR
+ VPWR _17963_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29949_ _35225_/Q _29086_/X _29965_/S VGND VGND VPWR VPWR _29950_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19702_ _34292_/Q _34228_/Q _34164_/Q _34100_/Q _19389_/X _19390_/X VGND VGND VPWR
+ VPWR _19702_/X sky130_fd_sc_hd__mux4_1
XFILLER_214_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16914_ _16842_/X _16912_/X _16913_/X _16847_/X VGND VGND VPWR VPWR _16914_/X sky130_fd_sc_hd__a22o_1
X_32960_ _36098_/CLK _32960_/D VGND VGND VPWR VPWR _32960_/Q sky130_fd_sc_hd__dfxtp_1
X_17894_ _17855_/X _17892_/X _17893_/X _17858_/X VGND VGND VPWR VPWR _17894_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31911_ _23286_/X _36155_/Q _31919_/S VGND VGND VPWR VPWR _31912_/A sky130_fd_sc_hd__mux2_1
X_19633_ _19495_/X _19631_/X _19632_/X _19500_/X VGND VGND VPWR VPWR _19633_/X sky130_fd_sc_hd__a22o_1
XFILLER_238_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16845_ _33764_/Q _33700_/Q _33636_/Q _33572_/Q _16843_/X _16844_/X VGND VGND VPWR
+ VPWR _16845_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32891_ _36027_/CLK _32891_/D VGND VGND VPWR VPWR _32891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34630_ _34822_/CLK _34630_/D VGND VGND VPWR VPWR _34630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19564_ _19564_/A VGND VGND VPWR VPWR _32111_/D sky130_fd_sc_hd__buf_2
X_31842_ _23124_/X _36122_/Q _31856_/S VGND VGND VPWR VPWR _31843_/A sky130_fd_sc_hd__mux2_1
X_16776_ _16769_/X _16774_/X _16775_/X VGND VGND VPWR VPWR _16810_/A sky130_fd_sc_hd__o21ba_1
XFILLER_19_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18515_ _33234_/Q _36114_/Q _33106_/Q _33042_/Q _18320_/X _18321_/X VGND VGND VPWR
+ VPWR _18515_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34561_ _35777_/CLK _34561_/D VGND VGND VPWR VPWR _34561_/Q sky130_fd_sc_hd__dfxtp_1
X_31773_ _31773_/A VGND VGND VPWR VPWR _36089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19495_ _20201_/A VGND VGND VPWR VPWR _19495_/X sky130_fd_sc_hd__buf_2
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33512_ _33512_/CLK _33512_/D VGND VGND VPWR VPWR _33512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30724_ _30724_/A VGND VGND VPWR VPWR _35592_/D sky130_fd_sc_hd__clkbuf_1
X_18446_ _20165_/A VGND VGND VPWR VPWR _18446_/X sky130_fd_sc_hd__buf_4
XFILLER_59_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34492_ _35772_/CLK _34492_/D VGND VGND VPWR VPWR _34492_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36231_ _36232_/CLK _36231_/D VGND VGND VPWR VPWR _36231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18377_ _34766_/Q _34702_/Q _34638_/Q _34574_/Q _18375_/X _18376_/X VGND VGND VPWR
+ VPWR _18377_/X sky130_fd_sc_hd__mux4_1
X_33443_ _33507_/CLK _33443_/D VGND VGND VPWR VPWR _33443_/Q sky130_fd_sc_hd__dfxtp_1
X_30655_ _30655_/A VGND VGND VPWR VPWR _35559_/D sky130_fd_sc_hd__clkbuf_1
X_17328_ _17324_/X _17327_/X _17161_/X VGND VGND VPWR VPWR _17329_/D sky130_fd_sc_hd__o21ba_1
X_36162_ _36165_/CLK _36162_/D VGND VGND VPWR VPWR _36162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33374_ _33946_/CLK _33374_/D VGND VGND VPWR VPWR _33374_/Q sky130_fd_sc_hd__dfxtp_1
X_30586_ _23327_/X _35527_/Q _30590_/S VGND VGND VPWR VPWR _30587_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1006 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35113_ _35879_/CLK _35113_/D VGND VGND VPWR VPWR _35113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32325_ _35781_/CLK _32325_/D VGND VGND VPWR VPWR _32325_/Q sky130_fd_sc_hd__dfxtp_1
X_17259_ _34543_/Q _32431_/Q _34415_/Q _34351_/Q _17225_/X _17226_/X VGND VGND VPWR
+ VPWR _17259_/X sky130_fd_sc_hd__mux4_1
X_36093_ _36095_/CLK _36093_/D VGND VGND VPWR VPWR _36093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32256_ _33922_/CLK _32256_/D VGND VGND VPWR VPWR _32256_/Q sky130_fd_sc_hd__dfxtp_1
X_20270_ _20270_/A VGND VGND VPWR VPWR _32131_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_146_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35044_ _35300_/CLK _35044_/D VGND VGND VPWR VPWR _35044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31207_ _35821_/Q input25/X _31223_/S VGND VGND VPWR VPWR _31208_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_170_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _34317_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_157_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32187_ _35811_/CLK _32187_/D VGND VGND VPWR VPWR _32187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31138_ _35789_/Q _29246_/X _31138_/S VGND VGND VPWR VPWR _31139_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23960_ _23059_/X _32520_/Q _23962_/S VGND VGND VPWR VPWR _23961_/A sky130_fd_sc_hd__mux2_1
XTAP_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31069_ _31138_/S VGND VGND VPWR VPWR _31088_/S sky130_fd_sc_hd__buf_4
X_35946_ _35946_/CLK _35946_/D VGND VGND VPWR VPWR _35946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22911_ _23075_/S VGND VGND VPWR VPWR _22939_/S sky130_fd_sc_hd__buf_4
XFILLER_116_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35877_ _35941_/CLK _35877_/D VGND VGND VPWR VPWR _35877_/Q sky130_fd_sc_hd__dfxtp_1
X_23891_ _22957_/X _32487_/Q _23899_/S VGND VGND VPWR VPWR _23892_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25630_ _25630_/A VGND VGND VPWR VPWR _33242_/D sky130_fd_sc_hd__clkbuf_1
X_34828_ _35340_/CLK _34828_/D VGND VGND VPWR VPWR _34828_/Q sky130_fd_sc_hd__dfxtp_1
X_22842_ _22838_/X _22841_/X _22467_/A VGND VGND VPWR VPWR _22843_/D sky130_fd_sc_hd__o21ba_1
XFILLER_140_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25561_ _25561_/A VGND VGND VPWR VPWR _33211_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34759_ _34822_/CLK _34759_/D VGND VGND VPWR VPWR _34759_/Q sky130_fd_sc_hd__dfxtp_1
X_22773_ _33226_/Q _32586_/Q _35978_/Q _35914_/Q _20675_/X _20676_/X VGND VGND VPWR
+ VPWR _22773_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27300_ _27300_/A VGND VGND VPWR VPWR _34001_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24512_ _24512_/A VGND VGND VPWR VPWR _32749_/D sky130_fd_sc_hd__clkbuf_1
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28280_ _28280_/A VGND VGND VPWR VPWR _34465_/D sky130_fd_sc_hd__clkbuf_1
X_21724_ _22430_/A VGND VGND VPWR VPWR _21724_/X sky130_fd_sc_hd__buf_4
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25492_ _25492_/A VGND VGND VPWR VPWR _33178_/D sky130_fd_sc_hd__clkbuf_1
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27231_ _26931_/X _33969_/Q _27239_/S VGND VGND VPWR VPWR _27232_/A sky130_fd_sc_hd__mux2_1
X_24443_ input85/X input84/X input83/X _23561_/B VGND VGND VPWR VPWR _24444_/A sky130_fd_sc_hd__or4b_1
XFILLER_24_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21655_ _22501_/A VGND VGND VPWR VPWR _21655_/X sky130_fd_sc_hd__buf_6
XFILLER_123_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27162_ _26829_/X _33936_/Q _27176_/S VGND VGND VPWR VPWR _27163_/A sky130_fd_sc_hd__mux2_1
X_20606_ _20659_/A VGND VGND VPWR VPWR _22557_/A sky130_fd_sc_hd__buf_12
X_24374_ _32695_/Q _24373_/X _24398_/S VGND VGND VPWR VPWR _24375_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21586_ _33256_/Q _36136_/Q _33128_/Q _33064_/Q _21305_/X _21306_/X VGND VGND VPWR
+ VPWR _21586_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26113_ _25143_/X _33471_/Q _26113_/S VGND VGND VPWR VPWR _26114_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23325_ _32226_/Q _23228_/X _23350_/S VGND VGND VPWR VPWR _23326_/A sky130_fd_sc_hd__mux2_1
X_20537_ _35340_/Q _35276_/Q _35212_/Q _32332_/Q _18388_/X _18390_/X VGND VGND VPWR
+ VPWR _20537_/X sky130_fd_sc_hd__mux4_1
X_27093_ _27093_/A VGND VGND VPWR VPWR _33903_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26044_ _25041_/X _33438_/Q _26050_/S VGND VGND VPWR VPWR _26045_/A sky130_fd_sc_hd__mux2_1
X_20468_ _20464_/X _20467_/X _20142_/A _20143_/A VGND VGND VPWR VPWR _20483_/B sky130_fd_sc_hd__o211a_1
X_23256_ input30/X VGND VGND VPWR VPWR _23256_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_180_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22207_ _21952_/X _22205_/X _22206_/X _21955_/X VGND VGND VPWR VPWR _22207_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_161_CLK clkbuf_6_30__f_CLK/X VGND VGND VPWR VPWR _35977_/CLK sky130_fd_sc_hd__clkbuf_16
X_20399_ _34056_/Q _33992_/Q _33928_/Q _32264_/Q _18358_/X _18360_/X VGND VGND VPWR
+ VPWR _20399_/X sky130_fd_sc_hd__mux4_1
X_23187_ _32176_/Q _23121_/X _23206_/S VGND VGND VPWR VPWR _23188_/A sky130_fd_sc_hd__mux2_1
XTAP_6601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29803_ _35156_/Q _29070_/X _29809_/S VGND VGND VPWR VPWR _29804_/A sky130_fd_sc_hd__mux2_1
XTAP_6634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22138_ _22134_/X _22137_/X _22100_/X VGND VGND VPWR VPWR _22146_/C sky130_fd_sc_hd__o21ba_1
XTAP_5900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27995_ _26860_/X _34330_/Q _28009_/S VGND VGND VPWR VPWR _27996_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29734_ _29734_/A VGND VGND VPWR VPWR _35123_/D sky130_fd_sc_hd__clkbuf_1
X_26946_ input35/X VGND VGND VPWR VPWR _26946_/X sky130_fd_sc_hd__buf_4
XTAP_6689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22069_ _21754_/X _22067_/X _22068_/X _21759_/X VGND VGND VPWR VPWR _22069_/X sky130_fd_sc_hd__a22o_1
XTAP_5955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29665_ _29665_/A VGND VGND VPWR VPWR _35090_/D sky130_fd_sc_hd__clkbuf_1
X_26877_ _26877_/A VGND VGND VPWR VPWR _33823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16630_ _16496_/X _16628_/X _16629_/X _16499_/X VGND VGND VPWR VPWR _16630_/X sky130_fd_sc_hd__a22o_1
X_28616_ _28616_/A VGND VGND VPWR VPWR _34624_/D sky130_fd_sc_hd__clkbuf_1
X_25828_ _25828_/A VGND VGND VPWR VPWR _33335_/D sky130_fd_sc_hd__clkbuf_1
X_29596_ _35058_/Q _29163_/X _29602_/S VGND VGND VPWR VPWR _29597_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16561_ _16489_/X _16559_/X _16560_/X _16494_/X VGND VGND VPWR VPWR _16561_/X sky130_fd_sc_hd__a22o_1
X_25759_ _25019_/X _33303_/Q _25759_/S VGND VGND VPWR VPWR _25760_/A sky130_fd_sc_hd__mux2_1
X_28547_ _26878_/X _34592_/Q _28549_/S VGND VGND VPWR VPWR _28548_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18300_ _33486_/Q _33422_/Q _33358_/Q _33294_/Q _18298_/X _18299_/X VGND VGND VPWR
+ VPWR _18300_/X sky130_fd_sc_hd__mux4_1
X_19280_ _19142_/X _19278_/X _19279_/X _19147_/X VGND VGND VPWR VPWR _19280_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_6_55__f_CLK clkbuf_5_27_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_55__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_28478_ _28478_/A VGND VGND VPWR VPWR _34559_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16492_ _33754_/Q _33690_/Q _33626_/Q _33562_/Q _16490_/X _16491_/X VGND VGND VPWR
+ VPWR _16492_/X sky130_fd_sc_hd__mux4_1
X_18231_ _15977_/X _18229_/X _18230_/X _15987_/X VGND VGND VPWR VPWR _18231_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27429_ _27429_/A VGND VGND VPWR VPWR _34062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18162_ _32778_/Q _32714_/Q _32650_/Q _36106_/Q _17978_/X _16873_/A VGND VGND VPWR
+ VPWR _18162_/X sky130_fd_sc_hd__mux4_1
X_30440_ _30440_/A VGND VGND VPWR VPWR _35457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17113_ _16796_/X _17111_/X _17112_/X _16799_/X VGND VGND VPWR VPWR _17113_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18093_ _18093_/A _18093_/B _18093_/C _18093_/D VGND VGND VPWR VPWR _18094_/A sky130_fd_sc_hd__or4_4
XFILLER_117_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30371_ _23145_/X _35425_/Q _30371_/S VGND VGND VPWR VPWR _30372_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32110_ _35552_/CLK _32110_/D VGND VGND VPWR VPWR _32110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17044_ _16801_/X _17042_/X _17043_/X _16806_/X VGND VGND VPWR VPWR _17044_/X sky130_fd_sc_hd__a22o_1
X_33090_ _36165_/CLK _33090_/D VGND VGND VPWR VPWR _33090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32041_ _36009_/CLK _32041_/D VGND VGND VPWR VPWR _32041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_152_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _35339_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_171_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _33760_/Q _33696_/Q _33632_/Q _33568_/Q _18790_/X _18791_/X VGND VGND VPWR
+ VPWR _18995_/X sky130_fd_sc_hd__mux4_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35800_ _36063_/CLK _35800_/D VGND VGND VPWR VPWR _35800_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17946_ _32771_/Q _32707_/Q _32643_/Q _36099_/Q _17625_/X _17762_/X VGND VGND VPWR
+ VPWR _17946_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33992_ _34243_/CLK _33992_/D VGND VGND VPWR VPWR _33992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35731_ _35733_/CLK _35731_/D VGND VGND VPWR VPWR _35731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32943_ _33007_/CLK _32943_/D VGND VGND VPWR VPWR _32943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17877_ _17873_/X _17876_/X _17834_/X VGND VGND VPWR VPWR _17899_/A sky130_fd_sc_hd__o21ba_1
XFILLER_61_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19616_ _35761_/Q _35121_/Q _34481_/Q _33841_/Q _19440_/X _19441_/X VGND VGND VPWR
+ VPWR _19616_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35662_ _35727_/CLK _35662_/D VGND VGND VPWR VPWR _35662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16828_ _16641_/X _16826_/X _16827_/X _16644_/X VGND VGND VPWR VPWR _16828_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32874_ _36075_/CLK _32874_/D VGND VGND VPWR VPWR _32874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34613_ _35250_/CLK _34613_/D VGND VGND VPWR VPWR _34613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31825_ _23099_/X _36114_/Q _31835_/S VGND VGND VPWR VPWR _31826_/A sky130_fd_sc_hd__mux2_1
X_19547_ _35823_/Q _32200_/Q _35695_/Q _35631_/Q _19260_/X _19261_/X VGND VGND VPWR
+ VPWR _19547_/X sky130_fd_sc_hd__mux4_1
X_35593_ _35975_/CLK _35593_/D VGND VGND VPWR VPWR _35593_/Q sky130_fd_sc_hd__dfxtp_1
X_16759_ _35297_/Q _35233_/Q _35169_/Q _32289_/Q _16653_/X _16654_/X VGND VGND VPWR
+ VPWR _16759_/X sky130_fd_sc_hd__mux4_1
XFILLER_241_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34544_ _35954_/CLK _34544_/D VGND VGND VPWR VPWR _34544_/Q sky130_fd_sc_hd__dfxtp_1
X_31756_ _31756_/A VGND VGND VPWR VPWR _36081_/D sky130_fd_sc_hd__clkbuf_1
X_19478_ _19474_/X _19477_/X _19436_/X _19437_/X VGND VGND VPWR VPWR _19493_/B sky130_fd_sc_hd__o211a_1
XFILLER_146_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18429_ _18374_/X _18427_/X _18428_/X _18384_/X VGND VGND VPWR VPWR _18429_/X sky130_fd_sc_hd__a22o_1
X_30707_ _35584_/Q _29206_/X _30725_/S VGND VGND VPWR VPWR _30708_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1019 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34475_ _35944_/CLK _34475_/D VGND VGND VPWR VPWR _34475_/Q sky130_fd_sc_hd__dfxtp_1
X_31687_ _31687_/A VGND VGND VPWR VPWR _36048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_222_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36214_ _36216_/CLK _36214_/D VGND VGND VPWR VPWR _36214_/Q sky130_fd_sc_hd__dfxtp_1
X_33426_ _33490_/CLK _33426_/D VGND VGND VPWR VPWR _33426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21440_ _21440_/A _21440_/B _21440_/C _21440_/D VGND VGND VPWR VPWR _21441_/A sky130_fd_sc_hd__or4_4
X_30638_ _30638_/A VGND VGND VPWR VPWR _35551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21371_ _22430_/A VGND VGND VPWR VPWR _21371_/X sky130_fd_sc_hd__clkbuf_4
X_36145_ _36147_/CLK _36145_/D VGND VGND VPWR VPWR _36145_/Q sky130_fd_sc_hd__dfxtp_1
X_33357_ _34060_/CLK _33357_/D VGND VGND VPWR VPWR _33357_/Q sky130_fd_sc_hd__dfxtp_1
X_30569_ _23300_/X _35519_/Q _30569_/S VGND VGND VPWR VPWR _30570_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_391_CLK clkbuf_6_34__f_CLK/X VGND VGND VPWR VPWR _35757_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23110_ _23110_/A VGND VGND VPWR VPWR _32149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20322_ _35589_/Q _35525_/Q _35461_/Q _35397_/Q _20256_/X _20257_/X VGND VGND VPWR
+ VPWR _20322_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32308_ _35574_/CLK _32308_/D VGND VGND VPWR VPWR _32308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24090_ _23050_/X _32581_/Q _24098_/S VGND VGND VPWR VPWR _24091_/A sky130_fd_sc_hd__mux2_1
X_36076_ _36076_/CLK _36076_/D VGND VGND VPWR VPWR _36076_/Q sky130_fd_sc_hd__dfxtp_1
X_33288_ _36168_/CLK _33288_/D VGND VGND VPWR VPWR _33288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20253_ _35843_/Q _32222_/Q _35715_/Q _35651_/Q _19966_/X _19967_/X VGND VGND VPWR
+ VPWR _20253_/X sky130_fd_sc_hd__mux4_1
X_23041_ input48/X VGND VGND VPWR VPWR _23041_/X sky130_fd_sc_hd__clkbuf_4
X_35027_ _36204_/CLK _35027_/D VGND VGND VPWR VPWR _35027_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_143_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _35853_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_190_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32239_ _34032_/CLK _32239_/D VGND VGND VPWR VPWR _32239_/Q sky130_fd_sc_hd__dfxtp_1
X_20184_ _20180_/X _20183_/X _20142_/X _20143_/X VGND VGND VPWR VPWR _20199_/B sky130_fd_sc_hd__o211a_1
XFILLER_62_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26800_ _26800_/A VGND VGND VPWR VPWR _33795_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27780_ _27780_/A VGND VGND VPWR VPWR _34228_/D sky130_fd_sc_hd__clkbuf_1
X_24992_ _25187_/S VGND VGND VPWR VPWR _25020_/S sky130_fd_sc_hd__buf_4
XFILLER_130_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26731_ _26731_/A VGND VGND VPWR VPWR _33762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23943_ _23970_/S VGND VGND VPWR VPWR _23962_/S sky130_fd_sc_hd__buf_6
XTAP_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35929_ _35929_/CLK _35929_/D VGND VGND VPWR VPWR _35929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_218_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29450_ _29450_/A VGND VGND VPWR VPWR _34988_/D sky130_fd_sc_hd__clkbuf_1
X_26662_ _26662_/A VGND VGND VPWR VPWR _33730_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23874_ _22932_/X _32479_/Q _23878_/S VGND VGND VPWR VPWR _23875_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_805 _22895_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25613_ _25613_/A VGND VGND VPWR VPWR _33234_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_816 _22929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28401_ _28401_/A VGND VGND VPWR VPWR _34522_/D sky130_fd_sc_hd__clkbuf_1
X_29381_ _29381_/A VGND VGND VPWR VPWR _34956_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_226_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22825_ _32524_/Q _32396_/Q _32076_/Q _36044_/Q _22582_/X _21607_/A VGND VGND VPWR
+ VPWR _22825_/X sky130_fd_sc_hd__mux4_1
XANTENNA_827 _23121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26593_ _26683_/S VGND VGND VPWR VPWR _26612_/S sky130_fd_sc_hd__buf_4
XANTENNA_838 _23280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_849 _24244_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28332_ _34490_/Q _24382_/X _28342_/S VGND VGND VPWR VPWR _28333_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25544_ _25544_/A VGND VGND VPWR VPWR _33203_/D sky130_fd_sc_hd__clkbuf_1
X_22756_ _34314_/Q _34250_/Q _34186_/Q _34122_/Q _20645_/X _20646_/X VGND VGND VPWR
+ VPWR _22756_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21707_ _35563_/Q _35499_/Q _35435_/Q _35371_/Q _21497_/X _21498_/X VGND VGND VPWR
+ VPWR _21707_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28263_ _34457_/Q _24280_/X _28279_/S VGND VGND VPWR VPWR _28264_/A sky130_fd_sc_hd__mux2_1
X_25475_ _25475_/A VGND VGND VPWR VPWR _33170_/D sky130_fd_sc_hd__clkbuf_1
X_22687_ _35335_/Q _35271_/Q _35207_/Q _32327_/Q _20688_/X _20690_/X VGND VGND VPWR
+ VPWR _22687_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27214_ _26906_/X _33961_/Q _27218_/S VGND VGND VPWR VPWR _27215_/A sky130_fd_sc_hd__mux2_1
X_24426_ _32712_/Q _24425_/X _24429_/S VGND VGND VPWR VPWR _24427_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28194_ _28194_/A VGND VGND VPWR VPWR _34424_/D sky130_fd_sc_hd__clkbuf_1
X_21638_ _21634_/X _21637_/X _21394_/X VGND VGND VPWR VPWR _21646_/C sky130_fd_sc_hd__o21ba_1
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27145_ _27145_/A VGND VGND VPWR VPWR _33928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24357_ input30/X VGND VGND VPWR VPWR _24357_/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_382_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _35889_/CLK sky130_fd_sc_hd__clkbuf_16
X_21569_ _34791_/Q _34727_/Q _34663_/Q _34599_/Q _21535_/X _21536_/X VGND VGND VPWR
+ VPWR _21569_/X sky130_fd_sc_hd__mux4_1
XFILLER_193_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_924 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23308_ _32220_/Q _23307_/X _23334_/S VGND VGND VPWR VPWR _23309_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27076_ _27076_/A VGND VGND VPWR VPWR _33895_/D sky130_fd_sc_hd__clkbuf_1
X_24288_ _24288_/A VGND VGND VPWR VPWR _32667_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26027_ _25016_/X _33430_/Q _26029_/S VGND VGND VPWR VPWR _26028_/A sky130_fd_sc_hd__mux2_1
XTAP_7110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_134_CLK clkbuf_6_22__f_CLK/X VGND VGND VPWR VPWR _35664_/CLK sky130_fd_sc_hd__clkbuf_16
X_23239_ _32197_/Q _23237_/X _23268_/S VGND VGND VPWR VPWR _23240_/A sky130_fd_sc_hd__mux2_1
XTAP_7121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1204 _23127_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1215 _23559_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1226 _24394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1237 _25314_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17800_ _34047_/Q _33983_/Q _33919_/Q _32255_/Q _17726_/X _17727_/X VGND VGND VPWR
+ VPWR _17800_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1248 _26497_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15992_ _34254_/Q _34190_/Q _34126_/Q _34062_/Q _15989_/X _15991_/X VGND VGND VPWR
+ VPWR _15992_/X sky130_fd_sc_hd__mux4_1
X_18780_ _34777_/Q _34713_/Q _34649_/Q _34585_/Q _18529_/X _18530_/X VGND VGND VPWR
+ VPWR _18780_/X sky130_fd_sc_hd__mux4_1
XTAP_6475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27978_ _26835_/X _34322_/Q _27988_/S VGND VGND VPWR VPWR _27979_/A sky130_fd_sc_hd__mux2_1
XANTENNA_1259 _28371_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17731_ _32765_/Q _32701_/Q _32637_/Q _36093_/Q _17625_/X _17409_/X VGND VGND VPWR
+ VPWR _17731_/X sky130_fd_sc_hd__mux4_1
X_29717_ _29717_/A VGND VGND VPWR VPWR _35115_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26929_ _26928_/X _33840_/Q _26944_/S VGND VGND VPWR VPWR _26930_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29648_ _35083_/Q _29240_/X _29652_/S VGND VGND VPWR VPWR _29649_/A sky130_fd_sc_hd__mux2_1
X_17662_ _32507_/Q _32379_/Q _32059_/Q _36027_/Q _17629_/X _17417_/X VGND VGND VPWR
+ VPWR _17662_/X sky130_fd_sc_hd__mux4_1
XFILLER_224_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19401_ _33003_/Q _32939_/Q _32875_/Q _32811_/Q _19289_/X _19290_/X VGND VGND VPWR
+ VPWR _19401_/X sky130_fd_sc_hd__mux4_1
X_16613_ _33181_/Q _32541_/Q _35933_/Q _35869_/Q _16368_/X _16369_/X VGND VGND VPWR
+ VPWR _16613_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17593_ _32761_/Q _32697_/Q _32633_/Q _36089_/Q _17272_/X _17409_/X VGND VGND VPWR
+ VPWR _17593_/X sky130_fd_sc_hd__mux4_1
X_29579_ _35050_/Q _29138_/X _29581_/S VGND VGND VPWR VPWR _29580_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16544_ _17956_/A VGND VGND VPWR VPWR _16544_/X sky130_fd_sc_hd__buf_4
X_31610_ _36012_/Q input24/X _31628_/S VGND VGND VPWR VPWR _31611_/A sky130_fd_sc_hd__mux2_1
X_19332_ _35817_/Q _32194_/Q _35689_/Q _35625_/Q _19260_/X _19261_/X VGND VGND VPWR
+ VPWR _19332_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32590_ _36050_/CLK _32590_/D VGND VGND VPWR VPWR _32590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31541_ _23342_/X _35980_/Q _31543_/S VGND VGND VPWR VPWR _31542_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19263_ _35751_/Q _35111_/Q _34471_/Q _33831_/Q _19087_/X _19088_/X VGND VGND VPWR
+ VPWR _19263_/X sky130_fd_sc_hd__mux4_1
X_16475_ _16288_/X _16473_/X _16474_/X _16291_/X VGND VGND VPWR VPWR _16475_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18214_ _18214_/A VGND VGND VPWR VPWR _32011_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34260_ _34260_/CLK _34260_/D VGND VGND VPWR VPWR _34260_/Q sky130_fd_sc_hd__dfxtp_1
X_31472_ _23234_/X _35947_/Q _31472_/S VGND VGND VPWR VPWR _31473_/A sky130_fd_sc_hd__mux2_1
X_19194_ _35813_/Q _32189_/Q _35685_/Q _35621_/Q _18907_/X _18908_/X VGND VGND VPWR
+ VPWR _19194_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33211_ _36027_/CLK _33211_/D VGND VGND VPWR VPWR _33211_/Q sky130_fd_sc_hd__dfxtp_1
X_30423_ _30423_/A VGND VGND VPWR VPWR _35449_/D sky130_fd_sc_hd__clkbuf_1
X_18145_ _18141_/X _18144_/X _17853_/X VGND VGND VPWR VPWR _18153_/C sky130_fd_sc_hd__o21ba_1
XFILLER_191_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34191_ _34256_/CLK _34191_/D VGND VGND VPWR VPWR _34191_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_373_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _36015_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_184_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18076_ _33031_/Q _32967_/Q _32903_/Q _32839_/Q _15980_/X _15983_/X VGND VGND VPWR
+ VPWR _18076_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30354_ _30354_/A VGND VGND VPWR VPWR _35416_/D sky130_fd_sc_hd__clkbuf_1
X_33142_ _36087_/CLK _33142_/D VGND VGND VPWR VPWR _33142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17027_ _16702_/X _17025_/X _17026_/X _16708_/X VGND VGND VPWR VPWR _17027_/X sky130_fd_sc_hd__a22o_1
X_33073_ _33520_/CLK _33073_/D VGND VGND VPWR VPWR _33073_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_125_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _34004_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30285_ _30285_/A VGND VGND VPWR VPWR _35384_/D sky130_fd_sc_hd__clkbuf_1
X_32024_ _35995_/CLK _32024_/D VGND VGND VPWR VPWR _32024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18978_ _18974_/X _18977_/X _18730_/X _18731_/X VGND VGND VPWR VPWR _18993_/B sky130_fd_sc_hd__o211a_2
XFILLER_246_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _35330_/Q _35266_/Q _35202_/Q _32322_/Q _17712_/X _17713_/X VGND VGND VPWR
+ VPWR _17929_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33975_ _36152_/CLK _33975_/D VGND VGND VPWR VPWR _33975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35714_ _35715_/CLK _35714_/D VGND VGND VPWR VPWR _35714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20940_ _20940_/A _20940_/B _20940_/C _20940_/D VGND VGND VPWR VPWR _20941_/A sky130_fd_sc_hd__or4_1
XFILLER_54_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32926_ _35481_/CLK _32926_/D VGND VGND VPWR VPWR _32926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35645_ _35709_/CLK _35645_/D VGND VGND VPWR VPWR _35645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20871_ _20871_/A VGND VGND VPWR VPWR _36179_/D sky130_fd_sc_hd__clkbuf_1
X_32857_ _35995_/CLK _32857_/D VGND VGND VPWR VPWR _32857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22610_ _22508_/X _22608_/X _22609_/X _22511_/X VGND VGND VPWR VPWR _22610_/X sky130_fd_sc_hd__a22o_1
X_31808_ _31808_/A VGND VGND VPWR VPWR _36106_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35576_ _35638_/CLK _35576_/D VGND VGND VPWR VPWR _35576_/Q sky130_fd_sc_hd__dfxtp_1
X_23590_ _32346_/Q _23124_/X _23604_/S VGND VGND VPWR VPWR _23591_/A sky130_fd_sc_hd__mux2_1
X_32788_ _35002_/CLK _32788_/D VGND VGND VPWR VPWR _32788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22541_ _22501_/X _22539_/X _22540_/X _22506_/X VGND VGND VPWR VPWR _22541_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34527_ _35039_/CLK _34527_/D VGND VGND VPWR VPWR _34527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31739_ _31739_/A VGND VGND VPWR VPWR _36073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25260_ _25094_/X _33071_/Q _25272_/S VGND VGND VPWR VPWR _25261_/A sky130_fd_sc_hd__mux2_1
X_22472_ _34305_/Q _34241_/Q _34177_/Q _34113_/Q _22395_/X _22396_/X VGND VGND VPWR
+ VPWR _22472_/X sky130_fd_sc_hd__mux4_1
X_34458_ _35803_/CLK _34458_/D VGND VGND VPWR VPWR _34458_/Q sky130_fd_sc_hd__dfxtp_1
X_24211_ _23028_/X _32638_/Q _24213_/S VGND VGND VPWR VPWR _24212_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33409_ _34305_/CLK _33409_/D VGND VGND VPWR VPWR _33409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21423_ _32995_/Q _32931_/Q _32867_/Q _32803_/Q _21236_/X _21237_/X VGND VGND VPWR
+ VPWR _21423_/X sky130_fd_sc_hd__mux4_1
X_25191_ _24989_/X _33038_/Q _25209_/S VGND VGND VPWR VPWR _25192_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_364_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _34033_/CLK sky130_fd_sc_hd__clkbuf_16
X_34389_ _36196_/CLK _34389_/D VGND VGND VPWR VPWR _34389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24142_ _22926_/X _32605_/Q _24150_/S VGND VGND VPWR VPWR _24143_/A sky130_fd_sc_hd__mux2_1
X_36128_ _36128_/CLK _36128_/D VGND VGND VPWR VPWR _36128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_958 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21354_ _35553_/Q _35489_/Q _35425_/Q _35361_/Q _21144_/X _21145_/X VGND VGND VPWR
+ VPWR _21354_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20305_ _33797_/Q _33733_/Q _33669_/Q _33605_/Q _20202_/X _20203_/X VGND VGND VPWR
+ VPWR _20305_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_116_CLK clkbuf_6_20__f_CLK/X VGND VGND VPWR VPWR _36220_/CLK sky130_fd_sc_hd__clkbuf_16
X_24073_ _23025_/X _32573_/Q _24077_/S VGND VGND VPWR VPWR _24074_/A sky130_fd_sc_hd__mux2_1
X_36059_ _36059_/CLK _36059_/D VGND VGND VPWR VPWR _36059_/Q sky130_fd_sc_hd__dfxtp_1
X_28950_ _34783_/Q _24298_/X _28954_/S VGND VGND VPWR VPWR _28951_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21285_ _21281_/X _21284_/X _21041_/X VGND VGND VPWR VPWR _21293_/C sky130_fd_sc_hd__o21ba_1
XFILLER_89_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23024_ _23024_/A VGND VGND VPWR VPWR _32060_/D sky130_fd_sc_hd__clkbuf_1
X_27901_ _27901_/A VGND VGND VPWR VPWR _34285_/D sky130_fd_sc_hd__clkbuf_1
X_20236_ _20230_/X _20235_/X _20167_/X VGND VGND VPWR VPWR _20237_/D sky130_fd_sc_hd__o21ba_1
X_28881_ _28881_/A VGND VGND VPWR VPWR _34750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20167_ _20167_/A VGND VGND VPWR VPWR _20167_/X sky130_fd_sc_hd__clkbuf_4
X_27832_ _27832_/A VGND VGND VPWR VPWR _34253_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24975_ _23056_/X _32967_/Q _24979_/S VGND VGND VPWR VPWR _24976_/A sky130_fd_sc_hd__mux2_1
X_20098_ _19848_/X _20094_/X _20097_/X _19853_/X VGND VGND VPWR VPWR _20098_/X sky130_fd_sc_hd__a22o_1
XTAP_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27763_ _34220_/Q _24338_/X _27781_/S VGND VGND VPWR VPWR _27764_/A sky130_fd_sc_hd__mux2_1
XTAP_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29502_ _29502_/A VGND VGND VPWR VPWR _35013_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26714_ _26714_/A VGND VGND VPWR VPWR _33754_/D sky130_fd_sc_hd__clkbuf_1
X_23926_ _23926_/A VGND VGND VPWR VPWR _32503_/D sky130_fd_sc_hd__clkbuf_1
X_27694_ _34188_/Q _24437_/X _27696_/S VGND VGND VPWR VPWR _27695_/A sky130_fd_sc_hd__mux2_1
XTAP_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_602 _20167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26645_ _26645_/A VGND VGND VPWR VPWR _33722_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29433_ _29433_/A VGND VGND VPWR VPWR _34980_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_613 _18505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23857_ _22907_/X _32471_/Q _23857_/S VGND VGND VPWR VPWR _23858_/A sky130_fd_sc_hd__mux2_1
XTAP_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_624 _18680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_635 _19111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_646 _19463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22808_ _20644_/X _22806_/X _22807_/X _20654_/X VGND VGND VPWR VPWR _22808_/X sky130_fd_sc_hd__a22o_1
XANTENNA_657 _20363_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29364_ _23316_/X _34948_/Q _29374_/S VGND VGND VPWR VPWR _29365_/A sky130_fd_sc_hd__mux2_1
X_26576_ _26576_/A VGND VGND VPWR VPWR _33689_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_668 _22460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23788_ _23788_/A VGND VGND VPWR VPWR _32438_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_679 _22556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25527_ _25527_/A VGND VGND VPWR VPWR _33195_/D sky130_fd_sc_hd__clkbuf_1
X_28315_ _34482_/Q _24357_/X _28321_/S VGND VGND VPWR VPWR _28316_/A sky130_fd_sc_hd__mux2_1
X_22739_ _35849_/Q _32229_/Q _35721_/Q _35657_/Q _20589_/X _20591_/X VGND VGND VPWR
+ VPWR _22739_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29295_ _23152_/X _34915_/Q _29311_/S VGND VGND VPWR VPWR _29296_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28246_ _34449_/Q _24255_/X _28258_/S VGND VGND VPWR VPWR _28247_/A sky130_fd_sc_hd__mux2_1
X_16260_ _33171_/Q _32531_/Q _35923_/Q _35859_/Q _16063_/X _16065_/X VGND VGND VPWR
+ VPWR _16260_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25458_ _25186_/X _33165_/Q _25458_/S VGND VGND VPWR VPWR _25459_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24409_ _24409_/A VGND VGND VPWR VPWR _32706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16191_ _17846_/A VGND VGND VPWR VPWR _16191_/X sky130_fd_sc_hd__buf_6
X_28177_ _28177_/A VGND VGND VPWR VPWR _34416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_355_CLK clkbuf_6_44__f_CLK/X VGND VGND VPWR VPWR _35829_/CLK sky130_fd_sc_hd__clkbuf_16
X_25389_ _25458_/S VGND VGND VPWR VPWR _25408_/S sky130_fd_sc_hd__buf_6
XFILLER_139_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27128_ _26977_/X _33920_/Q _27146_/S VGND VGND VPWR VPWR _27129_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_107_CLK clkbuf_6_22__f_CLK/X VGND VGND VPWR VPWR _35727_/CLK sky130_fd_sc_hd__clkbuf_16
X_19950_ _19950_/A _19950_/B _19950_/C _19950_/D VGND VGND VPWR VPWR _19951_/A sky130_fd_sc_hd__or4_4
X_27059_ _27059_/A VGND VGND VPWR VPWR _33887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18901_ _33245_/Q _36125_/Q _33117_/Q _33053_/Q _18652_/X _18653_/X VGND VGND VPWR
+ VPWR _18901_/X sky130_fd_sc_hd__mux4_1
X_30070_ _30070_/A VGND VGND VPWR VPWR _35282_/D sky130_fd_sc_hd__clkbuf_1
X_19881_ _35064_/Q _35000_/Q _34936_/Q _34872_/Q _19809_/X _19810_/X VGND VGND VPWR
+ VPWR _19881_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1001 _17957_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1023 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1012 _17842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1023 _17865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18832_ _18796_/X _18830_/X _18831_/X _18799_/X VGND VGND VPWR VPWR _18832_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1034 _17853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1045 _17159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1056 _16309_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1067 _17090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18763_ _34009_/Q _33945_/Q _33881_/Q _32153_/Q _18614_/X _18615_/X VGND VGND VPWR
+ VPWR _18763_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1078 _17164_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15975_ input67/X input68/X VGND VGND VPWR VPWR _17761_/A sky130_fd_sc_hd__nor2b_4
XFILLER_110_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1089 _17232_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17714_ _35324_/Q _35260_/Q _35196_/Q _32316_/Q _17712_/X _17713_/X VGND VGND VPWR
+ VPWR _17714_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33760_ _34080_/CLK _33760_/D VGND VGND VPWR VPWR _33760_/Q sky130_fd_sc_hd__dfxtp_1
X_30972_ _35710_/Q _29200_/X _30974_/S VGND VGND VPWR VPWR _30973_/A sky130_fd_sc_hd__mux2_1
X_18694_ _32471_/Q _32343_/Q _32023_/Q _35991_/Q _18517_/X _18658_/X VGND VGND VPWR
+ VPWR _18694_/X sky130_fd_sc_hd__mux4_1
XTAP_4870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32711_ _36167_/CLK _32711_/D VGND VGND VPWR VPWR _32711_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17645_ _17502_/X _17643_/X _17644_/X _17505_/X VGND VGND VPWR VPWR _17645_/X sky130_fd_sc_hd__a22o_1
X_33691_ _34266_/CLK _33691_/D VGND VGND VPWR VPWR _33691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35430_ _35814_/CLK _35430_/D VGND VGND VPWR VPWR _35430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32642_ _33026_/CLK _32642_/D VGND VGND VPWR VPWR _32642_/Q sky130_fd_sc_hd__dfxtp_1
X_17576_ _35320_/Q _35256_/Q _35192_/Q _32312_/Q _17359_/X _17360_/X VGND VGND VPWR
+ VPWR _17576_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19315_ _19315_/A VGND VGND VPWR VPWR _32104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16527_ _33755_/Q _33691_/Q _33627_/Q _33563_/Q _16490_/X _16491_/X VGND VGND VPWR
+ VPWR _16527_/X sky130_fd_sc_hd__mux4_1
X_35361_ _35744_/CLK _35361_/D VGND VGND VPWR VPWR _35361_/Q sky130_fd_sc_hd__dfxtp_1
X_32573_ _35965_/CLK _32573_/D VGND VGND VPWR VPWR _32573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34312_ _34312_/CLK _34312_/D VGND VGND VPWR VPWR _34312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31524_ _31524_/A VGND VGND VPWR VPWR _35971_/D sky130_fd_sc_hd__clkbuf_1
X_19246_ _33767_/Q _33703_/Q _33639_/Q _33575_/Q _19143_/X _19144_/X VGND VGND VPWR
+ VPWR _19246_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16458_ _16458_/A VGND VGND VPWR VPWR _31960_/D sky130_fd_sc_hd__clkbuf_1
X_35292_ _35292_/CLK _35292_/D VGND VGND VPWR VPWR _35292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34243_ _34243_/CLK _34243_/D VGND VGND VPWR VPWR _34243_/Q sky130_fd_sc_hd__dfxtp_1
X_16389_ _16143_/X _16387_/X _16388_/X _16146_/X VGND VGND VPWR VPWR _16389_/X sky130_fd_sc_hd__a22o_1
X_31455_ _31455_/A VGND VGND VPWR VPWR _35938_/D sky130_fd_sc_hd__clkbuf_1
X_19177_ _19171_/X _19176_/X _19108_/X VGND VGND VPWR VPWR _19178_/D sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_346_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _33780_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18128_ _33545_/Q _33481_/Q _33417_/Q _33353_/Q _17829_/X _17830_/X VGND VGND VPWR
+ VPWR _18128_/X sky130_fd_sc_hd__mux4_1
X_30406_ _30406_/A VGND VGND VPWR VPWR _35441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31386_ _35906_/Q input48/X _31400_/S VGND VGND VPWR VPWR _31387_/A sky130_fd_sc_hd__mux2_1
X_34174_ _34302_/CLK _34174_/D VGND VGND VPWR VPWR _34174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33125_ _36132_/CLK _33125_/D VGND VGND VPWR VPWR _33125_/Q sky130_fd_sc_hd__dfxtp_1
X_18059_ _34566_/Q _32454_/Q _34438_/Q _34374_/Q _17931_/X _17932_/X VGND VGND VPWR
+ VPWR _18059_/X sky130_fd_sc_hd__mux4_1
X_30337_ _30337_/A VGND VGND VPWR VPWR _35408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21070_ _32985_/Q _32921_/Q _32857_/Q _32793_/Q _20883_/X _20884_/X VGND VGND VPWR
+ VPWR _21070_/X sky130_fd_sc_hd__mux4_1
X_30268_ _30268_/A VGND VGND VPWR VPWR _35376_/D sky130_fd_sc_hd__clkbuf_1
X_33056_ _34146_/CLK _33056_/D VGND VGND VPWR VPWR _33056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20021_ _20021_/A VGND VGND VPWR VPWR _32124_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32007_ _36194_/CLK _32007_/D VGND VGND VPWR VPWR _32007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30199_ _30199_/A VGND VGND VPWR VPWR _35343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24760_ _22938_/X _32865_/Q _24760_/S VGND VGND VPWR VPWR _24761_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21972_ _33523_/Q _33459_/Q _33395_/Q _33331_/Q _21723_/X _21724_/X VGND VGND VPWR
+ VPWR _21972_/X sky130_fd_sc_hd__mux4_1
X_33958_ _34087_/CLK _33958_/D VGND VGND VPWR VPWR _33958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23711_ _22892_/X _32402_/Q _23721_/S VGND VGND VPWR VPWR _23712_/A sky130_fd_sc_hd__mux2_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32909_ _34317_/CLK _32909_/D VGND VGND VPWR VPWR _32909_/Q sky130_fd_sc_hd__dfxtp_1
X_20923_ _32981_/Q _32917_/Q _32853_/Q _32789_/Q _20883_/X _20884_/X VGND VGND VPWR
+ VPWR _20923_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24691_ _23038_/X _32833_/Q _24707_/S VGND VGND VPWR VPWR _24692_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33889_ _34017_/CLK _33889_/D VGND VGND VPWR VPWR _33889_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26430_ _25013_/X _33621_/Q _26434_/S VGND VGND VPWR VPWR _26431_/A sky130_fd_sc_hd__mux2_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35628_ _35950_/CLK _35628_/D VGND VGND VPWR VPWR _35628_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23642_ _32371_/Q _23261_/X _23646_/S VGND VGND VPWR VPWR _23643_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20854_ _22395_/A VGND VGND VPWR VPWR _20854_/X sky130_fd_sc_hd__buf_6
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26361_ _26361_/A VGND VGND VPWR VPWR _33588_/D sky130_fd_sc_hd__clkbuf_1
X_23573_ _32338_/Q _23099_/X _23583_/S VGND VGND VPWR VPWR _23574_/A sky130_fd_sc_hd__mux2_1
X_35559_ _35879_/CLK _35559_/D VGND VGND VPWR VPWR _35559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20785_ _32977_/Q _32913_/Q _32849_/Q _32785_/Q _20633_/X _20635_/X VGND VGND VPWR
+ VPWR _20785_/X sky130_fd_sc_hd__mux4_1
X_28100_ _28100_/A VGND VGND VPWR VPWR _34380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25312_ _25171_/X _33096_/Q _25314_/S VGND VGND VPWR VPWR _25313_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22524_ _35586_/Q _35522_/Q _35458_/Q _35394_/Q _22203_/X _22204_/X VGND VGND VPWR
+ VPWR _22524_/X sky130_fd_sc_hd__mux4_1
X_29080_ _34839_/Q _29079_/X _29080_/S VGND VGND VPWR VPWR _29081_/A sky130_fd_sc_hd__mux2_1
X_26292_ _26292_/A VGND VGND VPWR VPWR _33555_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28031_ _28031_/A VGND VGND VPWR VPWR _34347_/D sky130_fd_sc_hd__clkbuf_1
X_25243_ _25069_/X _33063_/Q _25251_/S VGND VGND VPWR VPWR _25244_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22455_ _22455_/A VGND VGND VPWR VPWR _22455_/X sky130_fd_sc_hd__buf_4
XFILLER_210_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_337_CLK clkbuf_6_47__f_CLK/X VGND VGND VPWR VPWR _36150_/CLK sky130_fd_sc_hd__clkbuf_16
X_21406_ _21759_/A VGND VGND VPWR VPWR _21406_/X sky130_fd_sc_hd__clkbuf_4
X_25174_ input55/X VGND VGND VPWR VPWR _25174_/X sky130_fd_sc_hd__clkbuf_8
X_22386_ _35326_/Q _35262_/Q _35198_/Q _32318_/Q _22312_/X _22313_/X VGND VGND VPWR
+ VPWR _22386_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_861 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24125_ _22901_/X _32597_/Q _24129_/S VGND VGND VPWR VPWR _24126_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21337_ _22557_/A VGND VGND VPWR VPWR _21337_/X sky130_fd_sc_hd__buf_4
XFILLER_190_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29982_ _35241_/Q _29135_/X _29986_/S VGND VGND VPWR VPWR _29983_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28933_ _34775_/Q _24273_/X _28933_/S VGND VGND VPWR VPWR _28934_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24056_ _23000_/X _32565_/Q _24056_/S VGND VGND VPWR VPWR _24057_/A sky130_fd_sc_hd__mux2_1
X_21268_ _22447_/A VGND VGND VPWR VPWR _21268_/X sky130_fd_sc_hd__buf_4
XFILLER_132_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23007_ input36/X VGND VGND VPWR VPWR _23007_/X sky130_fd_sc_hd__clkbuf_4
X_20219_ _20069_/X _20217_/X _20218_/X _20073_/X VGND VGND VPWR VPWR _20219_/X sky130_fd_sc_hd__a22o_1
X_28864_ _26946_/X _34742_/Q _28882_/S VGND VGND VPWR VPWR _28865_/A sky130_fd_sc_hd__mux2_1
X_21199_ _21195_/X _21198_/X _21022_/X VGND VGND VPWR VPWR _21223_/A sky130_fd_sc_hd__o21ba_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27815_ _34245_/Q _24416_/X _27823_/S VGND VGND VPWR VPWR _27816_/A sky130_fd_sc_hd__mux2_1
XTAP_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28795_ _28795_/A VGND VGND VPWR VPWR _34709_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24958_ _23031_/X _32959_/Q _24958_/S VGND VGND VPWR VPWR _24959_/A sky130_fd_sc_hd__mux2_1
XTAP_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27746_ _34212_/Q _24314_/X _27760_/S VGND VGND VPWR VPWR _27747_/A sky130_fd_sc_hd__mux2_1
XTAP_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23909_ _23909_/A VGND VGND VPWR VPWR _32495_/D sky130_fd_sc_hd__clkbuf_1
X_27677_ _27677_/A VGND VGND VPWR VPWR _34179_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24889_ _22929_/X _32926_/Q _24895_/S VGND VGND VPWR VPWR _24890_/A sky130_fd_sc_hd__mux2_1
XANTENNA_410 _36212_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_421 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29416_ _29416_/A VGND VGND VPWR VPWR _34972_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_432 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17430_ _17352_/X _17426_/X _17429_/X _17355_/X VGND VGND VPWR VPWR _17430_/X sky130_fd_sc_hd__a22o_1
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26628_ _26628_/A VGND VGND VPWR VPWR _33714_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_443 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_454 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_465 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_1160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_476 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29347_ _23289_/X _34940_/Q _29353_/S VGND VGND VPWR VPWR _29348_/A sky130_fd_sc_hd__mux2_1
X_17361_ _35314_/Q _35250_/Q _35186_/Q _32306_/Q _17359_/X _17360_/X VGND VGND VPWR
+ VPWR _17361_/X sky130_fd_sc_hd__mux4_1
XANTENNA_487 _31994_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26559_ _26559_/A VGND VGND VPWR VPWR _33681_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_498 _32008_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19100_ _19096_/X _19097_/X _19098_/X _19099_/X VGND VGND VPWR VPWR _19100_/X sky130_fd_sc_hd__a22o_1
X_16312_ _16136_/X _16310_/X _16311_/X _16141_/X VGND VGND VPWR VPWR _16312_/X sky130_fd_sc_hd__a22o_1
XFILLER_144_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17292_ _17149_/X _17290_/X _17291_/X _17152_/X VGND VGND VPWR VPWR _17292_/X sky130_fd_sc_hd__a22o_1
XFILLER_13_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29278_ _23127_/X _34907_/Q _29290_/S VGND VGND VPWR VPWR _29279_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16243_ _33491_/Q _33427_/Q _33363_/Q _33299_/Q _15998_/X _15999_/X VGND VGND VPWR
+ VPWR _16243_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19031_ _18748_/X _19029_/X _19030_/X _18753_/X VGND VGND VPWR VPWR _19031_/X sky130_fd_sc_hd__a22o_1
X_28229_ _28229_/A VGND VGND VPWR VPWR _34441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_328_CLK clkbuf_6_44__f_CLK/X VGND VGND VPWR VPWR _36085_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31240_ _35837_/Q input42/X _31244_/S VGND VGND VPWR VPWR _31241_/A sky130_fd_sc_hd__mux2_1
X_16174_ _33745_/Q _33681_/Q _33617_/Q _33553_/Q _16137_/X _16138_/X VGND VGND VPWR
+ VPWR _16174_/X sky130_fd_sc_hd__mux4_1
XFILLER_126_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput108 _31976_/Q VGND VGND VPWR VPWR D1[26] sky130_fd_sc_hd__buf_2
X_31171_ _35804_/Q input6/X _31181_/S VGND VGND VPWR VPWR _31172_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput119 _31986_/Q VGND VGND VPWR VPWR D1[36] sky130_fd_sc_hd__buf_2
XFILLER_141_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30122_ _30122_/A VGND VGND VPWR VPWR _35307_/D sky130_fd_sc_hd__clkbuf_1
X_19933_ _19928_/X _19932_/X _19789_/X _19790_/X VGND VGND VPWR VPWR _19950_/B sky130_fd_sc_hd__o211a_1
XFILLER_218_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30053_ _35275_/Q _29240_/X _30057_/S VGND VGND VPWR VPWR _30054_/A sky130_fd_sc_hd__mux2_1
X_34930_ _35826_/CLK _34930_/D VGND VGND VPWR VPWR _34930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19864_ _32504_/Q _32376_/Q _32056_/Q _36024_/Q _19576_/X _19717_/X VGND VGND VPWR
+ VPWR _19864_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_2__f_CLK clkbuf_5_1_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_2__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_229_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput90 _31950_/Q VGND VGND VPWR VPWR D1[0] sky130_fd_sc_hd__buf_2
XFILLER_95_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18815_ _18811_/X _18814_/X _18741_/X VGND VGND VPWR VPWR _18825_/C sky130_fd_sc_hd__o21ba_1
XTAP_6080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34861_ _35757_/CLK _34861_/D VGND VGND VPWR VPWR _34861_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19795_ _35766_/Q _35126_/Q _34486_/Q _33846_/Q _19793_/X _19794_/X VGND VGND VPWR
+ VPWR _19795_/X sky130_fd_sc_hd__mux4_1
XFILLER_231_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33812_ _35667_/CLK _33812_/D VGND VGND VPWR VPWR _33812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18746_ _19452_/A VGND VGND VPWR VPWR _18746_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34792_ _34792_/CLK _34792_/D VGND VGND VPWR VPWR _34792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33743_ _34256_/CLK _33743_/D VGND VGND VPWR VPWR _33743_/Q sky130_fd_sc_hd__dfxtp_1
X_18677_ _35030_/Q _34966_/Q _34902_/Q _34838_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _18677_/X sky130_fd_sc_hd__mux4_1
X_30955_ _31003_/S VGND VGND VPWR VPWR _30974_/S sky130_fd_sc_hd__buf_4
XFILLER_102_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17628_ _17408_/X _17626_/X _17627_/X _17414_/X VGND VGND VPWR VPWR _17628_/X sky130_fd_sc_hd__a22o_1
X_33674_ _34251_/CLK _33674_/D VGND VGND VPWR VPWR _33674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30886_ _35669_/Q _29073_/X _30890_/S VGND VGND VPWR VPWR _30887_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35413_ _35925_/CLK _35413_/D VGND VGND VPWR VPWR _35413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32625_ _33262_/CLK _32625_/D VGND VGND VPWR VPWR _32625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17559_ _17555_/X _17556_/X _17557_/X _17558_/X VGND VGND VPWR VPWR _17559_/X sky130_fd_sc_hd__a22o_1
X_35344_ _35793_/CLK _35344_/D VGND VGND VPWR VPWR _35344_/Q sky130_fd_sc_hd__dfxtp_1
X_20570_ _35085_/Q _35021_/Q _34957_/Q _34893_/Q _18379_/X _18381_/X VGND VGND VPWR
+ VPWR _20570_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32556_ _35949_/CLK _32556_/D VGND VGND VPWR VPWR _32556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31507_ _31507_/A VGND VGND VPWR VPWR _35963_/D sky130_fd_sc_hd__clkbuf_1
X_19229_ _35750_/Q _35110_/Q _34470_/Q _33830_/Q _19087_/X _19088_/X VGND VGND VPWR
+ VPWR _19229_/X sky130_fd_sc_hd__mux4_1
X_35275_ _35338_/CLK _35275_/D VGND VGND VPWR VPWR _35275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_319_CLK clkbuf_6_39__f_CLK/X VGND VGND VPWR VPWR _35638_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_191_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32487_ _34792_/CLK _32487_/D VGND VGND VPWR VPWR _32487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22240_ _22236_/X _22239_/X _22100_/X VGND VGND VPWR VPWR _22250_/C sky130_fd_sc_hd__o21ba_1
XFILLER_9_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34226_ _34291_/CLK _34226_/D VGND VGND VPWR VPWR _34226_/Q sky130_fd_sc_hd__dfxtp_1
X_31438_ _31438_/A VGND VGND VPWR VPWR _35930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34157_ _35252_/CLK _34157_/D VGND VGND VPWR VPWR _34157_/Q sky130_fd_sc_hd__dfxtp_1
X_22171_ _35576_/Q _35512_/Q _35448_/Q _35384_/Q _21850_/X _21851_/X VGND VGND VPWR
+ VPWR _22171_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31369_ _35898_/Q input39/X _31379_/S VGND VGND VPWR VPWR _31370_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33108_ _36117_/CLK _33108_/D VGND VGND VPWR VPWR _33108_/Q sky130_fd_sc_hd__dfxtp_1
X_21122_ _35034_/Q _34970_/Q _34906_/Q _34842_/Q _21050_/X _21051_/X VGND VGND VPWR
+ VPWR _21122_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34088_ _34153_/CLK _34088_/D VGND VGND VPWR VPWR _34088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33039_ _36112_/CLK _33039_/D VGND VGND VPWR VPWR _33039_/Q sky130_fd_sc_hd__dfxtp_1
X_25930_ _25072_/X _33384_/Q _25936_/S VGND VGND VPWR VPWR _25931_/A sky130_fd_sc_hd__mux2_1
X_21053_ _21759_/A VGND VGND VPWR VPWR _21053_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_119_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1062 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20004_ _20000_/X _20001_/X _20002_/X _20003_/X VGND VGND VPWR VPWR _20004_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25861_ _25861_/A VGND VGND VPWR VPWR _33351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24812_ _24812_/A VGND VGND VPWR VPWR _32889_/D sky130_fd_sc_hd__clkbuf_1
X_27600_ _34143_/Q _24298_/X _27604_/S VGND VGND VPWR VPWR _27601_/A sky130_fd_sc_hd__mux2_1
X_25792_ _25792_/A VGND VGND VPWR VPWR _33318_/D sky130_fd_sc_hd__clkbuf_1
X_28580_ _28580_/A VGND VGND VPWR VPWR _34607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27531_ _27531_/A VGND VGND VPWR VPWR _34111_/D sky130_fd_sc_hd__clkbuf_1
X_24743_ _24743_/A VGND VGND VPWR VPWR _32856_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21955_ _22465_/A VGND VGND VPWR VPWR _21955_/X sky130_fd_sc_hd__buf_4
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20906_ _20687_/X _20904_/X _20905_/X _20697_/X VGND VGND VPWR VPWR _20906_/X sky130_fd_sc_hd__a22o_1
XFILLER_27_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27462_ _27462_/A VGND VGND VPWR VPWR _34078_/D sky130_fd_sc_hd__clkbuf_1
X_24674_ _23013_/X _32825_/Q _24686_/S VGND VGND VPWR VPWR _24675_/A sky130_fd_sc_hd__mux2_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21886_ _21599_/X _21884_/X _21885_/X _21602_/X VGND VGND VPWR VPWR _21886_/X sky130_fd_sc_hd__a22o_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29201_ _34878_/Q _29200_/X _29204_/S VGND VGND VPWR VPWR _29202_/A sky130_fd_sc_hd__mux2_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26413_ _26413_/A VGND VGND VPWR VPWR _33613_/D sky130_fd_sc_hd__clkbuf_1
X_23625_ _32363_/Q _23234_/X _23625_/S VGND VGND VPWR VPWR _23626_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20837_ _20833_/X _20836_/X _20700_/X VGND VGND VPWR VPWR _20838_/D sky130_fd_sc_hd__o21ba_1
X_27393_ _34046_/Q _24394_/X _27395_/S VGND VGND VPWR VPWR _27394_/A sky130_fd_sc_hd__mux2_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29132_ input19/X VGND VGND VPWR VPWR _29132_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_35_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26344_ _25084_/X _33580_/Q _26362_/S VGND VGND VPWR VPWR _26345_/A sky130_fd_sc_hd__mux2_1
X_23556_ _23556_/A VGND VGND VPWR VPWR _32331_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20768_ _34512_/Q _32400_/Q _34384_/Q _34320_/Q _20766_/X _20767_/X VGND VGND VPWR
+ VPWR _20768_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22507_ _22501_/X _22504_/X _22505_/X _22506_/X VGND VGND VPWR VPWR _22507_/X sky130_fd_sc_hd__a22o_1
X_29063_ _29063_/A VGND VGND VPWR VPWR _34833_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26275_ _25183_/X _33548_/Q _26277_/S VGND VGND VPWR VPWR _26276_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23487_ _23487_/A VGND VGND VPWR VPWR _32298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20699_ input76/X input75/X VGND VGND VPWR VPWR _22467_/A sky130_fd_sc_hd__or2b_4
XFILLER_182_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28014_ _26888_/X _34339_/Q _28030_/S VGND VGND VPWR VPWR _28015_/A sky130_fd_sc_hd__mux2_1
X_25226_ _25044_/X _33055_/Q _25230_/S VGND VGND VPWR VPWR _25227_/A sky130_fd_sc_hd__mux2_1
X_22438_ _22361_/X _22436_/X _22437_/X _22367_/X VGND VGND VPWR VPWR _22438_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25157_ _25156_/X _33027_/Q _25175_/S VGND VGND VPWR VPWR _25158_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22369_ _22369_/A VGND VGND VPWR VPWR _22369_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_237_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24108_ _31680_/A input83/X _23561_/B VGND VGND VPWR VPWR _24109_/A sky130_fd_sc_hd__or3b_1
XFILLER_237_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29965_ _35233_/Q _29110_/X _29965_/S VGND VGND VPWR VPWR _29966_/A sky130_fd_sc_hd__mux2_1
X_25088_ input25/X VGND VGND VPWR VPWR _25088_/X sky130_fd_sc_hd__buf_6
XFILLER_123_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28916_ _28916_/A VGND VGND VPWR VPWR _34766_/D sky130_fd_sc_hd__clkbuf_1
X_16930_ _16641_/X _16928_/X _16929_/X _16644_/X VGND VGND VPWR VPWR _16930_/X sky130_fd_sc_hd__a22o_1
X_24039_ _24039_/A VGND VGND VPWR VPWR _32556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29896_ _35200_/Q _29206_/X _29914_/S VGND VGND VPWR VPWR _29897_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28847_ _26922_/X _34734_/Q _28861_/S VGND VGND VPWR VPWR _28848_/A sky130_fd_sc_hd__mux2_1
X_16861_ _16857_/X _16860_/X _16783_/X _16784_/X VGND VGND VPWR VPWR _16878_/B sky130_fd_sc_hd__o211a_1
XFILLER_77_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18600_ _20012_/A VGND VGND VPWR VPWR _18600_/X sky130_fd_sc_hd__buf_6
XFILLER_120_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19580_ _19575_/X _19579_/X _19436_/X _19437_/X VGND VGND VPWR VPWR _19597_/B sky130_fd_sc_hd__o211a_1
XFILLER_237_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28778_ _31815_/A _28778_/B VGND VGND VPWR VPWR _28911_/S sky130_fd_sc_hd__nand2_8
X_16792_ _33186_/Q _32546_/Q _35938_/Q _35874_/Q _16721_/X _16722_/X VGND VGND VPWR
+ VPWR _16792_/X sky130_fd_sc_hd__mux4_1
XFILLER_237_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_1211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18531_ _34770_/Q _34706_/Q _34642_/Q _34578_/Q _18529_/X _18530_/X VGND VGND VPWR
+ VPWR _18531_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27729_ _34204_/Q _24289_/X _27739_/S VGND VGND VPWR VPWR _27730_/A sky130_fd_sc_hd__mux2_1
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30740_ _30740_/A VGND VGND VPWR VPWR _35599_/D sky130_fd_sc_hd__clkbuf_1
X_18462_ _18458_/X _18461_/X _18371_/X VGND VGND VPWR VPWR _18472_/C sky130_fd_sc_hd__o21ba_1
XFILLER_18_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_240 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_251 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_262 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _33268_/Q _36148_/Q _33140_/Q _33076_/Q _17411_/X _17412_/X VGND VGND VPWR
+ VPWR _17413_/X sky130_fd_sc_hd__mux4_1
XANTENNA_273 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_284 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30671_ _35567_/Q _29154_/X _30683_/S VGND VGND VPWR VPWR _30672_/A sky130_fd_sc_hd__mux2_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18393_ _20070_/A VGND VGND VPWR VPWR _19457_/A sky130_fd_sc_hd__buf_12
XFILLER_92_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_295 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32410_ _34781_/CLK _32410_/D VGND VGND VPWR VPWR _32410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _33010_/Q _32946_/Q _32882_/Q _32818_/Q _17342_/X _17343_/X VGND VGND VPWR
+ VPWR _17344_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33390_ _36147_/CLK _33390_/D VGND VGND VPWR VPWR _33390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32341_ _36052_/CLK _32341_/D VGND VGND VPWR VPWR _32341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17275_ _17055_/X _17273_/X _17274_/X _17061_/X VGND VGND VPWR VPWR _17275_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19014_ _20211_/A VGND VGND VPWR VPWR _19014_/X sky130_fd_sc_hd__clkbuf_4
X_16226_ _33170_/Q _32530_/Q _35922_/Q _35858_/Q _16063_/X _16065_/X VGND VGND VPWR
+ VPWR _16226_/X sky130_fd_sc_hd__mux4_1
X_35060_ _35061_/CLK _35060_/D VGND VGND VPWR VPWR _35060_/Q sky130_fd_sc_hd__dfxtp_1
X_32272_ _35281_/CLK _32272_/D VGND VGND VPWR VPWR _32272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34011_ _34267_/CLK _34011_/D VGND VGND VPWR VPWR _34011_/Q sky130_fd_sc_hd__dfxtp_1
X_16157_ _35728_/Q _35088_/Q _34448_/Q _33808_/Q _16049_/X _16051_/X VGND VGND VPWR
+ VPWR _16157_/X sky130_fd_sc_hd__mux4_1
X_31223_ _35829_/Q input33/X _31223_/S VGND VGND VPWR VPWR _31224_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16088_ _17712_/A VGND VGND VPWR VPWR _16088_/X sky130_fd_sc_hd__buf_6
X_31154_ _35796_/Q input61/X _31160_/S VGND VGND VPWR VPWR _31155_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19916_ _19916_/A _19916_/B _19916_/C _19916_/D VGND VGND VPWR VPWR _19917_/A sky130_fd_sc_hd__or4_4
X_30105_ _35299_/Q _29117_/X _30121_/S VGND VGND VPWR VPWR _30106_/A sky130_fd_sc_hd__mux2_1
X_35962_ _35963_/CLK _35962_/D VGND VGND VPWR VPWR _35962_/Q sky130_fd_sc_hd__dfxtp_1
X_31085_ _31085_/A VGND VGND VPWR VPWR _35763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30036_ _30036_/A VGND VGND VPWR VPWR _35266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34913_ _35040_/CLK _34913_/D VGND VGND VPWR VPWR _34913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19847_ _19847_/A VGND VGND VPWR VPWR _32119_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35893_ _35958_/CLK _35893_/D VGND VGND VPWR VPWR _35893_/Q sky130_fd_sc_hd__dfxtp_1
X_34844_ _35036_/CLK _34844_/D VGND VGND VPWR VPWR _34844_/Q sky130_fd_sc_hd__dfxtp_1
X_19778_ _33526_/Q _33462_/Q _33398_/Q _33334_/Q _19776_/X _19777_/X VGND VGND VPWR
+ VPWR _19778_/X sky130_fd_sc_hd__mux4_1
XFILLER_216_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18729_ _18657_/X _18727_/X _18728_/X _18661_/X VGND VGND VPWR VPWR _18729_/X sky130_fd_sc_hd__a22o_1
X_34775_ _34775_/CLK _34775_/D VGND VGND VPWR VPWR _34775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1000 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31987_ _36201_/CLK _31987_/D VGND VGND VPWR VPWR _31987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33726_ _33729_/CLK _33726_/D VGND VGND VPWR VPWR _33726_/Q sky130_fd_sc_hd__dfxtp_1
X_21740_ _22594_/A VGND VGND VPWR VPWR _21740_/X sky130_fd_sc_hd__buf_6
XFILLER_184_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30938_ _30938_/A VGND VGND VPWR VPWR _35693_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33657_ _34296_/CLK _33657_/D VGND VGND VPWR VPWR _33657_/Q sky130_fd_sc_hd__dfxtp_1
X_21671_ _35754_/Q _35114_/Q _34474_/Q _33834_/Q _21387_/X _21388_/X VGND VGND VPWR
+ VPWR _21671_/X sky130_fd_sc_hd__mux4_1
X_30869_ _30869_/A VGND VGND VPWR VPWR _35661_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_96_CLK clkbuf_leaf_96_CLK/A VGND VGND VPWR VPWR _34706_/CLK sky130_fd_sc_hd__clkbuf_16
X_23410_ _23410_/A VGND VGND VPWR VPWR _32263_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20622_ _33230_/Q _36110_/Q _33102_/Q _33038_/Q _20620_/X _20621_/X VGND VGND VPWR
+ VPWR _20622_/X sky130_fd_sc_hd__mux4_1
X_32608_ _36128_/CLK _32608_/D VGND VGND VPWR VPWR _32608_/Q sky130_fd_sc_hd__dfxtp_1
X_24390_ _24390_/A VGND VGND VPWR VPWR _32700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33588_ _34292_/CLK _33588_/D VGND VGND VPWR VPWR _33588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23341_ _23341_/A VGND VGND VPWR VPWR _32231_/D sky130_fd_sc_hd__clkbuf_1
X_35327_ _35581_/CLK _35327_/D VGND VGND VPWR VPWR _35327_/Q sky130_fd_sc_hd__dfxtp_1
X_20553_ _33293_/Q _36173_/Q _33165_/Q _33101_/Q _18328_/X _19457_/A VGND VGND VPWR
+ VPWR _20553_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32539_ _35864_/CLK _32539_/D VGND VGND VPWR VPWR _32539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26060_ _26060_/A VGND VGND VPWR VPWR _33445_/D sky130_fd_sc_hd__clkbuf_1
X_35258_ _35578_/CLK _35258_/D VGND VGND VPWR VPWR _35258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23272_ _32208_/Q _23270_/X _23301_/S VGND VGND VPWR VPWR _23273_/A sky130_fd_sc_hd__mux2_1
X_20484_ _20484_/A VGND VGND VPWR VPWR _32138_/D sky130_fd_sc_hd__buf_4
XFILLER_146_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25011_ _25010_/X _32980_/Q _25020_/S VGND VGND VPWR VPWR _25012_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22223_ _22155_/X _22221_/X _22222_/X _22158_/X VGND VGND VPWR VPWR _22223_/X sky130_fd_sc_hd__a22o_1
X_34209_ _36123_/CLK _34209_/D VGND VGND VPWR VPWR _34209_/Q sky130_fd_sc_hd__dfxtp_1
X_35189_ _35315_/CLK _35189_/D VGND VGND VPWR VPWR _35189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22154_ _22148_/X _22151_/X _22152_/X _22153_/X VGND VGND VPWR VPWR _22154_/X sky130_fd_sc_hd__a22o_1
XTAP_6805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21105_ _32474_/Q _32346_/Q _32026_/Q _35994_/Q _20817_/X _20958_/X VGND VGND VPWR
+ VPWR _21105_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29750_ _35131_/Q _29191_/X _29758_/S VGND VGND VPWR VPWR _29751_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26962_ input40/X VGND VGND VPWR VPWR _26962_/X sky130_fd_sc_hd__clkbuf_4
X_22085_ _22008_/X _22083_/X _22084_/X _22014_/X VGND VGND VPWR VPWR _22085_/X sky130_fd_sc_hd__a22o_1
XFILLER_248_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_20_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _35226_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28701_ _26906_/X _34665_/Q _28705_/S VGND VGND VPWR VPWR _28702_/A sky130_fd_sc_hd__mux2_1
X_21036_ _35736_/Q _35096_/Q _34456_/Q _33816_/Q _21034_/X _21035_/X VGND VGND VPWR
+ VPWR _21036_/X sky130_fd_sc_hd__mux4_1
X_25913_ _25047_/X _33376_/Q _25915_/S VGND VGND VPWR VPWR _25914_/A sky130_fd_sc_hd__mux2_1
X_29681_ _35098_/Q _29089_/X _29695_/S VGND VGND VPWR VPWR _29682_/A sky130_fd_sc_hd__mux2_1
X_26893_ _26893_/A VGND VGND VPWR VPWR _33828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28632_ _28632_/A VGND VGND VPWR VPWR _34632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25844_ _25844_/A VGND VGND VPWR VPWR _33343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28563_ _28563_/A VGND VGND VPWR VPWR _34599_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22987_ _22987_/A VGND VGND VPWR VPWR _32048_/D sky130_fd_sc_hd__clkbuf_1
X_25775_ _25775_/A VGND VGND VPWR VPWR _33310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_1103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27514_ _26950_/X _34103_/Q _27530_/S VGND VGND VPWR VPWR _27515_/A sky130_fd_sc_hd__mux2_1
X_24726_ _24726_/A VGND VGND VPWR VPWR _32848_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21938_ _32754_/Q _32690_/Q _32626_/Q _36082_/Q _21872_/X _21656_/X VGND VGND VPWR
+ VPWR _21938_/X sky130_fd_sc_hd__mux4_1
X_28494_ _26999_/X _34567_/Q _28498_/S VGND VGND VPWR VPWR _28495_/A sky130_fd_sc_hd__mux2_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27445_ _27445_/A VGND VGND VPWR VPWR _34070_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24657_ _22988_/X _32817_/Q _24665_/S VGND VGND VPWR VPWR _24658_/A sky130_fd_sc_hd__mux2_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21869_ _34032_/Q _33968_/Q _33904_/Q _32240_/Q _21620_/X _21621_/X VGND VGND VPWR
+ VPWR _21869_/X sky130_fd_sc_hd__mux4_1
XFILLER_242_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_87_CLK clkbuf_leaf_87_CLK/A VGND VGND VPWR VPWR _35671_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23608_ _23608_/A VGND VGND VPWR VPWR _32354_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24588_ _22886_/X _32784_/Q _24602_/S VGND VGND VPWR VPWR _24589_/A sky130_fd_sc_hd__mux2_1
X_27376_ _27424_/S VGND VGND VPWR VPWR _27395_/S sky130_fd_sc_hd__buf_4
XFILLER_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29115_ _34850_/Q _29113_/X _29142_/S VGND VGND VPWR VPWR _29116_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23539_ _23044_/X _32323_/Q _23551_/S VGND VGND VPWR VPWR _23540_/A sky130_fd_sc_hd__mux2_1
X_26327_ _25060_/X _33572_/Q _26341_/S VGND VGND VPWR VPWR _26328_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17060_ _33258_/Q _36138_/Q _33130_/Q _33066_/Q _17058_/X _17059_/X VGND VGND VPWR
+ VPWR _17060_/X sky130_fd_sc_hd__mux4_1
X_29046_ _34829_/Q _24440_/X _29046_/S VGND VGND VPWR VPWR _29047_/A sky130_fd_sc_hd__mux2_1
X_26258_ _26258_/A VGND VGND VPWR VPWR _33539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16011_ _17834_/A VGND VGND VPWR VPWR _16011_/X sky130_fd_sc_hd__buf_2
XFILLER_6_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25209_ _25019_/X _33047_/Q _25209_/S VGND VGND VPWR VPWR _25210_/A sky130_fd_sc_hd__mux2_1
X_26189_ _26189_/A VGND VGND VPWR VPWR _33506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_15__f_CLK clkbuf_5_7_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_61_CLK/A sky130_fd_sc_hd__clkbuf_16
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _34819_/Q _34755_/Q _34691_/Q _34627_/Q _17641_/X _17642_/X VGND VGND VPWR
+ VPWR _17962_/X sky130_fd_sc_hd__mux4_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29948_ _29948_/A VGND VGND VPWR VPWR _35224_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_11_CLK clkbuf_6_3__f_CLK/X VGND VGND VPWR VPWR _35738_/CLK sky130_fd_sc_hd__clkbuf_16
X_19701_ _33780_/Q _33716_/Q _33652_/Q _33588_/Q _19496_/X _19497_/X VGND VGND VPWR
+ VPWR _19701_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16913_ _34278_/Q _34214_/Q _34150_/Q _34086_/Q _16736_/X _16737_/X VGND VGND VPWR
+ VPWR _16913_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17893_ _35329_/Q _35265_/Q _35201_/Q _32321_/Q _17712_/X _17713_/X VGND VGND VPWR
+ VPWR _17893_/X sky130_fd_sc_hd__mux4_1
X_29879_ _35192_/Q _29182_/X _29893_/S VGND VGND VPWR VPWR _29880_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31910_ _31910_/A VGND VGND VPWR VPWR _36154_/D sky130_fd_sc_hd__clkbuf_1
X_19632_ _34290_/Q _34226_/Q _34162_/Q _34098_/Q _19389_/X _19390_/X VGND VGND VPWR
+ VPWR _19632_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16844_ _17903_/A VGND VGND VPWR VPWR _16844_/X sky130_fd_sc_hd__clkbuf_4
X_32890_ _32954_/CLK _32890_/D VGND VGND VPWR VPWR _32890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31841_ _31841_/A VGND VGND VPWR VPWR _36121_/D sky130_fd_sc_hd__clkbuf_1
X_19563_ _19563_/A _19563_/B _19563_/C _19563_/D VGND VGND VPWR VPWR _19564_/A sky130_fd_sc_hd__or4_1
XFILLER_65_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16775_ _17834_/A VGND VGND VPWR VPWR _16775_/X sky130_fd_sc_hd__buf_2
XFILLER_98_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_1331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18514_ _32722_/Q _32658_/Q _32594_/Q _36050_/Q _18513_/X _20013_/A VGND VGND VPWR
+ VPWR _18514_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34560_ _35777_/CLK _34560_/D VGND VGND VPWR VPWR _34560_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31772_ _36089_/Q input38/X _31784_/S VGND VGND VPWR VPWR _31773_/A sky130_fd_sc_hd__mux2_1
X_19494_ _19494_/A VGND VGND VPWR VPWR _32109_/D sky130_fd_sc_hd__buf_2
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33511_ _33512_/CLK _33511_/D VGND VGND VPWR VPWR _33511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18445_ _34000_/Q _33936_/Q _33872_/Q _32144_/Q _18408_/X _18409_/X VGND VGND VPWR
+ VPWR _18445_/X sky130_fd_sc_hd__mux4_1
X_30723_ _35592_/Q _29231_/X _30725_/S VGND VGND VPWR VPWR _30724_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34491_ _35771_/CLK _34491_/D VGND VGND VPWR VPWR _34491_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_78_CLK clkbuf_leaf_80_CLK/A VGND VGND VPWR VPWR _35922_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_36230_ _36232_/CLK _36230_/D VGND VGND VPWR VPWR _36230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33442_ _33702_/CLK _33442_/D VGND VGND VPWR VPWR _33442_/Q sky130_fd_sc_hd__dfxtp_1
X_18376_ _20232_/A VGND VGND VPWR VPWR _18376_/X sky130_fd_sc_hd__buf_4
X_30654_ _35559_/Q _29129_/X _30662_/S VGND VGND VPWR VPWR _30655_/A sky130_fd_sc_hd__mux2_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36161_ _36161_/CLK _36161_/D VGND VGND VPWR VPWR _36161_/Q sky130_fd_sc_hd__dfxtp_1
X_17327_ _17154_/X _17325_/X _17326_/X _17159_/X VGND VGND VPWR VPWR _17327_/X sky130_fd_sc_hd__a22o_1
XFILLER_202_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33373_ _33946_/CLK _33373_/D VGND VGND VPWR VPWR _33373_/Q sky130_fd_sc_hd__dfxtp_1
X_30585_ _30585_/A VGND VGND VPWR VPWR _35526_/D sky130_fd_sc_hd__clkbuf_1
X_35112_ _35879_/CLK _35112_/D VGND VGND VPWR VPWR _35112_/Q sky130_fd_sc_hd__dfxtp_1
X_32324_ _35332_/CLK _32324_/D VGND VGND VPWR VPWR _32324_/Q sky130_fd_sc_hd__dfxtp_1
X_36092_ _36092_/CLK _36092_/D VGND VGND VPWR VPWR _36092_/Q sky130_fd_sc_hd__dfxtp_1
X_17258_ _17149_/X _17256_/X _17257_/X _17152_/X VGND VGND VPWR VPWR _17258_/X sky130_fd_sc_hd__a22o_1
XFILLER_70_1280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16209_ _33490_/Q _33426_/Q _33362_/Q _33298_/Q _15998_/X _15999_/X VGND VGND VPWR
+ VPWR _16209_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35043_ _35299_/CLK _35043_/D VGND VGND VPWR VPWR _35043_/Q sky130_fd_sc_hd__dfxtp_1
X_32255_ _34046_/CLK _32255_/D VGND VGND VPWR VPWR _32255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17189_ _34541_/Q _32429_/Q _34413_/Q _34349_/Q _16872_/X _16873_/X VGND VGND VPWR
+ VPWR _17189_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31206_ _31206_/A VGND VGND VPWR VPWR _35820_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32186_ _35748_/CLK _32186_/D VGND VGND VPWR VPWR _32186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31137_ _31137_/A VGND VGND VPWR VPWR _35788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35945_ _35945_/CLK _35945_/D VGND VGND VPWR VPWR _35945_/Q sky130_fd_sc_hd__dfxtp_1
X_31068_ _31068_/A VGND VGND VPWR VPWR _35755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22910_ input2/X VGND VGND VPWR VPWR _22910_/X sky130_fd_sc_hd__buf_4
XFILLER_151_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30019_ _30019_/A VGND VGND VPWR VPWR _35258_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35876_ _35876_/CLK _35876_/D VGND VGND VPWR VPWR _35876_/Q sky130_fd_sc_hd__dfxtp_1
X_23890_ _23890_/A VGND VGND VPWR VPWR _32486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_1087 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34827_ _35147_/CLK _34827_/D VGND VGND VPWR VPWR _34827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22841_ _20656_/X _22839_/X _22840_/X _20668_/X VGND VGND VPWR VPWR _22841_/X sky130_fd_sc_hd__a22o_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25560_ _33211_/Q _24385_/X _25568_/S VGND VGND VPWR VPWR _25561_/A sky130_fd_sc_hd__mux2_1
X_34758_ _34822_/CLK _34758_/D VGND VGND VPWR VPWR _34758_/Q sky130_fd_sc_hd__dfxtp_1
X_22772_ _35594_/Q _35530_/Q _35466_/Q _35402_/Q _22556_/X _22557_/X VGND VGND VPWR
+ VPWR _22772_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24511_ _22976_/X _32749_/Q _24527_/S VGND VGND VPWR VPWR _24512_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21723_ _22429_/A VGND VGND VPWR VPWR _21723_/X sky130_fd_sc_hd__buf_4
X_33709_ _34745_/CLK _33709_/D VGND VGND VPWR VPWR _33709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25491_ _33178_/Q _24283_/X _25505_/S VGND VGND VPWR VPWR _25492_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34689_ _35328_/CLK _34689_/D VGND VGND VPWR VPWR _34689_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_69_CLK clkbuf_leaf_73_CLK/A VGND VGND VPWR VPWR _36119_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24442_ _24442_/A VGND VGND VPWR VPWR _32717_/D sky130_fd_sc_hd__clkbuf_1
X_27230_ _27230_/A VGND VGND VPWR VPWR _33968_/D sky130_fd_sc_hd__clkbuf_1
X_21654_ _21650_/X _21653_/X _21375_/X VGND VGND VPWR VPWR _21686_/A sky130_fd_sc_hd__o21ba_1
XFILLER_244_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27161_ _27161_/A VGND VGND VPWR VPWR _33935_/D sky130_fd_sc_hd__clkbuf_1
X_20605_ _22556_/A VGND VGND VPWR VPWR _20605_/X sky130_fd_sc_hd__buf_6
XFILLER_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24373_ input36/X VGND VGND VPWR VPWR _24373_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_193_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21585_ _32744_/Q _32680_/Q _32616_/Q _36072_/Q _21519_/X _21303_/X VGND VGND VPWR
+ VPWR _21585_/X sky130_fd_sc_hd__mux4_1
XFILLER_228_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26112_ _26112_/A VGND VGND VPWR VPWR _33470_/D sky130_fd_sc_hd__clkbuf_1
X_23324_ _23324_/A VGND VGND VPWR VPWR _32225_/D sky130_fd_sc_hd__clkbuf_1
X_20536_ _34828_/Q _34764_/Q _34700_/Q _34636_/Q _20294_/X _20295_/X VGND VGND VPWR
+ VPWR _20536_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27092_ _26925_/X _33903_/Q _27104_/S VGND VGND VPWR VPWR _27093_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26043_ _26043_/A VGND VGND VPWR VPWR _33437_/D sky130_fd_sc_hd__clkbuf_1
X_23255_ _23255_/A VGND VGND VPWR VPWR _32202_/D sky130_fd_sc_hd__clkbuf_1
X_20467_ _19454_/A _20465_/X _20466_/X _19459_/A VGND VGND VPWR VPWR _20467_/X sky130_fd_sc_hd__a22o_1
XFILLER_165_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22206_ _33209_/Q _32569_/Q _35961_/Q _35897_/Q _22027_/X _22028_/X VGND VGND VPWR
+ VPWR _22206_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23186_ _23186_/A VGND VGND VPWR VPWR _32175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20398_ _33544_/Q _33480_/Q _33416_/Q _33352_/Q _20129_/X _20130_/X VGND VGND VPWR
+ VPWR _20398_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_5_3_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_3_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XTAP_6602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29802_ _29802_/A VGND VGND VPWR VPWR _35155_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22137_ _21952_/X _22135_/X _22136_/X _21955_/X VGND VGND VPWR VPWR _22137_/X sky130_fd_sc_hd__a22o_1
XTAP_6624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput280 _32086_/Q VGND VGND VPWR VPWR D3[8] sky130_fd_sc_hd__buf_2
X_27994_ _27994_/A VGND VGND VPWR VPWR _34329_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29733_ _35123_/Q _29166_/X _29737_/S VGND VGND VPWR VPWR _29734_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22068_ _35061_/Q _34997_/Q _34933_/Q _34869_/Q _21756_/X _21757_/X VGND VGND VPWR
+ VPWR _22068_/X sky130_fd_sc_hd__mux4_1
X_26945_ _26945_/A VGND VGND VPWR VPWR _33845_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21019_ _33496_/Q _33432_/Q _33368_/Q _33304_/Q _21017_/X _21018_/X VGND VGND VPWR
+ VPWR _21019_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29664_ _35090_/Q _29064_/X _29674_/S VGND VGND VPWR VPWR _29665_/A sky130_fd_sc_hd__mux2_1
XTAP_5978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26876_ _26875_/X _33823_/Q _26882_/S VGND VGND VPWR VPWR _26877_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28615_ _26977_/X _34624_/Q _28633_/S VGND VGND VPWR VPWR _28616_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25827_ _25119_/X _33335_/Q _25843_/S VGND VGND VPWR VPWR _25828_/A sky130_fd_sc_hd__mux2_1
X_29595_ _29595_/A VGND VGND VPWR VPWR _35057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28546_ _28546_/A VGND VGND VPWR VPWR _34591_/D sky130_fd_sc_hd__clkbuf_1
X_16560_ _34268_/Q _34204_/Q _34140_/Q _34076_/Q _16383_/X _16384_/X VGND VGND VPWR
+ VPWR _16560_/X sky130_fd_sc_hd__mux4_1
X_25758_ _25758_/A VGND VGND VPWR VPWR _33302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24709_ _23065_/X _32842_/Q _24715_/S VGND VGND VPWR VPWR _24710_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28477_ _26974_/X _34559_/Q _28477_/S VGND VGND VPWR VPWR _28478_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16491_ _17903_/A VGND VGND VPWR VPWR _16491_/X sky130_fd_sc_hd__buf_4
XFILLER_203_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25689_ _25689_/A VGND VGND VPWR VPWR _33270_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18230_ _35788_/Q _35148_/Q _34508_/Q _33868_/Q _16108_/X _16109_/X VGND VGND VPWR
+ VPWR _18230_/X sky130_fd_sc_hd__mux4_1
X_27428_ _26821_/X _34062_/Q _27446_/S VGND VGND VPWR VPWR _27429_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_0_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _35036_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18161_ _18157_/X _18160_/X _17834_/A VGND VGND VPWR VPWR _18183_/A sky130_fd_sc_hd__o21ba_1
XFILLER_12_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27359_ _27359_/A VGND VGND VPWR VPWR _34029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17112_ _35307_/Q _35243_/Q _35179_/Q _32299_/Q _17006_/X _17007_/X VGND VGND VPWR
+ VPWR _17112_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18092_ _18088_/X _18091_/X _17867_/X VGND VGND VPWR VPWR _18093_/D sky130_fd_sc_hd__o21ba_1
X_30370_ _30370_/A VGND VGND VPWR VPWR _35424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29029_ _29029_/A VGND VGND VPWR VPWR _34820_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17043_ _35049_/Q _34985_/Q _34921_/Q _34857_/Q _16803_/X _16804_/X VGND VGND VPWR
+ VPWR _17043_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32040_ _36072_/CLK _32040_/D VGND VGND VPWR VPWR _32040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1043 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18994_ _18994_/A VGND VGND VPWR VPWR _32095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _17941_/X _17944_/X _17834_/X VGND VGND VPWR VPWR _17969_/A sky130_fd_sc_hd__o21ba_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33991_ _34816_/CLK _33991_/D VGND VGND VPWR VPWR _33991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35730_ _35730_/CLK _35730_/D VGND VGND VPWR VPWR _35730_/Q sky130_fd_sc_hd__dfxtp_1
X_32942_ _33007_/CLK _32942_/D VGND VGND VPWR VPWR _32942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17876_ _17555_/X _17874_/X _17875_/X _17558_/X VGND VGND VPWR VPWR _17876_/X sky130_fd_sc_hd__a22o_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19615_ _35825_/Q _32202_/Q _35697_/Q _35633_/Q _19613_/X _19614_/X VGND VGND VPWR
+ VPWR _19615_/X sky130_fd_sc_hd__mux4_1
X_35661_ _35789_/CLK _35661_/D VGND VGND VPWR VPWR _35661_/Q sky130_fd_sc_hd__dfxtp_1
X_16827_ _35747_/Q _35107_/Q _34467_/Q _33827_/Q _16787_/X _16788_/X VGND VGND VPWR
+ VPWR _16827_/X sky130_fd_sc_hd__mux4_1
X_32873_ _36009_/CLK _32873_/D VGND VGND VPWR VPWR _32873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_998 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34612_ _35187_/CLK _34612_/D VGND VGND VPWR VPWR _34612_/Q sky130_fd_sc_hd__dfxtp_1
X_31824_ _31824_/A VGND VGND VPWR VPWR _36113_/D sky130_fd_sc_hd__clkbuf_1
X_19546_ _19542_/X _19545_/X _19436_/X _19437_/X VGND VGND VPWR VPWR _19563_/B sky130_fd_sc_hd__o211a_1
X_35592_ _35849_/CLK _35592_/D VGND VGND VPWR VPWR _35592_/Q sky130_fd_sc_hd__dfxtp_1
X_16758_ _34785_/Q _34721_/Q _34657_/Q _34593_/Q _16582_/X _16583_/X VGND VGND VPWR
+ VPWR _16758_/X sky130_fd_sc_hd__mux4_1
XFILLER_207_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34543_ _35954_/CLK _34543_/D VGND VGND VPWR VPWR _34543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31755_ _36081_/Q input29/X _31763_/S VGND VGND VPWR VPWR _31756_/A sky130_fd_sc_hd__mux2_1
X_19477_ _19363_/X _19475_/X _19476_/X _19367_/X VGND VGND VPWR VPWR _19477_/X sky130_fd_sc_hd__a22o_1
XFILLER_206_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16689_ _34527_/Q _32415_/Q _34399_/Q _34335_/Q _16519_/X _16520_/X VGND VGND VPWR
+ VPWR _16689_/X sky130_fd_sc_hd__mux4_1
XFILLER_222_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30706_ _30733_/S VGND VGND VPWR VPWR _30725_/S sky130_fd_sc_hd__buf_4
X_18428_ _35279_/Q _35215_/Q _35151_/Q _32271_/Q _18379_/X _18381_/X VGND VGND VPWR
+ VPWR _18428_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34474_ _35945_/CLK _34474_/D VGND VGND VPWR VPWR _34474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31686_ _36048_/Q input23/X _31700_/S VGND VGND VPWR VPWR _31687_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36213_ _36216_/CLK _36213_/D VGND VGND VPWR VPWR _36213_/Q sky130_fd_sc_hd__dfxtp_1
X_33425_ _36232_/CLK _33425_/D VGND VGND VPWR VPWR _33425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18359_ _18359_/A VGND VGND VPWR VPWR _20147_/A sky130_fd_sc_hd__buf_12
X_30637_ _35551_/Q _29104_/X _30641_/S VGND VGND VPWR VPWR _30638_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36144_ _36146_/CLK _36144_/D VGND VGND VPWR VPWR _36144_/Q sky130_fd_sc_hd__dfxtp_1
X_33356_ _33548_/CLK _33356_/D VGND VGND VPWR VPWR _33356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21370_ _22429_/A VGND VGND VPWR VPWR _21370_/X sky130_fd_sc_hd__buf_4
X_30568_ _30568_/A VGND VGND VPWR VPWR _35518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20321_ _20000_/X _20319_/X _20320_/X _20003_/X VGND VGND VPWR VPWR _20321_/X sky130_fd_sc_hd__a22o_1
X_32307_ _35700_/CLK _32307_/D VGND VGND VPWR VPWR _32307_/Q sky130_fd_sc_hd__dfxtp_1
X_36075_ _36075_/CLK _36075_/D VGND VGND VPWR VPWR _36075_/Q sky130_fd_sc_hd__dfxtp_1
X_33287_ _36167_/CLK _33287_/D VGND VGND VPWR VPWR _33287_/Q sky130_fd_sc_hd__dfxtp_1
X_30499_ _30499_/A VGND VGND VPWR VPWR _35485_/D sky130_fd_sc_hd__clkbuf_1
X_35026_ _35026_/CLK _35026_/D VGND VGND VPWR VPWR _35026_/Q sky130_fd_sc_hd__dfxtp_1
X_23040_ _23040_/A VGND VGND VPWR VPWR _32065_/D sky130_fd_sc_hd__clkbuf_1
X_20252_ _20248_/X _20251_/X _20142_/X _20143_/X VGND VGND VPWR VPWR _20269_/B sky130_fd_sc_hd__o211a_1
X_32238_ _34032_/CLK _32238_/D VGND VGND VPWR VPWR _32238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20183_ _20069_/X _20181_/X _20182_/X _20073_/X VGND VGND VPWR VPWR _20183_/X sky130_fd_sc_hd__a22o_1
X_32169_ _35797_/CLK _32169_/D VGND VGND VPWR VPWR _32169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_61__f_CLK clkbuf_5_30_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_61__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_24991_ _31815_/B _28373_/B VGND VGND VPWR VPWR _25187_/S sky130_fd_sc_hd__nand2_8
XTAP_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26730_ _33762_/Q _24307_/X _26748_/S VGND VGND VPWR VPWR _26731_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23942_ _23942_/A VGND VGND VPWR VPWR _32511_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35928_ _35928_/CLK _35928_/D VGND VGND VPWR VPWR _35928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26661_ _25153_/X _33730_/Q _26675_/S VGND VGND VPWR VPWR _26662_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23873_ _23873_/A VGND VGND VPWR VPWR _32478_/D sky130_fd_sc_hd__clkbuf_1
X_35859_ _35925_/CLK _35859_/D VGND VGND VPWR VPWR _35859_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28400_ _26860_/X _34522_/Q _28414_/S VGND VGND VPWR VPWR _28401_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22824_ _21749_/A _22822_/X _22823_/X _21752_/A VGND VGND VPWR VPWR _22824_/X sky130_fd_sc_hd__a22o_1
X_25612_ _33234_/Q _24258_/X _25622_/S VGND VGND VPWR VPWR _25613_/A sky130_fd_sc_hd__mux2_1
XANTENNA_806 _22898_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29380_ _23342_/X _34956_/Q _29382_/S VGND VGND VPWR VPWR _29381_/A sky130_fd_sc_hd__mux2_1
XANTENNA_817 _22938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26592_ _26592_/A VGND VGND VPWR VPWR _33697_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_828 _23124_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_839 _23294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_213_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28331_ _28331_/A VGND VGND VPWR VPWR _34489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22755_ _33802_/Q _33738_/Q _33674_/Q _33610_/Q _22502_/X _22503_/X VGND VGND VPWR
+ VPWR _22755_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25543_ _33203_/Q _24360_/X _25547_/S VGND VGND VPWR VPWR _25544_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21706_ _21594_/X _21704_/X _21705_/X _21597_/X VGND VGND VPWR VPWR _21706_/X sky130_fd_sc_hd__a22o_1
X_25474_ _33170_/Q _24258_/X _25484_/S VGND VGND VPWR VPWR _25475_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28262_ _28262_/A VGND VGND VPWR VPWR _34456_/D sky130_fd_sc_hd__clkbuf_1
X_22686_ _34823_/Q _34759_/Q _34695_/Q _34631_/Q _22594_/X _22595_/X VGND VGND VPWR
+ VPWR _22686_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24425_ input54/X VGND VGND VPWR VPWR _24425_/X sky130_fd_sc_hd__clkbuf_8
X_27213_ _27213_/A VGND VGND VPWR VPWR _33960_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21637_ _21599_/X _21635_/X _21636_/X _21602_/X VGND VGND VPWR VPWR _21637_/X sky130_fd_sc_hd__a22o_1
X_28193_ _26953_/X _34424_/Q _28207_/S VGND VGND VPWR VPWR _28194_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27144_ _27002_/X _33928_/Q _27146_/S VGND VGND VPWR VPWR _27145_/A sky130_fd_sc_hd__mux2_1
X_24356_ _24356_/A VGND VGND VPWR VPWR _32689_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21568_ _21564_/X _21567_/X _21394_/X VGND VGND VPWR VPWR _21576_/C sky130_fd_sc_hd__o21ba_1
XFILLER_219_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23307_ input47/X VGND VGND VPWR VPWR _23307_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_165_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20519_ _34060_/Q _33996_/Q _33932_/Q _32268_/Q _18358_/X _18360_/X VGND VGND VPWR
+ VPWR _20519_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27075_ _26900_/X _33895_/Q _27083_/S VGND VGND VPWR VPWR _27076_/A sky130_fd_sc_hd__mux2_1
X_24287_ _32667_/Q _24286_/X _24305_/S VGND VGND VPWR VPWR _24288_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21499_ _35557_/Q _35493_/Q _35429_/Q _35365_/Q _21497_/X _21498_/X VGND VGND VPWR
+ VPWR _21499_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26026_ _26026_/A VGND VGND VPWR VPWR _33429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23238_ _23346_/S VGND VGND VPWR VPWR _23268_/S sky130_fd_sc_hd__buf_6
XFILLER_107_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23169_ _32168_/Q _23099_/X _23182_/S VGND VGND VPWR VPWR _23170_/A sky130_fd_sc_hd__mux2_1
XTAP_6421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1205 _23133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1216 _23696_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1227 _24429_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1238 _25597_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ _17796_/A VGND VGND VPWR VPWR _15991_/X sky130_fd_sc_hd__buf_4
XTAP_5720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1249 _26683_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27977_ _27977_/A VGND VGND VPWR VPWR _34321_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17730_ _17724_/X _17729_/X _17481_/X VGND VGND VPWR VPWR _17752_/A sky130_fd_sc_hd__o21ba_1
XFILLER_121_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29716_ _35115_/Q _29141_/X _29716_/S VGND VGND VPWR VPWR _29717_/A sky130_fd_sc_hd__mux2_1
XTAP_6498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26928_ input28/X VGND VGND VPWR VPWR _26928_/X sky130_fd_sc_hd__buf_4
XFILLER_47_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29647_ _29647_/A VGND VGND VPWR VPWR _35082_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17661_ _17408_/X _17659_/X _17660_/X _17414_/X VGND VGND VPWR VPWR _17661_/X sky130_fd_sc_hd__a22o_1
XFILLER_236_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26859_ _26859_/A VGND VGND VPWR VPWR _33817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19400_ _32491_/Q _32363_/Q _32043_/Q _36011_/Q _19223_/X _19364_/X VGND VGND VPWR
+ VPWR _19400_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16612_ _35549_/Q _35485_/Q _35421_/Q _35357_/Q _16544_/X _16545_/X VGND VGND VPWR
+ VPWR _16612_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17592_ _17588_/X _17591_/X _17481_/X VGND VGND VPWR VPWR _17616_/A sky130_fd_sc_hd__o21ba_1
X_29578_ _29578_/A VGND VGND VPWR VPWR _35049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19331_ _19327_/X _19330_/X _19083_/X _19084_/X VGND VGND VPWR VPWR _19346_/B sky130_fd_sc_hd__o211a_1
X_28529_ _28529_/A VGND VGND VPWR VPWR _34583_/D sky130_fd_sc_hd__clkbuf_1
X_16543_ _16288_/X _16541_/X _16542_/X _16291_/X VGND VGND VPWR VPWR _16543_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31540_ _31540_/A VGND VGND VPWR VPWR _35979_/D sky130_fd_sc_hd__clkbuf_1
X_19262_ _35815_/Q _32191_/Q _35687_/Q _35623_/Q _19260_/X _19261_/X VGND VGND VPWR
+ VPWR _19262_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16474_ _35737_/Q _35097_/Q _34457_/Q _33817_/Q _16434_/X _16435_/X VGND VGND VPWR
+ VPWR _16474_/X sky130_fd_sc_hd__mux4_1
XFILLER_245_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18213_ _18213_/A _18213_/B _18213_/C _18213_/D VGND VGND VPWR VPWR _18214_/A sky130_fd_sc_hd__or4_4
XFILLER_188_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31471_ _31471_/A VGND VGND VPWR VPWR _35946_/D sky130_fd_sc_hd__clkbuf_1
X_19193_ _19189_/X _19192_/X _19083_/X _19084_/X VGND VGND VPWR VPWR _19210_/B sky130_fd_sc_hd__o211a_1
XFILLER_31_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33210_ _36027_/CLK _33210_/D VGND VGND VPWR VPWR _33210_/Q sky130_fd_sc_hd__dfxtp_1
X_18144_ _15997_/X _18142_/X _18143_/X _16003_/X VGND VGND VPWR VPWR _18144_/X sky130_fd_sc_hd__a22o_1
X_30422_ _23280_/X _35449_/Q _30434_/S VGND VGND VPWR VPWR _30423_/A sky130_fd_sc_hd__mux2_1
X_34190_ _34256_/CLK _34190_/D VGND VGND VPWR VPWR _34190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33141_ _36086_/CLK _33141_/D VGND VGND VPWR VPWR _33141_/Q sky130_fd_sc_hd__dfxtp_1
X_18075_ _32519_/Q _32391_/Q _32071_/Q _36039_/Q _17982_/X _17770_/X VGND VGND VPWR
+ VPWR _18075_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30353_ _23117_/X _35416_/Q _30371_/S VGND VGND VPWR VPWR _30354_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17026_ _33257_/Q _36137_/Q _33129_/Q _33065_/Q _16705_/X _16706_/X VGND VGND VPWR
+ VPWR _17026_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33072_ _36081_/CLK _33072_/D VGND VGND VPWR VPWR _33072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30284_ _35384_/Q _29182_/X _30298_/S VGND VGND VPWR VPWR _30285_/A sky130_fd_sc_hd__mux2_1
XFILLER_236_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32023_ _33507_/CLK _32023_/D VGND VGND VPWR VPWR _32023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _18657_/X _18975_/X _18976_/X _18661_/X VGND VGND VPWR VPWR _18977_/X sky130_fd_sc_hd__a22o_1
XFILLER_6_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _34818_/Q _34754_/Q _34690_/Q _34626_/Q _17641_/X _17642_/X VGND VGND VPWR
+ VPWR _17928_/X sky130_fd_sc_hd__mux4_1
XFILLER_234_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33974_ _36152_/CLK _33974_/D VGND VGND VPWR VPWR _33974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35713_ _35715_/CLK _35713_/D VGND VGND VPWR VPWR _35713_/Q sky130_fd_sc_hd__dfxtp_1
X_32925_ _34146_/CLK _32925_/D VGND VGND VPWR VPWR _32925_/Q sky130_fd_sc_hd__dfxtp_1
X_17859_ _17855_/X _17856_/X _17857_/X _17858_/X VGND VGND VPWR VPWR _17859_/X sky130_fd_sc_hd__a22o_1
XFILLER_27_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20870_ _20870_/A _20870_/B _20870_/C _20870_/D VGND VGND VPWR VPWR _20871_/A sky130_fd_sc_hd__or4_2
X_35644_ _35965_/CLK _35644_/D VGND VGND VPWR VPWR _35644_/Q sky130_fd_sc_hd__dfxtp_1
X_32856_ _35994_/CLK _32856_/D VGND VGND VPWR VPWR _32856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31807_ _36106_/Q input57/X _31813_/S VGND VGND VPWR VPWR _31808_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19529_ _19454_/X _19527_/X _19528_/X _19459_/X VGND VGND VPWR VPWR _19529_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35575_ _35575_/CLK _35575_/D VGND VGND VPWR VPWR _35575_/Q sky130_fd_sc_hd__dfxtp_1
X_32787_ _32978_/CLK _32787_/D VGND VGND VPWR VPWR _32787_/Q sky130_fd_sc_hd__dfxtp_1
X_22540_ _34307_/Q _34243_/Q _34179_/Q _34115_/Q _22395_/X _22396_/X VGND VGND VPWR
+ VPWR _22540_/X sky130_fd_sc_hd__mux4_1
X_34526_ _35038_/CLK _34526_/D VGND VGND VPWR VPWR _34526_/Q sky130_fd_sc_hd__dfxtp_1
X_31738_ _36073_/Q input20/X _31742_/S VGND VGND VPWR VPWR _31739_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_1431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22471_ _33793_/Q _33729_/Q _33665_/Q _33601_/Q _22149_/X _22150_/X VGND VGND VPWR
+ VPWR _22471_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34457_ _35803_/CLK _34457_/D VGND VGND VPWR VPWR _34457_/Q sky130_fd_sc_hd__dfxtp_1
X_31669_ _31669_/A VGND VGND VPWR VPWR _36040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24210_ _24210_/A VGND VGND VPWR VPWR _32637_/D sky130_fd_sc_hd__clkbuf_1
X_33408_ _34305_/CLK _33408_/D VGND VGND VPWR VPWR _33408_/Q sky130_fd_sc_hd__dfxtp_1
X_21422_ _32483_/Q _32355_/Q _32035_/Q _36003_/Q _21170_/X _21311_/X VGND VGND VPWR
+ VPWR _21422_/X sky130_fd_sc_hd__mux4_1
XFILLER_202_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25190_ _25322_/S VGND VGND VPWR VPWR _25209_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_175_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34388_ _34706_/CLK _34388_/D VGND VGND VPWR VPWR _34388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24141_ _24141_/A VGND VGND VPWR VPWR _32604_/D sky130_fd_sc_hd__clkbuf_1
X_36127_ _36127_/CLK _36127_/D VGND VGND VPWR VPWR _36127_/Q sky130_fd_sc_hd__dfxtp_1
X_33339_ _33723_/CLK _33339_/D VGND VGND VPWR VPWR _33339_/Q sky130_fd_sc_hd__dfxtp_1
X_21353_ _21241_/X _21351_/X _21352_/X _21244_/X VGND VGND VPWR VPWR _21353_/X sky130_fd_sc_hd__a22o_1
XFILLER_194_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20304_ _20304_/A VGND VGND VPWR VPWR _32132_/D sky130_fd_sc_hd__buf_4
XFILLER_135_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24072_ _24072_/A VGND VGND VPWR VPWR _32572_/D sky130_fd_sc_hd__clkbuf_1
X_36058_ _36121_/CLK _36058_/D VGND VGND VPWR VPWR _36058_/Q sky130_fd_sc_hd__dfxtp_1
X_21284_ _21246_/X _21282_/X _21283_/X _21249_/X VGND VGND VPWR VPWR _21284_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35009_ _35075_/CLK _35009_/D VGND VGND VPWR VPWR _35009_/Q sky130_fd_sc_hd__dfxtp_1
X_23023_ _23022_/X _32060_/Q _23032_/S VGND VGND VPWR VPWR _23024_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27900_ _34285_/Q _24342_/X _27916_/S VGND VGND VPWR VPWR _27901_/A sky130_fd_sc_hd__mux2_1
X_20235_ _20160_/X _20233_/X _20234_/X _20165_/X VGND VGND VPWR VPWR _20235_/X sky130_fd_sc_hd__a22o_1
X_28880_ _26971_/X _34750_/Q _28882_/S VGND VGND VPWR VPWR _28881_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27831_ _34253_/Q _24440_/X _27831_/S VGND VGND VPWR VPWR _27832_/A sky130_fd_sc_hd__mux2_1
XTAP_5005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20166_ _20160_/X _20161_/X _20164_/X _20165_/X VGND VGND VPWR VPWR _20166_/X sky130_fd_sc_hd__a22o_1
XTAP_5016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27762_ _27831_/S VGND VGND VPWR VPWR _27781_/S sky130_fd_sc_hd__buf_6
X_24974_ _24974_/A VGND VGND VPWR VPWR _32966_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20097_ _34303_/Q _34239_/Q _34175_/Q _34111_/Q _20095_/X _20096_/X VGND VGND VPWR
+ VPWR _20097_/X sky130_fd_sc_hd__mux4_1
XTAP_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29501_ _23319_/X _35013_/Q _29509_/S VGND VGND VPWR VPWR _29502_/A sky130_fd_sc_hd__mux2_1
XFILLER_218_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26713_ _33754_/Q _24283_/X _26727_/S VGND VGND VPWR VPWR _26714_/A sky130_fd_sc_hd__mux2_1
XTAP_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23925_ _23007_/X _32503_/Q _23941_/S VGND VGND VPWR VPWR _23926_/A sky130_fd_sc_hd__mux2_1
X_27693_ _27693_/A VGND VGND VPWR VPWR _34187_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29432_ _23175_/X _34980_/Q _29446_/S VGND VGND VPWR VPWR _29433_/A sky130_fd_sc_hd__mux2_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_603 _20167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26644_ _25128_/X _33722_/Q _26654_/S VGND VGND VPWR VPWR _26645_/A sky130_fd_sc_hd__mux2_1
XTAP_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23856_ _23856_/A VGND VGND VPWR VPWR _32470_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_614 _18505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_625 _18681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_636 _19141_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22807_ _35339_/Q _35275_/Q _35211_/Q _32331_/Q _20688_/X _20690_/X VGND VGND VPWR
+ VPWR _22807_/X sky130_fd_sc_hd__mux4_1
X_29363_ _29363_/A VGND VGND VPWR VPWR _34947_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_647 _19629_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_658 _20363_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26575_ _25026_/X _33689_/Q _26591_/S VGND VGND VPWR VPWR _26576_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20999_ _35735_/Q _35095_/Q _34455_/Q _33815_/Q _20649_/X _20651_/X VGND VGND VPWR
+ VPWR _20999_/X sky130_fd_sc_hd__mux4_1
XANTENNA_669 _22460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23787_ _23003_/X _32438_/Q _23805_/S VGND VGND VPWR VPWR _23788_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28314_ _28314_/A VGND VGND VPWR VPWR _34481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25526_ _33195_/Q _24335_/X _25526_/S VGND VGND VPWR VPWR _25527_/A sky130_fd_sc_hd__mux2_1
X_22738_ _22734_/X _22737_/X _22442_/X _22443_/X VGND VGND VPWR VPWR _22753_/B sky130_fd_sc_hd__o211a_1
X_29294_ _29294_/A VGND VGND VPWR VPWR _34914_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28245_ _28245_/A VGND VGND VPWR VPWR _34448_/D sky130_fd_sc_hd__clkbuf_1
X_22669_ _34055_/Q _33991_/Q _33927_/Q _32263_/Q _20658_/X _20660_/X VGND VGND VPWR
+ VPWR _22669_/X sky130_fd_sc_hd__mux4_1
X_25457_ _25457_/A VGND VGND VPWR VPWR _33164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24408_ _32706_/Q _24407_/X _24429_/S VGND VGND VPWR VPWR _24409_/A sky130_fd_sc_hd__mux2_1
X_16190_ _16044_/X _16188_/X _16189_/X _16054_/X VGND VGND VPWR VPWR _16190_/X sky130_fd_sc_hd__a22o_1
X_28176_ _26928_/X _34416_/Q _28186_/S VGND VGND VPWR VPWR _28177_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25388_ _25388_/A VGND VGND VPWR VPWR _33131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27127_ _27154_/S VGND VGND VPWR VPWR _27146_/S sky130_fd_sc_hd__buf_4
XFILLER_153_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24339_ _24401_/A VGND VGND VPWR VPWR _24367_/S sky130_fd_sc_hd__buf_4
XFILLER_153_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27058_ _26875_/X _33887_/Q _27062_/S VGND VGND VPWR VPWR _27059_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18900_ _32733_/Q _32669_/Q _32605_/Q _36061_/Q _18866_/X _18650_/X VGND VGND VPWR
+ VPWR _18900_/X sky130_fd_sc_hd__mux4_1
X_26009_ _30465_/B _26685_/B VGND VGND VPWR VPWR _26142_/S sky130_fd_sc_hd__nand2_8
X_19880_ _34552_/Q _32440_/Q _34424_/Q _34360_/Q _19878_/X _19879_/X VGND VGND VPWR
+ VPWR _19880_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1002 _17834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18831_ _34011_/Q _33947_/Q _33883_/Q _32155_/Q _18614_/X _18615_/X VGND VGND VPWR
+ VPWR _18831_/X sky130_fd_sc_hd__mux4_1
XANTENNA_1013 _17842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1024 _17865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1035 _17149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1046 _17159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1057 _16457_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18762_ _33497_/Q _33433_/Q _33369_/Q _33305_/Q _18717_/X _18718_/X VGND VGND VPWR
+ VPWR _18762_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1068 _17119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1079 _17194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17713_ _17713_/A VGND VGND VPWR VPWR _17713_/X sky130_fd_sc_hd__buf_6
XFILLER_62_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30971_ _30971_/A VGND VGND VPWR VPWR _35709_/D sky130_fd_sc_hd__clkbuf_1
X_18693_ _18649_/X _18691_/X _18692_/X _18655_/X VGND VGND VPWR VPWR _18693_/X sky130_fd_sc_hd__a22o_1
XFILLER_29_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32710_ _36103_/CLK _32710_/D VGND VGND VPWR VPWR _32710_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_291_CLK clkbuf_6_57__f_CLK/X VGND VGND VPWR VPWR _36031_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_1339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17644_ _35322_/Q _35258_/Q _35194_/Q _32314_/Q _17359_/X _17360_/X VGND VGND VPWR
+ VPWR _17644_/X sky130_fd_sc_hd__mux4_1
XTAP_4893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33690_ _33692_/CLK _33690_/D VGND VGND VPWR VPWR _33690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32641_ _36098_/CLK _32641_/D VGND VGND VPWR VPWR _32641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17575_ _34808_/Q _34744_/Q _34680_/Q _34616_/Q _17288_/X _17289_/X VGND VGND VPWR
+ VPWR _17575_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19314_ _19314_/A _19314_/B _19314_/C _19314_/D VGND VGND VPWR VPWR _19315_/A sky130_fd_sc_hd__or4_4
XFILLER_188_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16526_ _16526_/A VGND VGND VPWR VPWR _31962_/D sky130_fd_sc_hd__clkbuf_1
X_35360_ _35744_/CLK _35360_/D VGND VGND VPWR VPWR _35360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32572_ _36028_/CLK _32572_/D VGND VGND VPWR VPWR _32572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_1224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34311_ _34817_/CLK _34311_/D VGND VGND VPWR VPWR _34311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31523_ _23313_/X _35971_/Q _31535_/S VGND VGND VPWR VPWR _31524_/A sky130_fd_sc_hd__mux2_1
X_19245_ _19245_/A VGND VGND VPWR VPWR _32102_/D sky130_fd_sc_hd__clkbuf_1
X_16457_ _16457_/A _16457_/B _16457_/C _16457_/D VGND VGND VPWR VPWR _16458_/A sky130_fd_sc_hd__or4_2
X_35291_ _35293_/CLK _35291_/D VGND VGND VPWR VPWR _35291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34242_ _34243_/CLK _34242_/D VGND VGND VPWR VPWR _34242_/Q sky130_fd_sc_hd__dfxtp_1
X_31454_ _23148_/X _35938_/Q _31472_/S VGND VGND VPWR VPWR _31455_/A sky130_fd_sc_hd__mux2_1
X_19176_ _19101_/X _19174_/X _19175_/X _19106_/X VGND VGND VPWR VPWR _19176_/X sky130_fd_sc_hd__a22o_1
X_16388_ _34007_/Q _33943_/Q _33879_/Q _32151_/Q _16314_/X _16315_/X VGND VGND VPWR
+ VPWR _16388_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18127_ _17901_/X _18125_/X _18126_/X _17906_/X VGND VGND VPWR VPWR _18127_/X sky130_fd_sc_hd__a22o_1
XFILLER_185_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30405_ _23253_/X _35441_/Q _30413_/S VGND VGND VPWR VPWR _30406_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34173_ _36157_/CLK _34173_/D VGND VGND VPWR VPWR _34173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31385_ _31385_/A VGND VGND VPWR VPWR _35905_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33124_ _36132_/CLK _33124_/D VGND VGND VPWR VPWR _33124_/Q sky130_fd_sc_hd__dfxtp_1
X_18058_ _17855_/X _18056_/X _18057_/X _17858_/X VGND VGND VPWR VPWR _18058_/X sky130_fd_sc_hd__a22o_1
X_30336_ _23093_/X _35408_/Q _30350_/S VGND VGND VPWR VPWR _30337_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17009_ _16796_/X _17005_/X _17008_/X _16799_/X VGND VGND VPWR VPWR _17009_/X sky130_fd_sc_hd__a22o_1
X_33055_ _36124_/CLK _33055_/D VGND VGND VPWR VPWR _33055_/Q sky130_fd_sc_hd__dfxtp_1
X_30267_ _35376_/Q _29157_/X _30277_/S VGND VGND VPWR VPWR _30268_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20020_ _20020_/A _20020_/B _20020_/C _20020_/D VGND VGND VPWR VPWR _20021_/A sky130_fd_sc_hd__or4_4
X_32006_ _36194_/CLK _32006_/D VGND VGND VPWR VPWR _32006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30198_ _35343_/Q _29055_/X _30214_/S VGND VGND VPWR VPWR _30199_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_859 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21971_ _21795_/X _21969_/X _21970_/X _21800_/X VGND VGND VPWR VPWR _21971_/X sky130_fd_sc_hd__a22o_1
X_33957_ _36134_/CLK _33957_/D VGND VGND VPWR VPWR _33957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_282_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _33083_/CLK sky130_fd_sc_hd__clkbuf_16
X_23710_ _23710_/A VGND VGND VPWR VPWR _32401_/D sky130_fd_sc_hd__clkbuf_1
X_20922_ _32469_/Q _32341_/Q _32021_/Q _35989_/Q _20817_/X _22463_/A VGND VGND VPWR
+ VPWR _20922_/X sky130_fd_sc_hd__mux4_1
XFILLER_26_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32908_ _35919_/CLK _32908_/D VGND VGND VPWR VPWR _32908_/Q sky130_fd_sc_hd__dfxtp_1
X_24690_ _24690_/A VGND VGND VPWR VPWR _32832_/D sky130_fd_sc_hd__clkbuf_1
X_33888_ _34016_/CLK _33888_/D VGND VGND VPWR VPWR _33888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32839_ _34752_/CLK _32839_/D VGND VGND VPWR VPWR _32839_/Q sky130_fd_sc_hd__dfxtp_1
X_20853_ _20849_/X _20852_/X _20640_/X _20642_/X VGND VGND VPWR VPWR _20870_/B sky130_fd_sc_hd__o211a_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35627_ _35818_/CLK _35627_/D VGND VGND VPWR VPWR _35627_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23641_ _23641_/A VGND VGND VPWR VPWR _32370_/D sky130_fd_sc_hd__clkbuf_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23572_ _23572_/A VGND VGND VPWR VPWR _32337_/D sky130_fd_sc_hd__clkbuf_1
X_26360_ _25109_/X _33588_/Q _26362_/S VGND VGND VPWR VPWR _26361_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_922 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20784_ _32465_/Q _32337_/Q _32017_/Q _35985_/Q _20628_/X _22463_/A VGND VGND VPWR
+ VPWR _20784_/X sky130_fd_sc_hd__mux4_1
X_35558_ _35750_/CLK _35558_/D VGND VGND VPWR VPWR _35558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22523_ _22300_/X _22521_/X _22522_/X _22303_/X VGND VGND VPWR VPWR _22523_/X sky130_fd_sc_hd__a22o_1
X_25311_ _25311_/A VGND VGND VPWR VPWR _33095_/D sky130_fd_sc_hd__clkbuf_1
X_26291_ _25007_/X _33555_/Q _26299_/S VGND VGND VPWR VPWR _26292_/A sky130_fd_sc_hd__mux2_1
X_34509_ _35789_/CLK _34509_/D VGND VGND VPWR VPWR _34509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35489_ _35552_/CLK _35489_/D VGND VGND VPWR VPWR _35489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28030_ _26912_/X _34347_/Q _28030_/S VGND VGND VPWR VPWR _28031_/A sky130_fd_sc_hd__mux2_1
X_22454_ _22449_/X _22452_/X _22453_/X VGND VGND VPWR VPWR _22469_/C sky130_fd_sc_hd__o21ba_1
X_25242_ _25242_/A VGND VGND VPWR VPWR _33062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21405_ _35042_/Q _34978_/Q _34914_/Q _34850_/Q _21403_/X _21404_/X VGND VGND VPWR
+ VPWR _21405_/X sky130_fd_sc_hd__mux4_1
X_25173_ _25173_/A VGND VGND VPWR VPWR _33032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22385_ _34814_/Q _34750_/Q _34686_/Q _34622_/Q _22241_/X _22242_/X VGND VGND VPWR
+ VPWR _22385_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_1002 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24124_ _24124_/A VGND VGND VPWR VPWR _32596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21336_ _22556_/A VGND VGND VPWR VPWR _21336_/X sky130_fd_sc_hd__buf_4
XFILLER_191_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29981_ _29981_/A VGND VGND VPWR VPWR _35240_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28932_ _28932_/A VGND VGND VPWR VPWR _34774_/D sky130_fd_sc_hd__clkbuf_1
X_24055_ _24055_/A VGND VGND VPWR VPWR _32564_/D sky130_fd_sc_hd__clkbuf_1
X_21267_ _22446_/A VGND VGND VPWR VPWR _21267_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_151_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23006_ _23006_/A VGND VGND VPWR VPWR _32054_/D sky130_fd_sc_hd__clkbuf_1
X_20218_ _33026_/Q _32962_/Q _32898_/Q _32834_/Q _19995_/X _19996_/X VGND VGND VPWR
+ VPWR _20218_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28863_ _28911_/S VGND VGND VPWR VPWR _28882_/S sky130_fd_sc_hd__buf_4
X_21198_ _21096_/X _21196_/X _21197_/X _21099_/X VGND VGND VPWR VPWR _21198_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27814_ _27814_/A VGND VGND VPWR VPWR _34244_/D sky130_fd_sc_hd__clkbuf_1
X_20149_ _20000_/X _20145_/X _20148_/X _20003_/X VGND VGND VPWR VPWR _20149_/X sky130_fd_sc_hd__a22o_1
XTAP_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28794_ _26844_/X _34709_/Q _28798_/S VGND VGND VPWR VPWR _28795_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27745_ _27745_/A VGND VGND VPWR VPWR _34211_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24957_ _24957_/A VGND VGND VPWR VPWR _32958_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_273_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _36157_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23908_ _22982_/X _32495_/Q _23920_/S VGND VGND VPWR VPWR _23909_/A sky130_fd_sc_hd__mux2_1
XFILLER_246_896 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27676_ _34179_/Q _24410_/X _27688_/S VGND VGND VPWR VPWR _27677_/A sky130_fd_sc_hd__mux2_1
XTAP_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_400 _36210_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24888_ _24888_/A VGND VGND VPWR VPWR _32925_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_411 _36212_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29415_ _23130_/X _34972_/Q _29425_/S VGND VGND VPWR VPWR _29416_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_422 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26627_ _25103_/X _33714_/Q _26633_/S VGND VGND VPWR VPWR _26628_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_433 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23839_ _22875_/X _32462_/Q _23857_/S VGND VGND VPWR VPWR _23840_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_444 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_455 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_466 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29346_ _29346_/A VGND VGND VPWR VPWR _34939_/D sky130_fd_sc_hd__clkbuf_1
X_17360_ _17713_/A VGND VGND VPWR VPWR _17360_/X sky130_fd_sc_hd__buf_4
XFILLER_18_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_477 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26558_ _25001_/X _33681_/Q _26570_/S VGND VGND VPWR VPWR _26559_/A sky130_fd_sc_hd__mux2_1
XANTENNA_488 _31994_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_499 _32008_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16311_ _34261_/Q _34197_/Q _34133_/Q _34069_/Q _16005_/X _16007_/X VGND VGND VPWR
+ VPWR _16311_/X sky130_fd_sc_hd__mux4_1
X_25509_ _25509_/A VGND VGND VPWR VPWR _33186_/D sky130_fd_sc_hd__clkbuf_1
X_17291_ _35312_/Q _35248_/Q _35184_/Q _32304_/Q _17006_/X _17007_/X VGND VGND VPWR
+ VPWR _17291_/X sky130_fd_sc_hd__mux4_1
X_29277_ _29277_/A VGND VGND VPWR VPWR _34906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_1389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26489_ _25100_/X _33649_/Q _26497_/S VGND VGND VPWR VPWR _26490_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19030_ _35040_/Q _34976_/Q _34912_/Q _34848_/Q _18750_/X _18751_/X VGND VGND VPWR
+ VPWR _19030_/X sky130_fd_sc_hd__mux4_1
X_16242_ _16136_/X _16240_/X _16241_/X _16141_/X VGND VGND VPWR VPWR _16242_/X sky130_fd_sc_hd__a22o_1
X_28228_ _27005_/X _34441_/Q _28228_/S VGND VGND VPWR VPWR _28229_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16173_ _16173_/A VGND VGND VPWR VPWR _31952_/D sky130_fd_sc_hd__clkbuf_1
X_28159_ _26903_/X _34408_/Q _28165_/S VGND VGND VPWR VPWR _28160_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput109 _31977_/Q VGND VGND VPWR VPWR D1[27] sky130_fd_sc_hd__buf_2
X_31170_ _31170_/A VGND VGND VPWR VPWR _35803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30121_ _35307_/Q _29141_/X _30121_/S VGND VGND VPWR VPWR _30122_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19932_ _19716_/X _19930_/X _19931_/X _19720_/X VGND VGND VPWR VPWR _19932_/X sky130_fd_sc_hd__a22o_1
XFILLER_123_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30052_ _30052_/A VGND VGND VPWR VPWR _35274_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19863_ _19708_/X _19861_/X _19862_/X _19714_/X VGND VGND VPWR VPWR _19863_/X sky130_fd_sc_hd__a22o_1
XFILLER_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput91 _31960_/Q VGND VGND VPWR VPWR D1[10] sky130_fd_sc_hd__buf_2
XFILLER_96_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18814_ _18593_/X _18812_/X _18813_/X _18596_/X VGND VGND VPWR VPWR _18814_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19794_ _20147_/A VGND VGND VPWR VPWR _19794_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34860_ _35313_/CLK _34860_/D VGND VGND VPWR VPWR _34860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33811_ _35733_/CLK _33811_/D VGND VGND VPWR VPWR _33811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18745_ _35288_/Q _35224_/Q _35160_/Q _32280_/Q _18600_/X _18601_/X VGND VGND VPWR
+ VPWR _18745_/X sky130_fd_sc_hd__mux4_1
XTAP_5380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34791_ _34792_/CLK _34791_/D VGND VGND VPWR VPWR _34791_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_264_CLK clkbuf_6_57__f_CLK/X VGND VGND VPWR VPWR _36097_/CLK sky130_fd_sc_hd__clkbuf_16
X_33742_ _34256_/CLK _33742_/D VGND VGND VPWR VPWR _33742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18676_ _34518_/Q _32406_/Q _34390_/Q _34326_/Q _18466_/X _18467_/X VGND VGND VPWR
+ VPWR _18676_/X sky130_fd_sc_hd__mux4_1
X_30954_ _30954_/A VGND VGND VPWR VPWR _35701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17627_ _33274_/Q _36154_/Q _33146_/Q _33082_/Q _17411_/X _17412_/X VGND VGND VPWR
+ VPWR _17627_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33673_ _34752_/CLK _33673_/D VGND VGND VPWR VPWR _33673_/Q sky130_fd_sc_hd__dfxtp_1
X_30885_ _30885_/A VGND VGND VPWR VPWR _35668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35412_ _35927_/CLK _35412_/D VGND VGND VPWR VPWR _35412_/Q sky130_fd_sc_hd__dfxtp_1
X_32624_ _33262_/CLK _32624_/D VGND VGND VPWR VPWR _32624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17558_ _17911_/A VGND VGND VPWR VPWR _17558_/X sky130_fd_sc_hd__clkbuf_4
X_35343_ _35597_/CLK _35343_/D VGND VGND VPWR VPWR _35343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16509_ _35802_/Q _32177_/Q _35674_/Q _35610_/Q _16254_/X _16255_/X VGND VGND VPWR
+ VPWR _16509_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32555_ _35307_/CLK _32555_/D VGND VGND VPWR VPWR _32555_/Q sky130_fd_sc_hd__dfxtp_1
X_17489_ _17842_/A VGND VGND VPWR VPWR _17489_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_31_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31506_ _23286_/X _35963_/Q _31514_/S VGND VGND VPWR VPWR _31507_/A sky130_fd_sc_hd__mux2_1
X_19228_ _35814_/Q _32190_/Q _35686_/Q _35622_/Q _18907_/X _18908_/X VGND VGND VPWR
+ VPWR _19228_/X sky130_fd_sc_hd__mux4_1
X_35274_ _35340_/CLK _35274_/D VGND VGND VPWR VPWR _35274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32486_ _35303_/CLK _32486_/D VGND VGND VPWR VPWR _32486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34225_ _34227_/CLK _34225_/D VGND VGND VPWR VPWR _34225_/Q sky130_fd_sc_hd__dfxtp_1
X_31437_ _23124_/X _35930_/Q _31451_/S VGND VGND VPWR VPWR _31438_/A sky130_fd_sc_hd__mux2_1
X_19159_ _32996_/Q _32932_/Q _32868_/Q _32804_/Q _18936_/X _18937_/X VGND VGND VPWR
+ VPWR _19159_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22170_ _21947_/X _22168_/X _22169_/X _21950_/X VGND VGND VPWR VPWR _22170_/X sky130_fd_sc_hd__a22o_1
X_34156_ _36074_/CLK _34156_/D VGND VGND VPWR VPWR _34156_/Q sky130_fd_sc_hd__dfxtp_1
X_31368_ _31368_/A VGND VGND VPWR VPWR _35897_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33107_ _36115_/CLK _33107_/D VGND VGND VPWR VPWR _33107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21121_ _34522_/Q _32410_/Q _34394_/Q _34330_/Q _21119_/X _21120_/X VGND VGND VPWR
+ VPWR _21121_/X sky130_fd_sc_hd__mux4_1
X_30319_ _35401_/Q _29234_/X _30319_/S VGND VGND VPWR VPWR _30320_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_1339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34087_ _34087_/CLK _34087_/D VGND VGND VPWR VPWR _34087_/Q sky130_fd_sc_hd__dfxtp_1
X_31299_ _31299_/A VGND VGND VPWR VPWR _35864_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33038_ _36114_/CLK _33038_/D VGND VGND VPWR VPWR _33038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21052_ _35032_/Q _34968_/Q _34904_/Q _34840_/Q _21050_/X _21051_/X VGND VGND VPWR
+ VPWR _21052_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_1227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20003_ _20158_/A VGND VGND VPWR VPWR _20003_/X sky130_fd_sc_hd__buf_4
XFILLER_154_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25860_ _25168_/X _33351_/Q _25864_/S VGND VGND VPWR VPWR _25861_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24811_ _23013_/X _32889_/Q _24823_/S VGND VGND VPWR VPWR _24812_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25791_ _25066_/X _33318_/Q _25801_/S VGND VGND VPWR VPWR _25792_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34989_ _35054_/CLK _34989_/D VGND VGND VPWR VPWR _34989_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_255_CLK clkbuf_6_62__f_CLK/X VGND VGND VPWR VPWR _33922_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27530_ _26974_/X _34111_/Q _27530_/S VGND VGND VPWR VPWR _27531_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24742_ _22910_/X _32856_/Q _24760_/S VGND VGND VPWR VPWR _24743_/A sky130_fd_sc_hd__mux2_1
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21954_ _33202_/Q _32562_/Q _35954_/Q _35890_/Q _21674_/X _21675_/X VGND VGND VPWR
+ VPWR _21954_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20905_ _35028_/Q _34964_/Q _34900_/Q _34836_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _20905_/X sky130_fd_sc_hd__mux4_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27461_ _26872_/X _34078_/Q _27467_/S VGND VGND VPWR VPWR _27462_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24673_ _24673_/A VGND VGND VPWR VPWR _32824_/D sky130_fd_sc_hd__clkbuf_1
X_21885_ _33200_/Q _32560_/Q _35952_/Q _35888_/Q _21674_/X _21675_/X VGND VGND VPWR
+ VPWR _21885_/X sky130_fd_sc_hd__mux4_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29200_ input43/X VGND VGND VPWR VPWR _29200_/X sky130_fd_sc_hd__clkbuf_4
X_26412_ _25186_/X _33613_/Q _26412_/S VGND VGND VPWR VPWR _26413_/A sky130_fd_sc_hd__mux2_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20836_ _20687_/X _20834_/X _20835_/X _20697_/X VGND VGND VPWR VPWR _20836_/X sky130_fd_sc_hd__a22o_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23624_ _23624_/A VGND VGND VPWR VPWR _32362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27392_ _27392_/A VGND VGND VPWR VPWR _34045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_230_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29131_ _29131_/A VGND VGND VPWR VPWR _34855_/D sky130_fd_sc_hd__clkbuf_1
X_26343_ _26412_/S VGND VGND VPWR VPWR _26362_/S sky130_fd_sc_hd__buf_6
X_23555_ _23068_/X _32331_/Q _23559_/S VGND VGND VPWR VPWR _23556_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20767_ _21473_/A VGND VGND VPWR VPWR _20767_/X sky130_fd_sc_hd__buf_6
XFILLER_167_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22506_ _22506_/A VGND VGND VPWR VPWR _22506_/X sky130_fd_sc_hd__buf_4
X_29062_ _34833_/Q _29061_/X _29080_/S VGND VGND VPWR VPWR _29063_/A sky130_fd_sc_hd__mux2_1
X_26274_ _26274_/A VGND VGND VPWR VPWR _33547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23486_ _22966_/X _32298_/Q _23488_/S VGND VGND VPWR VPWR _23487_/A sky130_fd_sc_hd__mux2_1
X_20698_ _20687_/X _20691_/X _20695_/X _20697_/X VGND VGND VPWR VPWR _20698_/X sky130_fd_sc_hd__a22o_1
XFILLER_183_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28013_ _28013_/A VGND VGND VPWR VPWR _34338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22437_ _33280_/Q _36160_/Q _33152_/Q _33088_/Q _22364_/X _22365_/X VGND VGND VPWR
+ VPWR _22437_/X sky130_fd_sc_hd__mux4_1
X_25225_ _25225_/A VGND VGND VPWR VPWR _33054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25156_ input49/X VGND VGND VPWR VPWR _25156_/X sky130_fd_sc_hd__buf_2
X_22368_ _22361_/X _22363_/X _22366_/X _22367_/X VGND VGND VPWR VPWR _22368_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24107_ _24107_/A VGND VGND VPWR VPWR _32589_/D sky130_fd_sc_hd__clkbuf_1
X_21319_ _21241_/X _21317_/X _21318_/X _21244_/X VGND VGND VPWR VPWR _21319_/X sky130_fd_sc_hd__a22o_1
X_29964_ _29964_/A VGND VGND VPWR VPWR _35232_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25087_ _25087_/A VGND VGND VPWR VPWR _33004_/D sky130_fd_sc_hd__clkbuf_1
X_22299_ _22293_/X _22298_/X _22089_/X _22090_/X VGND VGND VPWR VPWR _22320_/B sky130_fd_sc_hd__o211a_1
XFILLER_85_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28915_ _34766_/Q _24244_/X _28933_/S VGND VGND VPWR VPWR _28916_/A sky130_fd_sc_hd__mux2_1
X_24038_ _22972_/X _32556_/Q _24056_/S VGND VGND VPWR VPWR _24039_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29895_ _29922_/S VGND VGND VPWR VPWR _29914_/S sky130_fd_sc_hd__buf_6
XFILLER_77_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_494_CLK clkbuf_leaf_2_CLK/A VGND VGND VPWR VPWR _35040_/CLK sky130_fd_sc_hd__clkbuf_16
X_28846_ _28846_/A VGND VGND VPWR VPWR _34733_/D sky130_fd_sc_hd__clkbuf_1
X_16860_ _16710_/X _16858_/X _16859_/X _16714_/X VGND VGND VPWR VPWR _16860_/X sky130_fd_sc_hd__a22o_1
XFILLER_172_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28777_ _28777_/A VGND VGND VPWR VPWR _34701_/D sky130_fd_sc_hd__clkbuf_1
X_16791_ _35554_/Q _35490_/Q _35426_/Q _35362_/Q _16544_/X _16545_/X VGND VGND VPWR
+ VPWR _16791_/X sky130_fd_sc_hd__mux4_1
X_25989_ _25159_/X _33412_/Q _25999_/S VGND VGND VPWR VPWR _25990_/A sky130_fd_sc_hd__mux2_1
XFILLER_203_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_246_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _33795_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_248_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_1193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18530_ _20295_/A VGND VGND VPWR VPWR _18530_/X sky130_fd_sc_hd__buf_4
XFILLER_20_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27728_ _27728_/A VGND VGND VPWR VPWR _34203_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _18356_/X _18459_/X _18460_/X _18368_/X VGND VGND VPWR VPWR _18461_/X sky130_fd_sc_hd__a22o_1
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27659_ _34171_/Q _24385_/X _27667_/S VGND VGND VPWR VPWR _27660_/A sky130_fd_sc_hd__mux2_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_230 _32136_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_241 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_252 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _17770_/A VGND VGND VPWR VPWR _17412_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_234_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_263 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18392_ _20162_/A VGND VGND VPWR VPWR _18392_/X sky130_fd_sc_hd__buf_4
X_30670_ _30670_/A VGND VGND VPWR VPWR _35566_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_274 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_296 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29329_ _29329_/A VGND VGND VPWR VPWR _34931_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_38__f_CLK clkbuf_5_19_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_38__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_17343_ _17830_/A VGND VGND VPWR VPWR _17343_/X sky130_fd_sc_hd__buf_4
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32340_ _35002_/CLK _32340_/D VGND VGND VPWR VPWR _32340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17274_ _33264_/Q _36144_/Q _33136_/Q _33072_/Q _17058_/X _17059_/X VGND VGND VPWR
+ VPWR _17274_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19013_ _32992_/Q _32928_/Q _32864_/Q _32800_/Q _18936_/X _18937_/X VGND VGND VPWR
+ VPWR _19013_/X sky130_fd_sc_hd__mux4_1
X_16225_ _35538_/Q _35474_/Q _35410_/Q _35346_/Q _16191_/X _16192_/X VGND VGND VPWR
+ VPWR _16225_/X sky130_fd_sc_hd__mux4_1
X_32271_ _34638_/CLK _32271_/D VGND VGND VPWR VPWR _32271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34010_ _34010_/CLK _34010_/D VGND VGND VPWR VPWR _34010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31222_ _31222_/A VGND VGND VPWR VPWR _35828_/D sky130_fd_sc_hd__clkbuf_1
X_16156_ _35792_/Q _32166_/Q _35664_/Q _35600_/Q _16045_/X _16046_/X VGND VGND VPWR
+ VPWR _16156_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31153_ _31153_/A VGND VGND VPWR VPWR _35795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16087_ _17154_/A VGND VGND VPWR VPWR _16087_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_142_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30104_ _30104_/A VGND VGND VPWR VPWR _35298_/D sky130_fd_sc_hd__clkbuf_1
X_19915_ _19911_/X _19914_/X _19814_/X VGND VGND VPWR VPWR _19916_/D sky130_fd_sc_hd__o21ba_1
X_35961_ _36027_/CLK _35961_/D VGND VGND VPWR VPWR _35961_/Q sky130_fd_sc_hd__dfxtp_1
X_31084_ _35763_/Q _29166_/X _31088_/S VGND VGND VPWR VPWR _31085_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_485_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _35935_/CLK sky130_fd_sc_hd__clkbuf_16
X_30035_ _35266_/Q _29213_/X _30049_/S VGND VGND VPWR VPWR _30036_/A sky130_fd_sc_hd__mux2_1
X_34912_ _35040_/CLK _34912_/D VGND VGND VPWR VPWR _34912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19846_ _19846_/A _19846_/B _19846_/C _19846_/D VGND VGND VPWR VPWR _19847_/A sky130_fd_sc_hd__or4_4
XFILLER_190_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_868 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35892_ _35956_/CLK _35892_/D VGND VGND VPWR VPWR _35892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34843_ _35166_/CLK _34843_/D VGND VGND VPWR VPWR _34843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19777_ _20130_/A VGND VGND VPWR VPWR _19777_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_113_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16989_ _17829_/A VGND VGND VPWR VPWR _16989_/X sky130_fd_sc_hd__buf_6
XFILLER_84_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_237_CLK clkbuf_6_61__f_CLK/X VGND VGND VPWR VPWR _35330_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_225_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18728_ _32984_/Q _32920_/Q _32856_/Q _32792_/Q _18583_/X _18584_/X VGND VGND VPWR
+ VPWR _18728_/X sky130_fd_sc_hd__mux4_1
X_34774_ _35669_/CLK _34774_/D VGND VGND VPWR VPWR _34774_/Q sky130_fd_sc_hd__dfxtp_1
X_31986_ _36201_/CLK _31986_/D VGND VGND VPWR VPWR _31986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33725_ _33789_/CLK _33725_/D VGND VGND VPWR VPWR _33725_/Q sky130_fd_sc_hd__dfxtp_1
X_18659_ _32470_/Q _32342_/Q _32022_/Q _35990_/Q _18517_/X _18658_/X VGND VGND VPWR
+ VPWR _18659_/X sky130_fd_sc_hd__mux4_1
X_30937_ _35693_/Q _29148_/X _30953_/S VGND VGND VPWR VPWR _30938_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21670_ _35818_/Q _32195_/Q _35690_/Q _35626_/Q _21560_/X _21561_/X VGND VGND VPWR
+ VPWR _21670_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30868_ _23345_/X _35661_/Q _30868_/S VGND VGND VPWR VPWR _30869_/A sky130_fd_sc_hd__mux2_1
X_33656_ _34296_/CLK _33656_/D VGND VGND VPWR VPWR _33656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20621_ _22503_/A VGND VGND VPWR VPWR _20621_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_71_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32607_ _35801_/CLK _32607_/D VGND VGND VPWR VPWR _32607_/Q sky130_fd_sc_hd__dfxtp_1
X_33587_ _34289_/CLK _33587_/D VGND VGND VPWR VPWR _33587_/Q sky130_fd_sc_hd__dfxtp_1
X_30799_ _30868_/S VGND VGND VPWR VPWR _30818_/S sky130_fd_sc_hd__buf_6
X_23340_ _32231_/Q _23339_/X _23346_/S VGND VGND VPWR VPWR _23341_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20552_ _32781_/Q _32717_/Q _32653_/Q _36109_/Q _20278_/X _19173_/A VGND VGND VPWR
+ VPWR _20552_/X sky130_fd_sc_hd__mux4_1
X_35326_ _35326_/CLK _35326_/D VGND VGND VPWR VPWR _35326_/Q sky130_fd_sc_hd__dfxtp_1
X_32538_ _35864_/CLK _32538_/D VGND VGND VPWR VPWR _32538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23271_ _23346_/S VGND VGND VPWR VPWR _23301_/S sky130_fd_sc_hd__buf_6
X_20483_ _20483_/A _20483_/B _20483_/C _20483_/D VGND VGND VPWR VPWR _20484_/A sky130_fd_sc_hd__or4_1
XFILLER_192_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32469_ _32983_/CLK _32469_/D VGND VGND VPWR VPWR _32469_/Q sky130_fd_sc_hd__dfxtp_1
X_35257_ _35257_/CLK _35257_/D VGND VGND VPWR VPWR _35257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25010_ input61/X VGND VGND VPWR VPWR _25010_/X sky130_fd_sc_hd__clkbuf_8
X_22222_ _34042_/Q _33978_/Q _33914_/Q _32250_/Q _21973_/X _21974_/X VGND VGND VPWR
+ VPWR _22222_/X sky130_fd_sc_hd__mux4_1
X_34208_ _34777_/CLK _34208_/D VGND VGND VPWR VPWR _34208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35188_ _35315_/CLK _35188_/D VGND VGND VPWR VPWR _35188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1084 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22153_ _22506_/A VGND VGND VPWR VPWR _22153_/X sky130_fd_sc_hd__clkbuf_4
X_34139_ _34267_/CLK _34139_/D VGND VGND VPWR VPWR _34139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21104_ _20949_/X _21102_/X _21103_/X _20955_/X VGND VGND VPWR VPWR _21104_/X sky130_fd_sc_hd__a22o_1
XTAP_6817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26961_ _26961_/A VGND VGND VPWR VPWR _33850_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22084_ _33270_/Q _36150_/Q _33142_/Q _33078_/Q _22011_/X _22012_/X VGND VGND VPWR
+ VPWR _22084_/X sky130_fd_sc_hd__mux4_1
XTAP_6839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_476_CLK clkbuf_6_8__f_CLK/X VGND VGND VPWR VPWR _35299_/CLK sky130_fd_sc_hd__clkbuf_16
X_28700_ _28700_/A VGND VGND VPWR VPWR _34664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21035_ _22595_/A VGND VGND VPWR VPWR _21035_/X sky130_fd_sc_hd__clkbuf_4
X_25912_ _25912_/A VGND VGND VPWR VPWR _33375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29680_ _29680_/A VGND VGND VPWR VPWR _35097_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26892_ _26891_/X _33828_/Q _26913_/S VGND VGND VPWR VPWR _26893_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28631_ _27002_/X _34632_/Q _28633_/S VGND VGND VPWR VPWR _28632_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_1300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25843_ _25143_/X _33343_/Q _25843_/S VGND VGND VPWR VPWR _25844_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_228_CLK clkbuf_6_54__f_CLK/X VGND VGND VPWR VPWR _32518_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_216_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28562_ _26900_/X _34599_/Q _28570_/S VGND VGND VPWR VPWR _28563_/A sky130_fd_sc_hd__mux2_1
X_25774_ _25041_/X _33310_/Q _25780_/S VGND VGND VPWR VPWR _25775_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22986_ _22985_/X _32048_/Q _23001_/S VGND VGND VPWR VPWR _22987_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27513_ _27513_/A VGND VGND VPWR VPWR _34102_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_215_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24725_ _22886_/X _32848_/Q _24739_/S VGND VGND VPWR VPWR _24726_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28493_ _28493_/A VGND VGND VPWR VPWR _34566_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21937_ _21933_/X _21936_/X _21728_/X VGND VGND VPWR VPWR _21967_/A sky130_fd_sc_hd__o21ba_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27444_ _26847_/X _34070_/Q _27446_/S VGND VGND VPWR VPWR _27445_/A sky130_fd_sc_hd__mux2_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24656_ _24656_/A VGND VGND VPWR VPWR _32816_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21868_ _33520_/Q _33456_/Q _33392_/Q _33328_/Q _21723_/X _21724_/X VGND VGND VPWR
+ VPWR _21868_/X sky130_fd_sc_hd__mux4_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23607_ _32354_/Q _23148_/X _23625_/S VGND VGND VPWR VPWR _23608_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20819_ _32978_/Q _32914_/Q _32850_/Q _32786_/Q _20633_/X _20635_/X VGND VGND VPWR
+ VPWR _20819_/X sky130_fd_sc_hd__mux4_1
X_27375_ _27375_/A VGND VGND VPWR VPWR _34037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24587_ _24587_/A VGND VGND VPWR VPWR _32783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21799_ _34286_/Q _34222_/Q _34158_/Q _34094_/Q _21689_/X _21690_/X VGND VGND VPWR
+ VPWR _21799_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_400_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _35946_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29114_ _29247_/S VGND VGND VPWR VPWR _29142_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_129_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26326_ _26326_/A VGND VGND VPWR VPWR _33571_/D sky130_fd_sc_hd__clkbuf_1
X_23538_ _23538_/A VGND VGND VPWR VPWR _32322_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29045_ _29045_/A VGND VGND VPWR VPWR _34828_/D sky130_fd_sc_hd__clkbuf_1
X_26257_ _25156_/X _33539_/Q _26269_/S VGND VGND VPWR VPWR _26258_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23469_ _23559_/S VGND VGND VPWR VPWR _23488_/S sky130_fd_sc_hd__buf_4
X_16010_ input69/X input70/X VGND VGND VPWR VPWR _17834_/A sky130_fd_sc_hd__or2b_4
XFILLER_183_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25208_ _25208_/A VGND VGND VPWR VPWR _33046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26188_ _25053_/X _33506_/Q _26206_/S VGND VGND VPWR VPWR _26189_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25139_ _25139_/A VGND VGND VPWR VPWR _33021_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17961_ _17955_/X _17960_/X _17853_/X VGND VGND VPWR VPWR _17969_/C sky130_fd_sc_hd__o21ba_1
XFILLER_69_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29947_ _35224_/Q _29082_/X _29965_/S VGND VGND VPWR VPWR _29948_/A sky130_fd_sc_hd__mux2_1
X_16912_ _33766_/Q _33702_/Q _33638_/Q _33574_/Q _16843_/X _16844_/X VGND VGND VPWR
+ VPWR _16912_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_467_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _35749_/CLK sky130_fd_sc_hd__clkbuf_16
X_19700_ _19700_/A VGND VGND VPWR VPWR _32115_/D sky130_fd_sc_hd__buf_2
XFILLER_2_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17892_ _34817_/Q _34753_/Q _34689_/Q _34625_/Q _17641_/X _17642_/X VGND VGND VPWR
+ VPWR _17892_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29878_ _29878_/A VGND VGND VPWR VPWR _35191_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19631_ _33778_/Q _33714_/Q _33650_/Q _33586_/Q _19496_/X _19497_/X VGND VGND VPWR
+ VPWR _19631_/X sky130_fd_sc_hd__mux4_1
X_16843_ _17902_/A VGND VGND VPWR VPWR _16843_/X sky130_fd_sc_hd__buf_4
XFILLER_120_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28829_ _28829_/A VGND VGND VPWR VPWR _34725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_219_CLK clkbuf_6_55__f_CLK/X VGND VGND VPWR VPWR _35779_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_226_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31840_ _23121_/X _36121_/Q _31856_/S VGND VGND VPWR VPWR _31841_/A sky130_fd_sc_hd__mux2_1
X_19562_ _19558_/X _19561_/X _19461_/X VGND VGND VPWR VPWR _19563_/D sky130_fd_sc_hd__o21ba_1
X_16774_ _16496_/X _16772_/X _16773_/X _16499_/X VGND VGND VPWR VPWR _16774_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_1294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18513_ _20278_/A VGND VGND VPWR VPWR _18513_/X sky130_fd_sc_hd__buf_6
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31771_ _31771_/A VGND VGND VPWR VPWR _36088_/D sky130_fd_sc_hd__clkbuf_1
X_19493_ _19493_/A _19493_/B _19493_/C _19493_/D VGND VGND VPWR VPWR _19494_/A sky130_fd_sc_hd__or4_1
XFILLER_34_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18444_ _33488_/Q _33424_/Q _33360_/Q _33296_/Q _18298_/X _18299_/X VGND VGND VPWR
+ VPWR _18444_/X sky130_fd_sc_hd__mux4_1
X_30722_ _30722_/A VGND VGND VPWR VPWR _35591_/D sky130_fd_sc_hd__clkbuf_1
X_33510_ _35991_/CLK _33510_/D VGND VGND VPWR VPWR _33510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34490_ _35771_/CLK _34490_/D VGND VGND VPWR VPWR _34490_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33441_ _34145_/CLK _33441_/D VGND VGND VPWR VPWR _33441_/Q sky130_fd_sc_hd__dfxtp_1
X_18375_ _20231_/A VGND VGND VPWR VPWR _18375_/X sky130_fd_sc_hd__buf_6
X_30653_ _30653_/A VGND VGND VPWR VPWR _35558_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17326_ _35057_/Q _34993_/Q _34929_/Q _34865_/Q _17156_/X _17157_/X VGND VGND VPWR
+ VPWR _17326_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36160_ _36160_/CLK _36160_/D VGND VGND VPWR VPWR _36160_/Q sky130_fd_sc_hd__dfxtp_1
X_33372_ _34074_/CLK _33372_/D VGND VGND VPWR VPWR _33372_/Q sky130_fd_sc_hd__dfxtp_1
X_30584_ _23322_/X _35526_/Q _30590_/S VGND VGND VPWR VPWR _30585_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32323_ _35330_/CLK _32323_/D VGND VGND VPWR VPWR _32323_/Q sky130_fd_sc_hd__dfxtp_1
X_35111_ _35750_/CLK _35111_/D VGND VGND VPWR VPWR _35111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36091_ _36156_/CLK _36091_/D VGND VGND VPWR VPWR _36091_/Q sky130_fd_sc_hd__dfxtp_1
X_17257_ _35311_/Q _35247_/Q _35183_/Q _32303_/Q _17006_/X _17007_/X VGND VGND VPWR
+ VPWR _17257_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16208_ _16136_/X _16206_/X _16207_/X _16141_/X VGND VGND VPWR VPWR _16208_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35042_ _35042_/CLK _35042_/D VGND VGND VPWR VPWR _35042_/Q sky130_fd_sc_hd__dfxtp_1
X_32254_ _34046_/CLK _32254_/D VGND VGND VPWR VPWR _32254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17188_ _17149_/X _17186_/X _17187_/X _17152_/X VGND VGND VPWR VPWR _17188_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31205_ _35820_/Q input24/X _31223_/S VGND VGND VPWR VPWR _31206_/A sky130_fd_sc_hd__mux2_1
X_16139_ _33744_/Q _33680_/Q _33616_/Q _33552_/Q _16137_/X _16138_/X VGND VGND VPWR
+ VPWR _16139_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_1434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32185_ _35807_/CLK _32185_/D VGND VGND VPWR VPWR _32185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31136_ _35788_/Q _29243_/X _31138_/S VGND VGND VPWR VPWR _31137_/A sky130_fd_sc_hd__mux2_1
XFILLER_216_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_458_CLK clkbuf_6_10__f_CLK/X VGND VGND VPWR VPWR _34987_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_151_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31067_ _35755_/Q _29141_/X _31067_/S VGND VGND VPWR VPWR _31068_/A sky130_fd_sc_hd__mux2_1
X_35944_ _35944_/CLK _35944_/D VGND VGND VPWR VPWR _35944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30018_ _35258_/Q _29188_/X _30028_/S VGND VGND VPWR VPWR _30019_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19829_ _33015_/Q _32951_/Q _32887_/Q _32823_/Q _19642_/X _19643_/X VGND VGND VPWR
+ VPWR _19829_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35875_ _35940_/CLK _35875_/D VGND VGND VPWR VPWR _35875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34826_ _35338_/CLK _34826_/D VGND VGND VPWR VPWR _34826_/Q sky130_fd_sc_hd__dfxtp_1
X_22840_ _35084_/Q _35020_/Q _34956_/Q _34892_/Q _20679_/X _20681_/X VGND VGND VPWR
+ VPWR _22840_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34757_ _35332_/CLK _34757_/D VGND VGND VPWR VPWR _34757_/Q sky130_fd_sc_hd__dfxtp_1
X_22771_ _20577_/X _22769_/X _22770_/X _20587_/X VGND VGND VPWR VPWR _22771_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31969_ _34970_/CLK _31969_/D VGND VGND VPWR VPWR _31969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24510_ _24510_/A VGND VGND VPWR VPWR _32748_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33708_ _36074_/CLK _33708_/D VGND VGND VPWR VPWR _33708_/Q sky130_fd_sc_hd__dfxtp_1
X_21722_ _21442_/X _21720_/X _21721_/X _21447_/X VGND VGND VPWR VPWR _21722_/X sky130_fd_sc_hd__a22o_1
XFILLER_225_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25490_ _25490_/A VGND VGND VPWR VPWR _33177_/D sky130_fd_sc_hd__clkbuf_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34688_ _35328_/CLK _34688_/D VGND VGND VPWR VPWR _34688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24441_ _32717_/Q _24440_/X _24441_/S VGND VGND VPWR VPWR _24442_/A sky130_fd_sc_hd__mux2_1
X_21653_ _21449_/X _21651_/X _21652_/X _21452_/X VGND VGND VPWR VPWR _21653_/X sky130_fd_sc_hd__a22o_1
X_33639_ _34278_/CLK _33639_/D VGND VGND VPWR VPWR _33639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_21__f_CLK clkbuf_5_10_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_21__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_27160_ _26826_/X _33935_/Q _27176_/S VGND VGND VPWR VPWR _27161_/A sky130_fd_sc_hd__mux2_1
X_20604_ _20657_/A VGND VGND VPWR VPWR _22556_/A sky130_fd_sc_hd__buf_12
X_21584_ _21580_/X _21583_/X _21375_/X VGND VGND VPWR VPWR _21614_/A sky130_fd_sc_hd__o21ba_1
X_24372_ _24372_/A VGND VGND VPWR VPWR _32694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26111_ _25140_/X _33470_/Q _26113_/S VGND VGND VPWR VPWR _26112_/A sky130_fd_sc_hd__mux2_1
X_23323_ _32225_/Q _23322_/X _23334_/S VGND VGND VPWR VPWR _23324_/A sky130_fd_sc_hd__mux2_1
X_20535_ _20531_/X _20534_/X _20153_/A VGND VGND VPWR VPWR _20543_/C sky130_fd_sc_hd__o21ba_1
X_35309_ _35500_/CLK _35309_/D VGND VGND VPWR VPWR _35309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27091_ _27091_/A VGND VGND VPWR VPWR _33902_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26042_ _25038_/X _33437_/Q _26050_/S VGND VGND VPWR VPWR _26043_/A sky130_fd_sc_hd__mux2_1
X_20466_ _33034_/Q _32970_/Q _32906_/Q _32842_/Q _18280_/X _18283_/X VGND VGND VPWR
+ VPWR _20466_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23254_ _32202_/Q _23253_/X _23268_/S VGND VGND VPWR VPWR _23255_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22205_ _35577_/Q _35513_/Q _35449_/Q _35385_/Q _22203_/X _22204_/X VGND VGND VPWR
+ VPWR _22205_/X sky130_fd_sc_hd__mux4_2
XFILLER_84_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23185_ _32175_/Q _23117_/X _23206_/S VGND VGND VPWR VPWR _23186_/A sky130_fd_sc_hd__mux2_1
X_20397_ _20201_/X _20395_/X _20396_/X _20206_/X VGND VGND VPWR VPWR _20397_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29801_ _35155_/Q _29067_/X _29809_/S VGND VGND VPWR VPWR _29802_/A sky130_fd_sc_hd__mux2_1
X_22136_ _33207_/Q _32567_/Q _35959_/Q _35895_/Q _22027_/X _22028_/X VGND VGND VPWR
+ VPWR _22136_/X sky130_fd_sc_hd__mux4_1
XTAP_6614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27993_ _26857_/X _34329_/Q _28009_/S VGND VGND VPWR VPWR _27994_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput270 _32135_/Q VGND VGND VPWR VPWR D3[57] sky130_fd_sc_hd__buf_2
XFILLER_245_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput281 _32087_/Q VGND VGND VPWR VPWR D3[9] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_449_CLK clkbuf_6_9__f_CLK/X VGND VGND VPWR VPWR _36003_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29732_ _29732_/A VGND VGND VPWR VPWR _35122_/D sky130_fd_sc_hd__clkbuf_1
X_22067_ _34549_/Q _32437_/Q _34421_/Q _34357_/Q _21825_/X _21826_/X VGND VGND VPWR
+ VPWR _22067_/X sky130_fd_sc_hd__mux4_1
X_26944_ _26943_/X _33845_/Q _26944_/S VGND VGND VPWR VPWR _26945_/A sky130_fd_sc_hd__mux2_1
XTAP_6669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21018_ _22396_/A VGND VGND VPWR VPWR _21018_/X sky130_fd_sc_hd__buf_4
XFILLER_236_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29663_ _29663_/A VGND VGND VPWR VPWR _35089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26875_ input9/X VGND VGND VPWR VPWR _26875_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28614_ _28641_/S VGND VGND VPWR VPWR _28633_/S sky130_fd_sc_hd__buf_4
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25826_ _25826_/A VGND VGND VPWR VPWR _33334_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29594_ _35057_/Q _29160_/X _29602_/S VGND VGND VPWR VPWR _29595_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28545_ _26875_/X _34591_/Q _28549_/S VGND VGND VPWR VPWR _28546_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25757_ _25016_/X _33302_/Q _25759_/S VGND VGND VPWR VPWR _25758_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22969_ input22/X VGND VGND VPWR VPWR _22969_/X sky130_fd_sc_hd__buf_2
XFILLER_245_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24708_ _24708_/A VGND VGND VPWR VPWR _32841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28476_ _28476_/A VGND VGND VPWR VPWR _34558_/D sky130_fd_sc_hd__clkbuf_1
X_16490_ _17902_/A VGND VGND VPWR VPWR _16490_/X sky130_fd_sc_hd__clkbuf_8
X_25688_ _33270_/Q _24369_/X _25706_/S VGND VGND VPWR VPWR _25689_/A sky130_fd_sc_hd__mux2_1
XFILLER_188_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27427_ _27559_/S VGND VGND VPWR VPWR _27446_/S sky130_fd_sc_hd__buf_4
XFILLER_231_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24639_ _24639_/A VGND VGND VPWR VPWR _32808_/D sky130_fd_sc_hd__clkbuf_1
X_18160_ _17908_/X _18158_/X _18159_/X _17911_/X VGND VGND VPWR VPWR _18160_/X sky130_fd_sc_hd__a22o_1
XFILLER_141_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27358_ _34029_/Q _24342_/X _27374_/S VGND VGND VPWR VPWR _27359_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17111_ _34795_/Q _34731_/Q _34667_/Q _34603_/Q _16935_/X _16936_/X VGND VGND VPWR
+ VPWR _17111_/X sky130_fd_sc_hd__mux4_1
X_26309_ _26309_/A VGND VGND VPWR VPWR _33563_/D sky130_fd_sc_hd__clkbuf_1
X_18091_ _17860_/X _18089_/X _18090_/X _17865_/X VGND VGND VPWR VPWR _18091_/X sky130_fd_sc_hd__a22o_1
XFILLER_141_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27289_ _27017_/X _33997_/Q _27289_/S VGND VGND VPWR VPWR _27290_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29028_ _34820_/Q _24413_/X _29038_/S VGND VGND VPWR VPWR _29029_/A sky130_fd_sc_hd__mux2_1
X_17042_ _34537_/Q _32425_/Q _34409_/Q _34345_/Q _16872_/X _16873_/X VGND VGND VPWR
+ VPWR _17042_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18993_ _18993_/A _18993_/B _18993_/C _18993_/D VGND VGND VPWR VPWR _18994_/A sky130_fd_sc_hd__or4_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17944_ _17908_/X _17942_/X _17943_/X _17911_/X VGND VGND VPWR VPWR _17944_/X sky130_fd_sc_hd__a22o_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33990_ _34243_/CLK _33990_/D VGND VGND VPWR VPWR _33990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17875_ _34049_/Q _33985_/Q _33921_/Q _32257_/Q _17726_/X _17727_/X VGND VGND VPWR
+ VPWR _17875_/X sky130_fd_sc_hd__mux4_1
X_32941_ _36015_/CLK _32941_/D VGND VGND VPWR VPWR _32941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19614_ _20096_/A VGND VGND VPWR VPWR _19614_/X sky130_fd_sc_hd__buf_4
XFILLER_241_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35660_ _35853_/CLK _35660_/D VGND VGND VPWR VPWR _35660_/Q sky130_fd_sc_hd__dfxtp_1
X_16826_ _35811_/Q _32187_/Q _35683_/Q _35619_/Q _16607_/X _16608_/X VGND VGND VPWR
+ VPWR _16826_/X sky130_fd_sc_hd__mux4_1
X_32872_ _36009_/CLK _32872_/D VGND VGND VPWR VPWR _32872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34611_ _35242_/CLK _34611_/D VGND VGND VPWR VPWR _34611_/Q sky130_fd_sc_hd__dfxtp_1
X_31823_ _23096_/X _36113_/Q _31835_/S VGND VGND VPWR VPWR _31824_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16757_ _16753_/X _16756_/X _16441_/X VGND VGND VPWR VPWR _16765_/C sky130_fd_sc_hd__o21ba_1
X_19545_ _19363_/X _19543_/X _19544_/X _19367_/X VGND VGND VPWR VPWR _19545_/X sky130_fd_sc_hd__a22o_1
X_35591_ _35845_/CLK _35591_/D VGND VGND VPWR VPWR _35591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31754_ _31754_/A VGND VGND VPWR VPWR _36080_/D sky130_fd_sc_hd__clkbuf_1
X_34542_ _35052_/CLK _34542_/D VGND VGND VPWR VPWR _34542_/Q sky130_fd_sc_hd__dfxtp_1
X_19476_ _33005_/Q _32941_/Q _32877_/Q _32813_/Q _19289_/X _19290_/X VGND VGND VPWR
+ VPWR _19476_/X sky130_fd_sc_hd__mux4_1
X_16688_ _16443_/X _16686_/X _16687_/X _16446_/X VGND VGND VPWR VPWR _16688_/X sky130_fd_sc_hd__a22o_1
X_30705_ _30705_/A VGND VGND VPWR VPWR _35583_/D sky130_fd_sc_hd__clkbuf_1
X_18427_ _34767_/Q _34703_/Q _34639_/Q _34575_/Q _18375_/X _18376_/X VGND VGND VPWR
+ VPWR _18427_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31685_ _31685_/A VGND VGND VPWR VPWR _36047_/D sky130_fd_sc_hd__clkbuf_1
X_34473_ _34859_/CLK _34473_/D VGND VGND VPWR VPWR _34473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36212_ _36216_/CLK _36212_/D VGND VGND VPWR VPWR _36212_/Q sky130_fd_sc_hd__dfxtp_1
X_33424_ _33940_/CLK _33424_/D VGND VGND VPWR VPWR _33424_/Q sky130_fd_sc_hd__dfxtp_1
X_18358_ _20146_/A VGND VGND VPWR VPWR _18358_/X sky130_fd_sc_hd__buf_8
XFILLER_221_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30636_ _30636_/A VGND VGND VPWR VPWR _35550_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_19_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_19_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_17309_ _32497_/Q _32369_/Q _32049_/Q _36017_/Q _17276_/X _17064_/X VGND VGND VPWR
+ VPWR _17309_/X sky130_fd_sc_hd__mux4_1
X_33355_ _33548_/CLK _33355_/D VGND VGND VPWR VPWR _33355_/Q sky130_fd_sc_hd__dfxtp_1
X_36143_ _36146_/CLK _36143_/D VGND VGND VPWR VPWR _36143_/Q sky130_fd_sc_hd__dfxtp_1
X_18289_ _20095_/A VGND VGND VPWR VPWR _18289_/X sky130_fd_sc_hd__clkbuf_8
X_30567_ _23297_/X _35518_/Q _30569_/S VGND VGND VPWR VPWR _30568_/A sky130_fd_sc_hd__mux2_1
X_20320_ _35781_/Q _35141_/Q _34501_/Q _33861_/Q _20146_/X _20147_/X VGND VGND VPWR
+ VPWR _20320_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32306_ _35700_/CLK _32306_/D VGND VGND VPWR VPWR _32306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33286_ _36166_/CLK _33286_/D VGND VGND VPWR VPWR _33286_/Q sky130_fd_sc_hd__dfxtp_1
X_36074_ _36074_/CLK _36074_/D VGND VGND VPWR VPWR _36074_/Q sky130_fd_sc_hd__dfxtp_1
X_30498_ _23133_/X _35485_/Q _30506_/S VGND VGND VPWR VPWR _30499_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20251_ _20069_/X _20249_/X _20250_/X _20073_/X VGND VGND VPWR VPWR _20251_/X sky130_fd_sc_hd__a22o_1
X_35025_ _35281_/CLK _35025_/D VGND VGND VPWR VPWR _35025_/Q sky130_fd_sc_hd__dfxtp_1
X_32237_ _35955_/CLK _32237_/D VGND VGND VPWR VPWR _32237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32168_ _35921_/CLK _32168_/D VGND VGND VPWR VPWR _32168_/Q sky130_fd_sc_hd__dfxtp_1
X_20182_ _33025_/Q _32961_/Q _32897_/Q _32833_/Q _19995_/X _19996_/X VGND VGND VPWR
+ VPWR _20182_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31119_ _31119_/A VGND VGND VPWR VPWR _35779_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24990_ _25462_/A _27561_/B VGND VGND VPWR VPWR _28373_/B sky130_fd_sc_hd__nor2_8
XFILLER_131_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32099_ _35808_/CLK _32099_/D VGND VGND VPWR VPWR _32099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23941_ _23031_/X _32511_/Q _23941_/S VGND VGND VPWR VPWR _23942_/A sky130_fd_sc_hd__mux2_1
XTAP_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35927_ _35927_/CLK _35927_/D VGND VGND VPWR VPWR _35927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26660_ _26660_/A VGND VGND VPWR VPWR _33729_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35858_ _35921_/CLK _35858_/D VGND VGND VPWR VPWR _35858_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23872_ _22929_/X _32478_/Q _23878_/S VGND VGND VPWR VPWR _23873_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25611_ _25611_/A VGND VGND VPWR VPWR _33233_/D sky130_fd_sc_hd__clkbuf_1
X_22823_ _33292_/Q _36172_/Q _33164_/Q _33100_/Q _20628_/X _21757_/A VGND VGND VPWR
+ VPWR _22823_/X sky130_fd_sc_hd__mux4_1
XANTENNA_807 _22901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_34809_ _34809_/CLK _34809_/D VGND VGND VPWR VPWR _34809_/Q sky130_fd_sc_hd__dfxtp_1
X_26591_ _25050_/X _33697_/Q _26591_/S VGND VGND VPWR VPWR _26592_/A sky130_fd_sc_hd__mux2_1
XANTENNA_818 _22988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35789_ _35789_/CLK _35789_/D VGND VGND VPWR VPWR _35789_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_829 _23127_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28330_ _34489_/Q _24379_/X _28342_/S VGND VGND VPWR VPWR _28331_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25542_ _25542_/A VGND VGND VPWR VPWR _33202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22754_ _22754_/A VGND VGND VPWR VPWR _36233_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21705_ _35755_/Q _35115_/Q _34475_/Q _33835_/Q _21387_/X _21388_/X VGND VGND VPWR
+ VPWR _21705_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28261_ _34456_/Q _24276_/X _28279_/S VGND VGND VPWR VPWR _28262_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25473_ _25473_/A VGND VGND VPWR VPWR _33169_/D sky130_fd_sc_hd__clkbuf_1
X_22685_ _22681_/X _22684_/X _22453_/X VGND VGND VPWR VPWR _22693_/C sky130_fd_sc_hd__o21ba_1
XFILLER_90_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27212_ _26903_/X _33960_/Q _27218_/S VGND VGND VPWR VPWR _27213_/A sky130_fd_sc_hd__mux2_1
X_24424_ _24424_/A VGND VGND VPWR VPWR _32711_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28192_ _28192_/A VGND VGND VPWR VPWR _34423_/D sky130_fd_sc_hd__clkbuf_1
X_21636_ _33193_/Q _32553_/Q _35945_/Q _35881_/Q _21321_/X _21322_/X VGND VGND VPWR
+ VPWR _21636_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27143_ _27143_/A VGND VGND VPWR VPWR _33927_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24355_ _32689_/Q _24354_/X _24367_/S VGND VGND VPWR VPWR _24356_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21567_ _21246_/X _21565_/X _21566_/X _21249_/X VGND VGND VPWR VPWR _21567_/X sky130_fd_sc_hd__a22o_1
X_23306_ _23306_/A VGND VGND VPWR VPWR _32219_/D sky130_fd_sc_hd__clkbuf_1
X_20518_ _33548_/Q _33484_/Q _33420_/Q _33356_/Q _18333_/X _18335_/X VGND VGND VPWR
+ VPWR _20518_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27074_ _27074_/A VGND VGND VPWR VPWR _33894_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21498_ _22557_/A VGND VGND VPWR VPWR _21498_/X sky130_fd_sc_hd__buf_4
X_24286_ input5/X VGND VGND VPWR VPWR _24286_/X sky130_fd_sc_hd__buf_4
XFILLER_181_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26025_ _25013_/X _33429_/Q _26029_/S VGND VGND VPWR VPWR _26026_/A sky130_fd_sc_hd__mux2_1
X_20449_ _34569_/Q _32457_/Q _34441_/Q _34377_/Q _20231_/X _20232_/X VGND VGND VPWR
+ VPWR _20449_/X sky130_fd_sc_hd__mux4_1
X_23237_ input24/X VGND VGND VPWR VPWR _23237_/X sky130_fd_sc_hd__buf_4
XTAP_7101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23168_ _23168_/A VGND VGND VPWR VPWR _32167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1206 _23136_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1217 _24261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1228 _24410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22119_ _34295_/Q _34231_/Q _34167_/Q _34103_/Q _22042_/X _22043_/X VGND VGND VPWR
+ VPWR _22119_/X sky130_fd_sc_hd__mux4_1
X_15990_ _16059_/A VGND VGND VPWR VPWR _17796_/A sky130_fd_sc_hd__buf_12
XTAP_5710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1239 _25735_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27976_ _26832_/X _34321_/Q _27988_/S VGND VGND VPWR VPWR _27977_/A sky130_fd_sc_hd__mux2_1
X_23099_ input45/X VGND VGND VPWR VPWR _23099_/X sky130_fd_sc_hd__buf_4
XFILLER_95_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26927_ _26927_/A VGND VGND VPWR VPWR _33839_/D sky130_fd_sc_hd__clkbuf_1
X_29715_ _29715_/A VGND VGND VPWR VPWR _35114_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17660_ _33275_/Q _36155_/Q _33147_/Q _33083_/Q _17411_/X _17412_/X VGND VGND VPWR
+ VPWR _17660_/X sky130_fd_sc_hd__mux4_1
X_29646_ _35082_/Q _29237_/X _29652_/S VGND VGND VPWR VPWR _29647_/A sky130_fd_sc_hd__mux2_1
XTAP_5798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26858_ _26857_/X _33817_/Q _26882_/S VGND VGND VPWR VPWR _26859_/A sky130_fd_sc_hd__mux2_1
X_16611_ _16288_/X _16609_/X _16610_/X _16291_/X VGND VGND VPWR VPWR _16611_/X sky130_fd_sc_hd__a22o_1
X_25809_ _25809_/A VGND VGND VPWR VPWR _33326_/D sky130_fd_sc_hd__clkbuf_1
X_17591_ _17555_/X _17589_/X _17590_/X _17558_/X VGND VGND VPWR VPWR _17591_/X sky130_fd_sc_hd__a22o_1
X_29577_ _35049_/Q _29135_/X _29581_/S VGND VGND VPWR VPWR _29578_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26789_ _26789_/A VGND VGND VPWR VPWR _33790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28528_ _26850_/X _34583_/Q _28528_/S VGND VGND VPWR VPWR _28529_/A sky130_fd_sc_hd__mux2_1
X_16542_ _35739_/Q _35099_/Q _34459_/Q _33819_/Q _16434_/X _16435_/X VGND VGND VPWR
+ VPWR _16542_/X sky130_fd_sc_hd__mux4_1
X_19330_ _19010_/X _19328_/X _19329_/X _19014_/X VGND VGND VPWR VPWR _19330_/X sky130_fd_sc_hd__a22o_1
XFILLER_204_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19261_ _20096_/A VGND VGND VPWR VPWR _19261_/X sky130_fd_sc_hd__buf_4
XFILLER_206_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28459_ _26946_/X _34550_/Q _28477_/S VGND VGND VPWR VPWR _28460_/A sky130_fd_sc_hd__mux2_1
X_16473_ _35801_/Q _32176_/Q _35673_/Q _35609_/Q _16254_/X _16255_/X VGND VGND VPWR
+ VPWR _16473_/X sky130_fd_sc_hd__mux4_1
X_18212_ _18208_/X _18211_/X _17867_/A VGND VGND VPWR VPWR _18213_/D sky130_fd_sc_hd__o21ba_1
XFILLER_223_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31470_ _23231_/X _35946_/Q _31472_/S VGND VGND VPWR VPWR _31471_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19192_ _19010_/X _19190_/X _19191_/X _19014_/X VGND VGND VPWR VPWR _19192_/X sky130_fd_sc_hd__a22o_1
XFILLER_223_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18143_ _33225_/Q _32585_/Q _35977_/Q _35913_/Q _16075_/X _16076_/X VGND VGND VPWR
+ VPWR _18143_/X sky130_fd_sc_hd__mux4_1
X_30421_ _30421_/A VGND VGND VPWR VPWR _35448_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33140_ _36149_/CLK _33140_/D VGND VGND VPWR VPWR _33140_/Q sky130_fd_sc_hd__dfxtp_1
X_18074_ _17761_/X _18072_/X _18073_/X _17767_/X VGND VGND VPWR VPWR _18074_/X sky130_fd_sc_hd__a22o_1
X_30352_ _30463_/S VGND VGND VPWR VPWR _30371_/S sky130_fd_sc_hd__buf_4
XFILLER_145_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17025_ _32745_/Q _32681_/Q _32617_/Q _36073_/Q _16919_/X _16703_/X VGND VGND VPWR
+ VPWR _17025_/X sky130_fd_sc_hd__mux4_1
XFILLER_171_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33071_ _36081_/CLK _33071_/D VGND VGND VPWR VPWR _33071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30283_ _30283_/A VGND VGND VPWR VPWR _35383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32022_ _33507_/CLK _32022_/D VGND VGND VPWR VPWR _32022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18976_ _32991_/Q _32927_/Q _32863_/Q _32799_/Q _18936_/X _18937_/X VGND VGND VPWR
+ VPWR _18976_/X sky130_fd_sc_hd__mux4_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _17923_/X _17926_/X _17853_/X VGND VGND VPWR VPWR _17937_/C sky130_fd_sc_hd__o21ba_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33973_ _34229_/CLK _33973_/D VGND VGND VPWR VPWR _33973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35712_ _35715_/CLK _35712_/D VGND VGND VPWR VPWR _35712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32924_ _34146_/CLK _32924_/D VGND VGND VPWR VPWR _32924_/Q sky130_fd_sc_hd__dfxtp_1
X_17858_ _17858_/A VGND VGND VPWR VPWR _17858_/X sky130_fd_sc_hd__buf_4
XFILLER_82_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35643_ _35772_/CLK _35643_/D VGND VGND VPWR VPWR _35643_/Q sky130_fd_sc_hd__dfxtp_1
X_16809_ _16800_/X _16807_/X _16808_/X VGND VGND VPWR VPWR _16810_/D sky130_fd_sc_hd__o21ba_1
XFILLER_54_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32855_ _33507_/CLK _32855_/D VGND VGND VPWR VPWR _32855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17789_ _35070_/Q _35006_/Q _34942_/Q _34878_/Q _17509_/X _17510_/X VGND VGND VPWR
+ VPWR _17789_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31806_ _31806_/A VGND VGND VPWR VPWR _36105_/D sky130_fd_sc_hd__clkbuf_1
X_19528_ _35054_/Q _34990_/Q _34926_/Q _34862_/Q _19456_/X _19457_/X VGND VGND VPWR
+ VPWR _19528_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35574_ _35574_/CLK _35574_/D VGND VGND VPWR VPWR _35574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32786_ _36052_/CLK _32786_/D VGND VGND VPWR VPWR _32786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_2_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_2_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_223_975 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34525_ _35036_/CLK _34525_/D VGND VGND VPWR VPWR _34525_/Q sky130_fd_sc_hd__dfxtp_1
X_19459_ _19459_/A VGND VGND VPWR VPWR _19459_/X sky130_fd_sc_hd__clkbuf_4
X_31737_ _31737_/A VGND VGND VPWR VPWR _36072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22470_ _22470_/A VGND VGND VPWR VPWR _36224_/D sky130_fd_sc_hd__clkbuf_1
X_34456_ _35738_/CLK _34456_/D VGND VGND VPWR VPWR _34456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31668_ _36040_/Q input54/X _31670_/S VGND VGND VPWR VPWR _31669_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33407_ _33789_/CLK _33407_/D VGND VGND VPWR VPWR _33407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21421_ _21302_/X _21419_/X _21420_/X _21308_/X VGND VGND VPWR VPWR _21421_/X sky130_fd_sc_hd__a22o_1
X_30619_ _30619_/A VGND VGND VPWR VPWR _35542_/D sky130_fd_sc_hd__clkbuf_1
X_34387_ _34967_/CLK _34387_/D VGND VGND VPWR VPWR _34387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31599_ _36007_/Q input18/X _31607_/S VGND VGND VPWR VPWR _31600_/A sky130_fd_sc_hd__mux2_1
X_21352_ _35745_/Q _35105_/Q _34465_/Q _33825_/Q _21034_/X _21035_/X VGND VGND VPWR
+ VPWR _21352_/X sky130_fd_sc_hd__mux4_1
X_24140_ _22923_/X _32604_/Q _24150_/S VGND VGND VPWR VPWR _24141_/A sky130_fd_sc_hd__mux2_1
X_36126_ _36127_/CLK _36126_/D VGND VGND VPWR VPWR _36126_/Q sky130_fd_sc_hd__dfxtp_1
X_33338_ _33787_/CLK _33338_/D VGND VGND VPWR VPWR _33338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20303_ _20303_/A _20303_/B _20303_/C _20303_/D VGND VGND VPWR VPWR _20304_/A sky130_fd_sc_hd__or4_2
X_24071_ _23022_/X _32572_/Q _24077_/S VGND VGND VPWR VPWR _24072_/A sky130_fd_sc_hd__mux2_1
X_36057_ _36121_/CLK _36057_/D VGND VGND VPWR VPWR _36057_/Q sky130_fd_sc_hd__dfxtp_1
X_21283_ _33183_/Q _32543_/Q _35935_/Q _35871_/Q _20968_/X _20969_/X VGND VGND VPWR
+ VPWR _21283_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33269_ _36149_/CLK _33269_/D VGND VGND VPWR VPWR _33269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20234_ _35074_/Q _35010_/Q _34946_/Q _34882_/Q _20162_/X _20163_/X VGND VGND VPWR
+ VPWR _20234_/X sky130_fd_sc_hd__mux4_1
X_35008_ _35075_/CLK _35008_/D VGND VGND VPWR VPWR _35008_/Q sky130_fd_sc_hd__dfxtp_1
X_23022_ input41/X VGND VGND VPWR VPWR _23022_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_190_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27830_ _27830_/A VGND VGND VPWR VPWR _34252_/D sky130_fd_sc_hd__clkbuf_1
X_20165_ _20165_/A VGND VGND VPWR VPWR _20165_/X sky130_fd_sc_hd__buf_4
XFILLER_131_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27761_ _27761_/A VGND VGND VPWR VPWR _34219_/D sky130_fd_sc_hd__clkbuf_1
X_20096_ _20096_/A VGND VGND VPWR VPWR _20096_/X sky130_fd_sc_hd__buf_4
X_24973_ _23053_/X _32966_/Q _24979_/S VGND VGND VPWR VPWR _24974_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29500_ _29500_/A VGND VGND VPWR VPWR _35012_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26712_ _26712_/A VGND VGND VPWR VPWR _33753_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23924_ _23924_/A VGND VGND VPWR VPWR _32502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27692_ _34187_/Q _24434_/X _27696_/S VGND VGND VPWR VPWR _27693_/A sky130_fd_sc_hd__mux2_1
XTAP_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29431_ _29431_/A VGND VGND VPWR VPWR _34979_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26643_ _26643_/A VGND VGND VPWR VPWR _33721_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23855_ _22904_/X _32470_/Q _23857_/S VGND VGND VPWR VPWR _23856_/A sky130_fd_sc_hd__mux2_1
XTAP_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_604 _18435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_615 _18505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_626 _18685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22806_ _34827_/Q _34763_/Q _34699_/Q _34635_/Q _22594_/X _22595_/X VGND VGND VPWR
+ VPWR _22806_/X sky130_fd_sc_hd__mux4_1
X_29362_ _23313_/X _34947_/Q _29374_/S VGND VGND VPWR VPWR _29363_/A sky130_fd_sc_hd__mux2_1
XANTENNA_637 _19211_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26574_ _26574_/A VGND VGND VPWR VPWR _33688_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23786_ _23834_/S VGND VGND VPWR VPWR _23805_/S sky130_fd_sc_hd__buf_4
XANTENNA_648 _19771_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_659 _20363_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20998_ _35799_/Q _32174_/Q _35671_/Q _35607_/Q _20854_/X _20855_/X VGND VGND VPWR
+ VPWR _20998_/X sky130_fd_sc_hd__mux4_1
X_28313_ _34481_/Q _24354_/X _28321_/S VGND VGND VPWR VPWR _28314_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25525_ _25525_/A VGND VGND VPWR VPWR _33194_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22737_ _21754_/A _22735_/X _22736_/X _21759_/A VGND VGND VPWR VPWR _22737_/X sky130_fd_sc_hd__a22o_1
X_29293_ _23148_/X _34914_/Q _29311_/S VGND VGND VPWR VPWR _29294_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28244_ _34448_/Q _24252_/X _28258_/S VGND VGND VPWR VPWR _28245_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25456_ _25183_/X _33164_/Q _25458_/S VGND VGND VPWR VPWR _25457_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22668_ _33543_/Q _33479_/Q _33415_/Q _33351_/Q _22429_/X _22430_/X VGND VGND VPWR
+ VPWR _22668_/X sky130_fd_sc_hd__mux4_2
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24407_ input48/X VGND VGND VPWR VPWR _24407_/X sky130_fd_sc_hd__buf_6
XFILLER_187_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21619_ _33513_/Q _33449_/Q _33385_/Q _33321_/Q _21370_/X _21371_/X VGND VGND VPWR
+ VPWR _21619_/X sky130_fd_sc_hd__mux4_1
X_28175_ _28175_/A VGND VGND VPWR VPWR _34415_/D sky130_fd_sc_hd__clkbuf_1
X_25387_ _25081_/X _33131_/Q _25387_/S VGND VGND VPWR VPWR _25388_/A sky130_fd_sc_hd__mux2_1
X_22599_ _34564_/Q _32452_/Q _34436_/Q _34372_/Q _22531_/X _22532_/X VGND VGND VPWR
+ VPWR _22599_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27126_ _27126_/A VGND VGND VPWR VPWR _33919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24338_ input24/X VGND VGND VPWR VPWR _24338_/X sky130_fd_sc_hd__clkbuf_8
X_27057_ _27057_/A VGND VGND VPWR VPWR _33886_/D sky130_fd_sc_hd__clkbuf_1
X_24269_ _24269_/A VGND VGND VPWR VPWR _32661_/D sky130_fd_sc_hd__clkbuf_1
X_26008_ _26008_/A VGND VGND VPWR VPWR _33421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1003 _17834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18830_ _33499_/Q _33435_/Q _33371_/Q _33307_/Q _18717_/X _18718_/X VGND VGND VPWR
+ VPWR _18830_/X sky130_fd_sc_hd__mux4_1
XTAP_6230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1014 _17842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1025 _17865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1036 _17152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1047 _17159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1058 _16458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18761_ _18436_/X _18759_/X _18760_/X _18441_/X VGND VGND VPWR VPWR _18761_/X sky130_fd_sc_hd__a22o_1
XTAP_6285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27959_ _27959_/A VGND VGND VPWR VPWR _34313_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1069 _17119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17712_ _17712_/A VGND VGND VPWR VPWR _17712_/X sky130_fd_sc_hd__buf_6
XFILLER_23_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30970_ _35709_/Q _29197_/X _30974_/S VGND VGND VPWR VPWR _30971_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18692_ _33239_/Q _36119_/Q _33111_/Q _33047_/Q _18652_/X _18653_/X VGND VGND VPWR
+ VPWR _18692_/X sky130_fd_sc_hd__mux4_1
XTAP_5595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29629_ _29629_/A VGND VGND VPWR VPWR _35073_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17643_ _34810_/Q _34746_/Q _34682_/Q _34618_/Q _17641_/X _17642_/X VGND VGND VPWR
+ VPWR _17643_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32640_ _36098_/CLK _32640_/D VGND VGND VPWR VPWR _32640_/Q sky130_fd_sc_hd__dfxtp_1
X_17574_ _17570_/X _17573_/X _17500_/X VGND VGND VPWR VPWR _17584_/C sky130_fd_sc_hd__o21ba_1
XFILLER_147_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19313_ _19309_/X _19312_/X _19108_/X VGND VGND VPWR VPWR _19314_/D sky130_fd_sc_hd__o21ba_1
X_16525_ _16525_/A _16525_/B _16525_/C _16525_/D VGND VGND VPWR VPWR _16526_/A sky130_fd_sc_hd__or4_2
XFILLER_205_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32571_ _35963_/CLK _32571_/D VGND VGND VPWR VPWR _32571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34310_ _34310_/CLK _34310_/D VGND VGND VPWR VPWR _34310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31522_ _31522_/A VGND VGND VPWR VPWR _35970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19244_ _19244_/A _19244_/B _19244_/C _19244_/D VGND VGND VPWR VPWR _19245_/A sky130_fd_sc_hd__or4_4
X_16456_ _16447_/X _16454_/X _16455_/X VGND VGND VPWR VPWR _16457_/D sky130_fd_sc_hd__o21ba_1
X_35290_ _35292_/CLK _35290_/D VGND VGND VPWR VPWR _35290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34241_ _36160_/CLK _34241_/D VGND VGND VPWR VPWR _34241_/Q sky130_fd_sc_hd__dfxtp_1
X_31453_ _31543_/S VGND VGND VPWR VPWR _31472_/S sky130_fd_sc_hd__buf_4
X_19175_ _35044_/Q _34980_/Q _34916_/Q _34852_/Q _19103_/X _19104_/X VGND VGND VPWR
+ VPWR _19175_/X sky130_fd_sc_hd__mux4_1
X_16387_ _33495_/Q _33431_/Q _33367_/Q _33303_/Q _15998_/X _15999_/X VGND VGND VPWR
+ VPWR _16387_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18126_ _34313_/Q _34249_/Q _34185_/Q _34121_/Q _16045_/X _16046_/X VGND VGND VPWR
+ VPWR _18126_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30404_ _30404_/A VGND VGND VPWR VPWR _35440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_247_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34172_ _36157_/CLK _34172_/D VGND VGND VPWR VPWR _34172_/Q sky130_fd_sc_hd__dfxtp_1
X_31384_ _35905_/Q input47/X _31400_/S VGND VGND VPWR VPWR _31385_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18057_ _35334_/Q _35270_/Q _35206_/Q _32326_/Q _16088_/X _16090_/X VGND VGND VPWR
+ VPWR _18057_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30335_ _30335_/A VGND VGND VPWR VPWR _35407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33123_ _36128_/CLK _33123_/D VGND VGND VPWR VPWR _33123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17008_ _35304_/Q _35240_/Q _35176_/Q _32296_/Q _17006_/X _17007_/X VGND VGND VPWR
+ VPWR _17008_/X sky130_fd_sc_hd__mux4_1
X_33054_ _36124_/CLK _33054_/D VGND VGND VPWR VPWR _33054_/Q sky130_fd_sc_hd__dfxtp_1
X_30266_ _30266_/A VGND VGND VPWR VPWR _35375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32005_ _36194_/CLK _32005_/D VGND VGND VPWR VPWR _32005_/Q sky130_fd_sc_hd__dfxtp_1
X_30197_ _30197_/A VGND VGND VPWR VPWR _35342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18959_ _18748_/X _18957_/X _18958_/X _18753_/X VGND VGND VPWR VPWR _18959_/X sky130_fd_sc_hd__a22o_1
XFILLER_230_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21970_ _34291_/Q _34227_/Q _34163_/Q _34099_/Q _21689_/X _21690_/X VGND VGND VPWR
+ VPWR _21970_/X sky130_fd_sc_hd__mux4_1
X_33956_ _34149_/CLK _33956_/D VGND VGND VPWR VPWR _33956_/Q sky130_fd_sc_hd__dfxtp_1
X_32907_ _36170_/CLK _32907_/D VGND VGND VPWR VPWR _32907_/Q sky130_fd_sc_hd__dfxtp_1
X_20921_ _20614_/X _20919_/X _20920_/X _20623_/X VGND VGND VPWR VPWR _20921_/X sky130_fd_sc_hd__a22o_1
XFILLER_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33887_ _34016_/CLK _33887_/D VGND VGND VPWR VPWR _33887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35626_ _35818_/CLK _35626_/D VGND VGND VPWR VPWR _35626_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23640_ _32370_/Q _23256_/X _23646_/S VGND VGND VPWR VPWR _23641_/A sky130_fd_sc_hd__mux2_1
X_32838_ _36039_/CLK _32838_/D VGND VGND VPWR VPWR _32838_/Q sky130_fd_sc_hd__dfxtp_1
X_20852_ _20626_/X _20850_/X _20851_/X _20637_/X VGND VGND VPWR VPWR _20852_/X sky130_fd_sc_hd__a22o_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23571_ _32337_/Q _23096_/X _23583_/S VGND VGND VPWR VPWR _23572_/A sky130_fd_sc_hd__mux2_1
X_35557_ _35749_/CLK _35557_/D VGND VGND VPWR VPWR _35557_/Q sky130_fd_sc_hd__dfxtp_1
X_32769_ _36098_/CLK _32769_/D VGND VGND VPWR VPWR _32769_/Q sky130_fd_sc_hd__dfxtp_1
X_20783_ _20614_/X _20781_/X _20782_/X _20623_/X VGND VGND VPWR VPWR _20783_/X sky130_fd_sc_hd__a22o_1
XFILLER_195_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25310_ _25168_/X _33095_/Q _25314_/S VGND VGND VPWR VPWR _25311_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34508_ _35853_/CLK _34508_/D VGND VGND VPWR VPWR _34508_/Q sky130_fd_sc_hd__dfxtp_1
X_22522_ _35778_/Q _35138_/Q _34498_/Q _33858_/Q _22446_/X _22447_/X VGND VGND VPWR
+ VPWR _22522_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26290_ _26290_/A VGND VGND VPWR VPWR _33554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35488_ _35552_/CLK _35488_/D VGND VGND VPWR VPWR _35488_/Q sky130_fd_sc_hd__dfxtp_1
X_25241_ _25066_/X _33062_/Q _25251_/S VGND VGND VPWR VPWR _25242_/A sky130_fd_sc_hd__mux2_1
X_34439_ _35078_/CLK _34439_/D VGND VGND VPWR VPWR _34439_/Q sky130_fd_sc_hd__dfxtp_1
X_22453_ _22453_/A VGND VGND VPWR VPWR _22453_/X sky130_fd_sc_hd__buf_2
XFILLER_206_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21404_ _21757_/A VGND VGND VPWR VPWR _21404_/X sky130_fd_sc_hd__buf_4
X_25172_ _25171_/X _33032_/Q _25175_/S VGND VGND VPWR VPWR _25173_/A sky130_fd_sc_hd__mux2_1
XFILLER_202_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22384_ _22378_/X _22383_/X _22100_/X VGND VGND VPWR VPWR _22392_/C sky130_fd_sc_hd__o21ba_1
XFILLER_159_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36109_ _36109_/CLK _36109_/D VGND VGND VPWR VPWR _36109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24123_ _22898_/X _32596_/Q _24129_/S VGND VGND VPWR VPWR _24124_/A sky130_fd_sc_hd__mux2_1
X_21335_ _33761_/Q _33697_/Q _33633_/Q _33569_/Q _21090_/X _21091_/X VGND VGND VPWR
+ VPWR _21335_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29980_ _35240_/Q _29132_/X _29986_/S VGND VGND VPWR VPWR _29981_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28931_ _34774_/Q _24270_/X _28933_/S VGND VGND VPWR VPWR _28932_/A sky130_fd_sc_hd__mux2_1
X_24054_ _22997_/X _32564_/Q _24056_/S VGND VGND VPWR VPWR _24055_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21266_ _33503_/Q _33439_/Q _33375_/Q _33311_/Q _21017_/X _21018_/X VGND VGND VPWR
+ VPWR _21266_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23005_ _23003_/X _32054_/Q _23032_/S VGND VGND VPWR VPWR _23006_/A sky130_fd_sc_hd__mux2_1
X_20217_ _32514_/Q _32386_/Q _32066_/Q _36034_/Q _19929_/X _20070_/X VGND VGND VPWR
+ VPWR _20217_/X sky130_fd_sc_hd__mux4_1
X_28862_ _28862_/A VGND VGND VPWR VPWR _34741_/D sky130_fd_sc_hd__clkbuf_1
X_21197_ _34013_/Q _33949_/Q _33885_/Q _32157_/Q _20914_/X _20915_/X VGND VGND VPWR
+ VPWR _21197_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27813_ _34244_/Q _24413_/X _27823_/S VGND VGND VPWR VPWR _27814_/A sky130_fd_sc_hd__mux2_1
X_20148_ _35776_/Q _35136_/Q _34496_/Q _33856_/Q _20146_/X _20147_/X VGND VGND VPWR
+ VPWR _20148_/X sky130_fd_sc_hd__mux4_1
X_28793_ _28793_/A VGND VGND VPWR VPWR _34708_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20079_ _35582_/Q _35518_/Q _35454_/Q _35390_/Q _19903_/X _19904_/X VGND VGND VPWR
+ VPWR _20079_/X sky130_fd_sc_hd__mux4_1
X_24956_ _23028_/X _32958_/Q _24958_/S VGND VGND VPWR VPWR _24957_/A sky130_fd_sc_hd__mux2_1
XTAP_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27744_ _34211_/Q _24311_/X _27760_/S VGND VGND VPWR VPWR _27745_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23907_ _23907_/A VGND VGND VPWR VPWR _32494_/D sky130_fd_sc_hd__clkbuf_1
X_27675_ _27675_/A VGND VGND VPWR VPWR _34178_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24887_ _22926_/X _32925_/Q _24895_/S VGND VGND VPWR VPWR _24888_/A sky130_fd_sc_hd__mux2_1
XANTENNA_401 _36210_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_412 _36212_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29414_ _29414_/A VGND VGND VPWR VPWR _34971_/D sky130_fd_sc_hd__clkbuf_1
X_26626_ _26626_/A VGND VGND VPWR VPWR _33713_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23838_ _23970_/S VGND VGND VPWR VPWR _23857_/S sky130_fd_sc_hd__buf_4
XTAP_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_423 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_434 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_445 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_456 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_467 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26557_ _26557_/A VGND VGND VPWR VPWR _33680_/D sky130_fd_sc_hd__clkbuf_1
X_29345_ _23286_/X _34939_/Q _29353_/S VGND VGND VPWR VPWR _29346_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23769_ _23769_/A VGND VGND VPWR VPWR _32429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_478 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_489 _31994_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16310_ _33749_/Q _33685_/Q _33621_/Q _33557_/Q _16137_/X _16138_/X VGND VGND VPWR
+ VPWR _16310_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25508_ _33186_/Q _24307_/X _25526_/S VGND VGND VPWR VPWR _25509_/A sky130_fd_sc_hd__mux2_1
XFILLER_242_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29276_ _23124_/X _34906_/Q _29290_/S VGND VGND VPWR VPWR _29277_/A sky130_fd_sc_hd__mux2_1
X_17290_ _34800_/Q _34736_/Q _34672_/Q _34608_/Q _17288_/X _17289_/X VGND VGND VPWR
+ VPWR _17290_/X sky130_fd_sc_hd__mux4_1
X_26488_ _26488_/A VGND VGND VPWR VPWR _33648_/D sky130_fd_sc_hd__clkbuf_1
X_28227_ _28227_/A VGND VGND VPWR VPWR _34440_/D sky130_fd_sc_hd__clkbuf_1
X_16241_ _34259_/Q _34195_/Q _34131_/Q _34067_/Q _16005_/X _16007_/X VGND VGND VPWR
+ VPWR _16241_/X sky130_fd_sc_hd__mux4_1
X_25439_ _25439_/A VGND VGND VPWR VPWR _33155_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16172_ _16172_/A _16172_/B _16172_/C _16172_/D VGND VGND VPWR VPWR _16173_/A sky130_fd_sc_hd__or4_4
X_28158_ _28158_/A VGND VGND VPWR VPWR _34407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27109_ _26950_/X _33911_/Q _27125_/S VGND VGND VPWR VPWR _27110_/A sky130_fd_sc_hd__mux2_1
X_28089_ _26999_/X _34375_/Q _28093_/S VGND VGND VPWR VPWR _28090_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30120_ _30120_/A VGND VGND VPWR VPWR _35306_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19931_ _33018_/Q _32954_/Q _32890_/Q _32826_/Q _19642_/X _19643_/X VGND VGND VPWR
+ VPWR _19931_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30051_ _35274_/Q _29237_/X _30057_/S VGND VGND VPWR VPWR _30052_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19862_ _33272_/Q _36152_/Q _33144_/Q _33080_/Q _19711_/X _19712_/X VGND VGND VPWR
+ VPWR _19862_/X sky130_fd_sc_hd__mux4_1
XFILLER_218_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput92 _31961_/Q VGND VGND VPWR VPWR D1[11] sky130_fd_sc_hd__buf_2
X_18813_ _33178_/Q _32538_/Q _35930_/Q _35866_/Q _18668_/X _18669_/X VGND VGND VPWR
+ VPWR _18813_/X sky130_fd_sc_hd__mux4_1
XTAP_6060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19793_ _20146_/A VGND VGND VPWR VPWR _19793_/X sky130_fd_sc_hd__buf_4
XTAP_6082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33810_ _35730_/CLK _33810_/D VGND VGND VPWR VPWR _33810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18744_ _34776_/Q _34712_/Q _34648_/Q _34584_/Q _18529_/X _18530_/X VGND VGND VPWR
+ VPWR _18744_/X sky130_fd_sc_hd__mux4_1
XTAP_5370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34790_ _34922_/CLK _34790_/D VGND VGND VPWR VPWR _34790_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33741_ _36112_/CLK _33741_/D VGND VGND VPWR VPWR _33741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18675_ _18374_/X _18673_/X _18674_/X _18384_/X VGND VGND VPWR VPWR _18675_/X sky130_fd_sc_hd__a22o_1
X_30953_ _35701_/Q _29172_/X _30953_/S VGND VGND VPWR VPWR _30954_/A sky130_fd_sc_hd__mux2_1
XFILLER_237_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17626_ _32762_/Q _32698_/Q _32634_/Q _36090_/Q _17625_/X _17409_/X VGND VGND VPWR
+ VPWR _17626_/X sky130_fd_sc_hd__mux4_1
X_33672_ _34817_/CLK _33672_/D VGND VGND VPWR VPWR _33672_/Q sky130_fd_sc_hd__dfxtp_1
X_30884_ _35668_/Q _29070_/X _30890_/S VGND VGND VPWR VPWR _30885_/A sky130_fd_sc_hd__mux2_1
XTAP_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35411_ _35922_/CLK _35411_/D VGND VGND VPWR VPWR _35411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32623_ _36078_/CLK _32623_/D VGND VGND VPWR VPWR _32623_/Q sky130_fd_sc_hd__dfxtp_1
X_17557_ _34040_/Q _33976_/Q _33912_/Q _32248_/Q _17373_/X _17374_/X VGND VGND VPWR
+ VPWR _17557_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_990 _17860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35342_ _35793_/CLK _35342_/D VGND VGND VPWR VPWR _35342_/Q sky130_fd_sc_hd__dfxtp_1
X_16508_ _16504_/X _16507_/X _16430_/X _16431_/X VGND VGND VPWR VPWR _16525_/B sky130_fd_sc_hd__o211a_2
X_32554_ _35947_/CLK _32554_/D VGND VGND VPWR VPWR _32554_/Q sky130_fd_sc_hd__dfxtp_1
X_17488_ _17416_/X _17486_/X _17487_/X _17420_/X VGND VGND VPWR VPWR _17488_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31505_ _31505_/A VGND VGND VPWR VPWR _35962_/D sky130_fd_sc_hd__clkbuf_1
X_19227_ _19222_/X _19226_/X _19083_/X _19084_/X VGND VGND VPWR VPWR _19244_/B sky130_fd_sc_hd__o211a_1
X_35273_ _35273_/CLK _35273_/D VGND VGND VPWR VPWR _35273_/Q sky130_fd_sc_hd__dfxtp_1
X_16439_ _33176_/Q _32536_/Q _35928_/Q _35864_/Q _16368_/X _16369_/X VGND VGND VPWR
+ VPWR _16439_/X sky130_fd_sc_hd__mux4_1
X_32485_ _36005_/CLK _32485_/D VGND VGND VPWR VPWR _32485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34224_ _34291_/CLK _34224_/D VGND VGND VPWR VPWR _34224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31436_ _31436_/A VGND VGND VPWR VPWR _35929_/D sky130_fd_sc_hd__clkbuf_1
X_19158_ _32484_/Q _32356_/Q _32036_/Q _36004_/Q _18870_/X _19011_/X VGND VGND VPWR
+ VPWR _19158_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18109_ _35848_/Q _32228_/Q _35720_/Q _35656_/Q _15989_/X _15991_/X VGND VGND VPWR
+ VPWR _18109_/X sky130_fd_sc_hd__mux4_1
X_31367_ _35897_/Q input38/X _31379_/S VGND VGND VPWR VPWR _31368_/A sky130_fd_sc_hd__mux2_1
X_34155_ _34282_/CLK _34155_/D VGND VGND VPWR VPWR _34155_/Q sky130_fd_sc_hd__dfxtp_1
X_19089_ _35746_/Q _35106_/Q _34466_/Q _33826_/Q _19087_/X _19088_/X VGND VGND VPWR
+ VPWR _19089_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30318_ _30318_/A VGND VGND VPWR VPWR _35400_/D sky130_fd_sc_hd__clkbuf_1
X_33106_ _36114_/CLK _33106_/D VGND VGND VPWR VPWR _33106_/Q sky130_fd_sc_hd__dfxtp_1
X_21120_ _21473_/A VGND VGND VPWR VPWR _21120_/X sky130_fd_sc_hd__buf_4
X_31298_ _35864_/Q input2/X _31316_/S VGND VGND VPWR VPWR _31299_/A sky130_fd_sc_hd__mux2_1
X_34086_ _34087_/CLK _34086_/D VGND VGND VPWR VPWR _34086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21051_ _21757_/A VGND VGND VPWR VPWR _21051_/X sky130_fd_sc_hd__buf_4
X_33037_ _34317_/CLK _33037_/D VGND VGND VPWR VPWR _33037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30249_ _30249_/A VGND VGND VPWR VPWR _35367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20002_ _35772_/Q _35132_/Q _34492_/Q _33852_/Q _19793_/X _19794_/X VGND VGND VPWR
+ VPWR _20002_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_1239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24810_ _24810_/A VGND VGND VPWR VPWR _32888_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25790_ _25790_/A VGND VGND VPWR VPWR _33317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_246_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34988_ _35052_/CLK _34988_/D VGND VGND VPWR VPWR _34988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24741_ _24852_/S VGND VGND VPWR VPWR _24760_/S sky130_fd_sc_hd__buf_4
X_33939_ _36228_/CLK _33939_/D VGND VGND VPWR VPWR _33939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21953_ _35570_/Q _35506_/Q _35442_/Q _35378_/Q _21850_/X _21851_/X VGND VGND VPWR
+ VPWR _21953_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20904_ _34516_/Q _32404_/Q _34388_/Q _34324_/Q _20766_/X _20767_/X VGND VGND VPWR
+ VPWR _20904_/X sky130_fd_sc_hd__mux4_1
X_27460_ _27460_/A VGND VGND VPWR VPWR _34077_/D sky130_fd_sc_hd__clkbuf_1
X_24672_ _23010_/X _32824_/Q _24686_/S VGND VGND VPWR VPWR _24673_/A sky130_fd_sc_hd__mux2_1
X_21884_ _35568_/Q _35504_/Q _35440_/Q _35376_/Q _21850_/X _21851_/X VGND VGND VPWR
+ VPWR _21884_/X sky130_fd_sc_hd__mux4_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26411_ _26411_/A VGND VGND VPWR VPWR _33612_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23623_ _32362_/Q _23231_/X _23625_/S VGND VGND VPWR VPWR _23624_/A sky130_fd_sc_hd__mux2_1
X_35609_ _36063_/CLK _35609_/D VGND VGND VPWR VPWR _35609_/Q sky130_fd_sc_hd__dfxtp_1
X_20835_ _35026_/Q _34962_/Q _34898_/Q _34834_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _20835_/X sky130_fd_sc_hd__mux4_1
X_27391_ _34045_/Q _24391_/X _27395_/S VGND VGND VPWR VPWR _27392_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29130_ _34855_/Q _29129_/X _29142_/S VGND VGND VPWR VPWR _29131_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26342_ _26342_/A VGND VGND VPWR VPWR _33579_/D sky130_fd_sc_hd__clkbuf_1
X_23554_ _23554_/A VGND VGND VPWR VPWR _32330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20766_ _22312_/A VGND VGND VPWR VPWR _20766_/X sky130_fd_sc_hd__buf_6
X_22505_ _34306_/Q _34242_/Q _34178_/Q _34114_/Q _22395_/X _22396_/X VGND VGND VPWR
+ VPWR _22505_/X sky130_fd_sc_hd__mux4_1
X_29061_ input34/X VGND VGND VPWR VPWR _29061_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26273_ _25180_/X _33547_/Q _26277_/S VGND VGND VPWR VPWR _26274_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23485_ _23485_/A VGND VGND VPWR VPWR _32297_/D sky130_fd_sc_hd__clkbuf_1
X_20697_ _21759_/A VGND VGND VPWR VPWR _20697_/X sky130_fd_sc_hd__clkbuf_4
X_28012_ _26884_/X _34338_/Q _28030_/S VGND VGND VPWR VPWR _28013_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25224_ _25041_/X _33054_/Q _25230_/S VGND VGND VPWR VPWR _25225_/A sky130_fd_sc_hd__mux2_1
X_22436_ _32768_/Q _32704_/Q _32640_/Q _36096_/Q _22225_/X _22362_/X VGND VGND VPWR
+ VPWR _22436_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25155_ _25155_/A VGND VGND VPWR VPWR _33026_/D sky130_fd_sc_hd__clkbuf_1
X_22367_ _22367_/A VGND VGND VPWR VPWR _22367_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_191_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _35583_/CLK sky130_fd_sc_hd__clkbuf_16
X_24106_ _23074_/X _32589_/Q _24106_/S VGND VGND VPWR VPWR _24107_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21318_ _35744_/Q _35104_/Q _34464_/Q _33824_/Q _21034_/X _21035_/X VGND VGND VPWR
+ VPWR _21318_/X sky130_fd_sc_hd__mux4_1
X_29963_ _35232_/Q _29107_/X _29965_/S VGND VGND VPWR VPWR _29964_/A sky130_fd_sc_hd__mux2_1
X_25086_ _25084_/X _33004_/Q _25113_/S VGND VGND VPWR VPWR _25087_/A sky130_fd_sc_hd__mux2_1
X_22298_ _22016_/X _22294_/X _22297_/X _22020_/X VGND VGND VPWR VPWR _22298_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28914_ _29046_/S VGND VGND VPWR VPWR _28933_/S sky130_fd_sc_hd__buf_4
X_24037_ _24106_/S VGND VGND VPWR VPWR _24056_/S sky130_fd_sc_hd__buf_6
XFILLER_85_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21249_ _22465_/A VGND VGND VPWR VPWR _21249_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_105_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29894_ _29894_/A VGND VGND VPWR VPWR _35199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28845_ _26919_/X _34733_/Q _28861_/S VGND VGND VPWR VPWR _28846_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16790_ _16641_/X _16786_/X _16789_/X _16644_/X VGND VGND VPWR VPWR _16790_/X sky130_fd_sc_hd__a22o_1
X_28776_ _27017_/X _34701_/Q _28776_/S VGND VGND VPWR VPWR _28777_/A sky130_fd_sc_hd__mux2_1
X_25988_ _25988_/A VGND VGND VPWR VPWR _33411_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_891 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24939_ _24987_/S VGND VGND VPWR VPWR _24958_/S sky130_fd_sc_hd__buf_4
X_27727_ _34203_/Q _24286_/X _27739_/S VGND VGND VPWR VPWR _27728_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18460_ _33168_/Q _32528_/Q _35920_/Q _35856_/Q _18363_/X _18365_/X VGND VGND VPWR
+ VPWR _18460_/X sky130_fd_sc_hd__mux4_1
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27658_ _27658_/A VGND VGND VPWR VPWR _34170_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_220 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_231 _32136_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_242 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _17982_/A VGND VGND VPWR VPWR _17411_/X sky130_fd_sc_hd__buf_4
X_18391_ _34510_/Q _32398_/Q _34382_/Q _34318_/Q _18388_/X _18390_/X VGND VGND VPWR
+ VPWR _18391_/X sky130_fd_sc_hd__mux4_1
X_26609_ _26609_/A VGND VGND VPWR VPWR _33705_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_253 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_264 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27589_ _27589_/A VGND VGND VPWR VPWR _34137_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_275 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_286 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17829_/A VGND VGND VPWR VPWR _17342_/X sky130_fd_sc_hd__buf_4
XANTENNA_297 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29328_ _23261_/X _34931_/Q _29332_/S VGND VGND VPWR VPWR _29329_/A sky130_fd_sc_hd__mux2_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17273_ _32752_/Q _32688_/Q _32624_/Q _36080_/Q _17272_/X _17056_/X VGND VGND VPWR
+ VPWR _17273_/X sky130_fd_sc_hd__mux4_1
X_29259_ _23099_/X _34898_/Q _29269_/S VGND VGND VPWR VPWR _29260_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16224_ _16044_/X _16222_/X _16223_/X _16054_/X VGND VGND VPWR VPWR _16224_/X sky130_fd_sc_hd__a22o_1
X_19012_ _32480_/Q _32352_/Q _32032_/Q _36000_/Q _18870_/X _19011_/X VGND VGND VPWR
+ VPWR _19012_/X sky130_fd_sc_hd__mux4_1
X_32270_ _36216_/CLK _32270_/D VGND VGND VPWR VPWR _32270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31221_ _35828_/Q input32/X _31223_/S VGND VGND VPWR VPWR _31222_/A sky130_fd_sc_hd__mux2_1
X_16155_ _16151_/X _16154_/X _16040_/X _16042_/X VGND VGND VPWR VPWR _16172_/B sky130_fd_sc_hd__o211a_1
XFILLER_31_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_182_CLK clkbuf_leaf_66_CLK/A VGND VGND VPWR VPWR _32978_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_115_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31152_ _35795_/Q input56/X _31160_/S VGND VGND VPWR VPWR _31153_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16086_ _17769_/A VGND VGND VPWR VPWR _17154_/A sky130_fd_sc_hd__buf_12
XFILLER_138_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30103_ _35298_/Q _29113_/X _30121_/S VGND VGND VPWR VPWR _30104_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19914_ _19807_/X _19912_/X _19913_/X _19812_/X VGND VGND VPWR VPWR _19914_/X sky130_fd_sc_hd__a22o_1
X_35960_ _36024_/CLK _35960_/D VGND VGND VPWR VPWR _35960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31083_ _31083_/A VGND VGND VPWR VPWR _35762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30034_ _30034_/A VGND VGND VPWR VPWR _35265_/D sky130_fd_sc_hd__clkbuf_1
X_34911_ _35040_/CLK _34911_/D VGND VGND VPWR VPWR _34911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19845_ _19841_/X _19844_/X _19814_/X VGND VGND VPWR VPWR _19846_/D sky130_fd_sc_hd__o21ba_1
XFILLER_155_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35891_ _35955_/CLK _35891_/D VGND VGND VPWR VPWR _35891_/Q sky130_fd_sc_hd__dfxtp_1
X_34842_ _35034_/CLK _34842_/D VGND VGND VPWR VPWR _34842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19776_ _20129_/A VGND VGND VPWR VPWR _19776_/X sky130_fd_sc_hd__buf_4
X_16988_ _32488_/Q _32360_/Q _32040_/Q _36008_/Q _16923_/X _16711_/X VGND VGND VPWR
+ VPWR _16988_/X sky130_fd_sc_hd__mux4_1
X_18727_ _32472_/Q _32344_/Q _32024_/Q _35992_/Q _18517_/X _18658_/X VGND VGND VPWR
+ VPWR _18727_/X sky130_fd_sc_hd__mux4_1
XFILLER_225_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34773_ _34775_/CLK _34773_/D VGND VGND VPWR VPWR _34773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31985_ _36201_/CLK _31985_/D VGND VGND VPWR VPWR _31985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33724_ _34044_/CLK _33724_/D VGND VGND VPWR VPWR _33724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18658_ _20070_/A VGND VGND VPWR VPWR _18658_/X sky130_fd_sc_hd__buf_4
X_30936_ _30936_/A VGND VGND VPWR VPWR _35692_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17609_ _34809_/Q _34745_/Q _34681_/Q _34617_/Q _17288_/X _17289_/X VGND VGND VPWR
+ VPWR _17609_/X sky130_fd_sc_hd__mux4_1
X_33655_ _34295_/CLK _33655_/D VGND VGND VPWR VPWR _33655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30867_ _30867_/A VGND VGND VPWR VPWR _35660_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18589_ _35796_/Q _32170_/Q _35668_/Q _35604_/Q _18554_/X _18555_/X VGND VGND VPWR
+ VPWR _18589_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20620_ _22502_/A VGND VGND VPWR VPWR _20620_/X sky130_fd_sc_hd__buf_4
X_32606_ _36062_/CLK _32606_/D VGND VGND VPWR VPWR _32606_/Q sky130_fd_sc_hd__dfxtp_1
X_33586_ _34289_/CLK _33586_/D VGND VGND VPWR VPWR _33586_/Q sky130_fd_sc_hd__dfxtp_1
X_30798_ _30798_/A VGND VGND VPWR VPWR _35627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35325_ _35326_/CLK _35325_/D VGND VGND VPWR VPWR _35325_/Q sky130_fd_sc_hd__dfxtp_1
X_20551_ _20547_/X _20550_/X _20134_/A VGND VGND VPWR VPWR _20573_/A sky130_fd_sc_hd__o21ba_1
XFILLER_123_1328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32537_ _35929_/CLK _32537_/D VGND VGND VPWR VPWR _32537_/Q sky130_fd_sc_hd__dfxtp_1
X_35256_ _35320_/CLK _35256_/D VGND VGND VPWR VPWR _35256_/Q sky130_fd_sc_hd__dfxtp_1
X_23270_ input35/X VGND VGND VPWR VPWR _23270_/X sky130_fd_sc_hd__buf_4
X_20482_ _20478_/X _20481_/X _20167_/A VGND VGND VPWR VPWR _20483_/D sky130_fd_sc_hd__o21ba_1
X_32468_ _35989_/CLK _32468_/D VGND VGND VPWR VPWR _32468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22221_ _33530_/Q _33466_/Q _33402_/Q _33338_/Q _22076_/X _22077_/X VGND VGND VPWR
+ VPWR _22221_/X sky130_fd_sc_hd__mux4_1
X_34207_ _35675_/CLK _34207_/D VGND VGND VPWR VPWR _34207_/Q sky130_fd_sc_hd__dfxtp_1
X_31419_ _31419_/A VGND VGND VPWR VPWR _35921_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_173_CLK clkbuf_leaf_76_CLK/A VGND VGND VPWR VPWR _36048_/CLK sky130_fd_sc_hd__clkbuf_16
X_35187_ _35187_/CLK _35187_/D VGND VGND VPWR VPWR _35187_/Q sky130_fd_sc_hd__dfxtp_1
X_32399_ _34638_/CLK _32399_/D VGND VGND VPWR VPWR _32399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22152_ _34296_/Q _34232_/Q _34168_/Q _34104_/Q _22042_/X _22043_/X VGND VGND VPWR
+ VPWR _22152_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34138_ _34202_/CLK _34138_/D VGND VGND VPWR VPWR _34138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21103_ _33242_/Q _36122_/Q _33114_/Q _33050_/Q _20952_/X _20953_/X VGND VGND VPWR
+ VPWR _21103_/X sky130_fd_sc_hd__mux4_1
XTAP_6818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34069_ _34197_/CLK _34069_/D VGND VGND VPWR VPWR _34069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26960_ _26959_/X _33850_/Q _26975_/S VGND VGND VPWR VPWR _26961_/A sky130_fd_sc_hd__mux2_1
X_22083_ _32758_/Q _32694_/Q _32630_/Q _36086_/Q _21872_/X _22009_/X VGND VGND VPWR
+ VPWR _22083_/X sky130_fd_sc_hd__mux4_1
XTAP_6829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21034_ _22594_/A VGND VGND VPWR VPWR _21034_/X sky130_fd_sc_hd__buf_6
X_25911_ _25044_/X _33375_/Q _25915_/S VGND VGND VPWR VPWR _25912_/A sky130_fd_sc_hd__mux2_1
X_26891_ input15/X VGND VGND VPWR VPWR _26891_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_248_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28630_ _28630_/A VGND VGND VPWR VPWR _34631_/D sky130_fd_sc_hd__clkbuf_1
X_25842_ _25842_/A VGND VGND VPWR VPWR _33342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_44__f_CLK clkbuf_5_22_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_44__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_75_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28561_ _28561_/A VGND VGND VPWR VPWR _34598_/D sky130_fd_sc_hd__clkbuf_1
X_25773_ _25773_/A VGND VGND VPWR VPWR _33309_/D sky130_fd_sc_hd__clkbuf_1
X_22985_ input28/X VGND VGND VPWR VPWR _22985_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_167_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24724_ _24724_/A VGND VGND VPWR VPWR _32847_/D sky130_fd_sc_hd__clkbuf_1
X_27512_ _26946_/X _34102_/Q _27530_/S VGND VGND VPWR VPWR _27513_/A sky130_fd_sc_hd__mux2_1
X_28492_ _26996_/X _34566_/Q _28498_/S VGND VGND VPWR VPWR _28493_/A sky130_fd_sc_hd__mux2_1
X_21936_ _21802_/X _21934_/X _21935_/X _21805_/X VGND VGND VPWR VPWR _21936_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27443_ _27443_/A VGND VGND VPWR VPWR _34069_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24655_ _22985_/X _32816_/Q _24665_/S VGND VGND VPWR VPWR _24656_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21867_ _21795_/X _21865_/X _21866_/X _21800_/X VGND VGND VPWR VPWR _21867_/X sky130_fd_sc_hd__a22o_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23606_ _23696_/S VGND VGND VPWR VPWR _23625_/S sky130_fd_sc_hd__buf_4
XFILLER_243_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20818_ _32466_/Q _32338_/Q _32018_/Q _35986_/Q _20817_/X _22463_/A VGND VGND VPWR
+ VPWR _20818_/X sky130_fd_sc_hd__mux4_1
X_27374_ _34037_/Q _24366_/X _27374_/S VGND VGND VPWR VPWR _27375_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24586_ _22883_/X _32783_/Q _24602_/S VGND VGND VPWR VPWR _24587_/A sky130_fd_sc_hd__mux2_1
X_21798_ _33774_/Q _33710_/Q _33646_/Q _33582_/Q _21796_/X _21797_/X VGND VGND VPWR
+ VPWR _21798_/X sky130_fd_sc_hd__mux4_1
X_26325_ _25057_/X _33571_/Q _26341_/S VGND VGND VPWR VPWR _26326_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29113_ input13/X VGND VGND VPWR VPWR _29113_/X sky130_fd_sc_hd__buf_2
X_23537_ _23041_/X _32322_/Q _23551_/S VGND VGND VPWR VPWR _23538_/A sky130_fd_sc_hd__mux2_1
XFILLER_204_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20749_ _32720_/Q _32656_/Q _32592_/Q _36048_/Q _22462_/A _22313_/A VGND VGND VPWR
+ VPWR _20749_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29044_ _34828_/Q _24437_/X _29046_/S VGND VGND VPWR VPWR _29045_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26256_ _26256_/A VGND VGND VPWR VPWR _33538_/D sky130_fd_sc_hd__clkbuf_1
X_23468_ _23468_/A VGND VGND VPWR VPWR _32289_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25207_ _25016_/X _33046_/Q _25209_/S VGND VGND VPWR VPWR _25208_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22419_ _22102_/X _22417_/X _22418_/X _22105_/X VGND VGND VPWR VPWR _22419_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_164_CLK clkbuf_6_30__f_CLK/X VGND VGND VPWR VPWR _36170_/CLK sky130_fd_sc_hd__clkbuf_16
X_26187_ _26277_/S VGND VGND VPWR VPWR _26206_/S sky130_fd_sc_hd__buf_4
XFILLER_6_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23399_ _32258_/Q _23310_/X _23413_/S VGND VGND VPWR VPWR _23400_/A sky130_fd_sc_hd__mux2_1
X_25138_ _25137_/X _33021_/Q _25144_/S VGND VGND VPWR VPWR _25139_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_1324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17960_ _17705_/X _17958_/X _17959_/X _17708_/X VGND VGND VPWR VPWR _17960_/X sky130_fd_sc_hd__a22o_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29946_ _30057_/S VGND VGND VPWR VPWR _29965_/S sky130_fd_sc_hd__buf_4
X_25069_ input18/X VGND VGND VPWR VPWR _25069_/X sky130_fd_sc_hd__buf_2
XFILLER_78_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16911_ _16911_/A VGND VGND VPWR VPWR _31973_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17891_ _17887_/X _17890_/X _17853_/X VGND VGND VPWR VPWR _17899_/C sky130_fd_sc_hd__o21ba_1
XFILLER_120_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29877_ _35191_/Q _29179_/X _29893_/S VGND VGND VPWR VPWR _29878_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19630_ _19630_/A VGND VGND VPWR VPWR _32113_/D sky130_fd_sc_hd__buf_2
XFILLER_215_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28828_ _26894_/X _34725_/Q _28840_/S VGND VGND VPWR VPWR _28829_/A sky130_fd_sc_hd__mux2_1
X_16842_ _17901_/A VGND VGND VPWR VPWR _16842_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_93_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19561_ _19454_/X _19559_/X _19560_/X _19459_/X VGND VGND VPWR VPWR _19561_/X sky130_fd_sc_hd__a22o_1
X_28759_ _28759_/A VGND VGND VPWR VPWR _34692_/D sky130_fd_sc_hd__clkbuf_1
X_16773_ _34018_/Q _33954_/Q _33890_/Q _32162_/Q _16667_/X _16668_/X VGND VGND VPWR
+ VPWR _16773_/X sky130_fd_sc_hd__mux4_1
XFILLER_234_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18512_ _18508_/X _18511_/X _18311_/X VGND VGND VPWR VPWR _18538_/A sky130_fd_sc_hd__o21ba_1
XFILLER_59_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31770_ _36088_/Q input37/X _31784_/S VGND VGND VPWR VPWR _31771_/A sky130_fd_sc_hd__mux2_1
X_19492_ _19488_/X _19491_/X _19461_/X VGND VGND VPWR VPWR _19493_/D sky130_fd_sc_hd__o21ba_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30721_ _35591_/Q _29228_/X _30725_/S VGND VGND VPWR VPWR _30722_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18443_ _20160_/A VGND VGND VPWR VPWR _18443_/X sky130_fd_sc_hd__buf_4
XFILLER_18_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33440_ _34017_/CLK _33440_/D VGND VGND VPWR VPWR _33440_/Q sky130_fd_sc_hd__dfxtp_1
X_18374_ _19449_/A VGND VGND VPWR VPWR _18374_/X sky130_fd_sc_hd__buf_4
X_30652_ _35558_/Q _29126_/X _30662_/S VGND VGND VPWR VPWR _30653_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _34545_/Q _32433_/Q _34417_/Q _34353_/Q _17225_/X _17226_/X VGND VGND VPWR
+ VPWR _17325_/X sky130_fd_sc_hd__mux4_1
X_30583_ _30583_/A VGND VGND VPWR VPWR _35525_/D sky130_fd_sc_hd__clkbuf_1
X_33371_ _36194_/CLK _33371_/D VGND VGND VPWR VPWR _33371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35110_ _35750_/CLK _35110_/D VGND VGND VPWR VPWR _35110_/Q sky130_fd_sc_hd__dfxtp_1
X_32322_ _35330_/CLK _32322_/D VGND VGND VPWR VPWR _32322_/Q sky130_fd_sc_hd__dfxtp_1
X_36090_ _36090_/CLK _36090_/D VGND VGND VPWR VPWR _36090_/Q sky130_fd_sc_hd__dfxtp_1
X_17256_ _34799_/Q _34735_/Q _34671_/Q _34607_/Q _16935_/X _16936_/X VGND VGND VPWR
+ VPWR _17256_/X sky130_fd_sc_hd__mux4_1
X_16207_ _34258_/Q _34194_/Q _34130_/Q _34066_/Q _16005_/X _16007_/X VGND VGND VPWR
+ VPWR _16207_/X sky130_fd_sc_hd__mux4_1
X_35041_ _35807_/CLK _35041_/D VGND VGND VPWR VPWR _35041_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_155_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _35337_/CLK sky130_fd_sc_hd__clkbuf_16
X_32253_ _34046_/CLK _32253_/D VGND VGND VPWR VPWR _32253_/Q sky130_fd_sc_hd__dfxtp_1
X_17187_ _35309_/Q _35245_/Q _35181_/Q _32301_/Q _17006_/X _17007_/X VGND VGND VPWR
+ VPWR _17187_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16138_ _17903_/A VGND VGND VPWR VPWR _16138_/X sky130_fd_sc_hd__buf_6
X_31204_ _31273_/S VGND VGND VPWR VPWR _31223_/S sky130_fd_sc_hd__buf_4
X_32184_ _35808_/CLK _32184_/D VGND VGND VPWR VPWR _32184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31135_ _31135_/A VGND VGND VPWR VPWR _35787_/D sky130_fd_sc_hd__clkbuf_1
X_16069_ _16056_/X _16061_/X _16066_/X _16068_/X VGND VGND VPWR VPWR _16069_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_931 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35943_ _35943_/CLK _35943_/D VGND VGND VPWR VPWR _35943_/Q sky130_fd_sc_hd__dfxtp_1
X_31066_ _31066_/A VGND VGND VPWR VPWR _35754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30017_ _30017_/A VGND VGND VPWR VPWR _35257_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19828_ _32503_/Q _32375_/Q _32055_/Q _36023_/Q _19576_/X _19717_/X VGND VGND VPWR
+ VPWR _19828_/X sky130_fd_sc_hd__mux4_1
X_35874_ _35938_/CLK _35874_/D VGND VGND VPWR VPWR _35874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34825_ _35848_/CLK _34825_/D VGND VGND VPWR VPWR _34825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19759_ _19647_/X _19757_/X _19758_/X _19650_/X VGND VGND VPWR VPWR _19759_/X sky130_fd_sc_hd__a22o_1
XFILLER_204_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34756_ _35332_/CLK _34756_/D VGND VGND VPWR VPWR _34756_/Q sky130_fd_sc_hd__dfxtp_1
X_22770_ _35786_/Q _35146_/Q _34506_/Q _33866_/Q _20708_/X _20709_/X VGND VGND VPWR
+ VPWR _22770_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31968_ _34970_/CLK _31968_/D VGND VGND VPWR VPWR _31968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33707_ _35320_/CLK _33707_/D VGND VGND VPWR VPWR _33707_/Q sky130_fd_sc_hd__dfxtp_1
X_21721_ _34284_/Q _34220_/Q _34156_/Q _34092_/Q _21689_/X _21690_/X VGND VGND VPWR
+ VPWR _21721_/X sky130_fd_sc_hd__mux4_1
XFILLER_92_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30919_ _30919_/A VGND VGND VPWR VPWR _35684_/D sky130_fd_sc_hd__clkbuf_1
X_34687_ _35837_/CLK _34687_/D VGND VGND VPWR VPWR _34687_/Q sky130_fd_sc_hd__dfxtp_1
X_31899_ _31899_/A VGND VGND VPWR VPWR _36149_/D sky130_fd_sc_hd__clkbuf_1
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24440_ input60/X VGND VGND VPWR VPWR _24440_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_244_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33638_ _33702_/CLK _33638_/D VGND VGND VPWR VPWR _33638_/Q sky130_fd_sc_hd__dfxtp_1
X_21652_ _34026_/Q _33962_/Q _33898_/Q _32234_/Q _21620_/X _21621_/X VGND VGND VPWR
+ VPWR _21652_/X sky130_fd_sc_hd__mux4_1
XFILLER_244_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20603_ _22511_/A VGND VGND VPWR VPWR _20603_/X sky130_fd_sc_hd__buf_4
X_24371_ _32694_/Q _24369_/X _24398_/S VGND VGND VPWR VPWR _24372_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33569_ _34145_/CLK _33569_/D VGND VGND VPWR VPWR _33569_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_394_CLK clkbuf_6_34__f_CLK/X VGND VGND VPWR VPWR _35822_/CLK sky130_fd_sc_hd__clkbuf_16
X_21583_ _21449_/X _21581_/X _21582_/X _21452_/X VGND VGND VPWR VPWR _21583_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26110_ _26110_/A VGND VGND VPWR VPWR _33469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23322_ input52/X VGND VGND VPWR VPWR _23322_/X sky130_fd_sc_hd__buf_4
XFILLER_14_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35308_ _35308_/CLK _35308_/D VGND VGND VPWR VPWR _35308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20534_ _18297_/X _20532_/X _20533_/X _18303_/X VGND VGND VPWR VPWR _20534_/X sky130_fd_sc_hd__a22o_1
X_27090_ _26922_/X _33902_/Q _27104_/S VGND VGND VPWR VPWR _27091_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_1450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26041_ _26041_/A VGND VGND VPWR VPWR _33436_/D sky130_fd_sc_hd__clkbuf_1
X_23253_ input29/X VGND VGND VPWR VPWR _23253_/X sky130_fd_sc_hd__clkbuf_4
X_35239_ _35239_/CLK _35239_/D VGND VGND VPWR VPWR _35239_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_146_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _35341_/CLK sky130_fd_sc_hd__clkbuf_16
X_20465_ _32522_/Q _32394_/Q _32074_/Q _36042_/Q _20282_/X _19307_/A VGND VGND VPWR
+ VPWR _20465_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22204_ _22557_/A VGND VGND VPWR VPWR _22204_/X sky130_fd_sc_hd__buf_4
XFILLER_3_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23184_ _23346_/S VGND VGND VPWR VPWR _23206_/S sky130_fd_sc_hd__clkbuf_8
X_20396_ _34312_/Q _34248_/Q _34184_/Q _34120_/Q _20095_/X _20096_/X VGND VGND VPWR
+ VPWR _20396_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29800_ _29800_/A VGND VGND VPWR VPWR _35154_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22135_ _35575_/Q _35511_/Q _35447_/Q _35383_/Q _21850_/X _21851_/X VGND VGND VPWR
+ VPWR _22135_/X sky130_fd_sc_hd__mux4_1
XTAP_6604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput260 _32126_/Q VGND VGND VPWR VPWR D3[48] sky130_fd_sc_hd__buf_2
X_27992_ _27992_/A VGND VGND VPWR VPWR _34328_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput271 _32136_/Q VGND VGND VPWR VPWR D3[58] sky130_fd_sc_hd__buf_2
XTAP_6637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29731_ _35122_/Q _29163_/X _29737_/S VGND VGND VPWR VPWR _29732_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22066_ _21749_/X _22064_/X _22065_/X _21752_/X VGND VGND VPWR VPWR _22066_/X sky130_fd_sc_hd__a22o_1
X_26943_ input33/X VGND VGND VPWR VPWR _26943_/X sky130_fd_sc_hd__clkbuf_4
XTAP_6659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21017_ _22395_/A VGND VGND VPWR VPWR _21017_/X sky130_fd_sc_hd__buf_4
XFILLER_43_1137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29662_ _35089_/Q _29061_/X _29674_/S VGND VGND VPWR VPWR _29663_/A sky130_fd_sc_hd__mux2_1
X_26874_ _26874_/A VGND VGND VPWR VPWR _33822_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28613_ _28613_/A VGND VGND VPWR VPWR _34623_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25825_ _25115_/X _33334_/Q _25843_/S VGND VGND VPWR VPWR _25826_/A sky130_fd_sc_hd__mux2_1
X_29593_ _29593_/A VGND VGND VPWR VPWR _35056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25756_ _25756_/A VGND VGND VPWR VPWR _33301_/D sky130_fd_sc_hd__clkbuf_1
X_28544_ _28544_/A VGND VGND VPWR VPWR _34590_/D sky130_fd_sc_hd__clkbuf_1
X_22968_ _22968_/A VGND VGND VPWR VPWR _32042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24707_ _23062_/X _32841_/Q _24707_/S VGND VGND VPWR VPWR _24708_/A sky130_fd_sc_hd__mux2_1
X_21919_ _33201_/Q _32561_/Q _35953_/Q _35889_/Q _21674_/X _21675_/X VGND VGND VPWR
+ VPWR _21919_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25687_ _25735_/S VGND VGND VPWR VPWR _25706_/S sky130_fd_sc_hd__buf_4
X_28475_ _26971_/X _34558_/Q _28477_/S VGND VGND VPWR VPWR _28476_/A sky130_fd_sc_hd__mux2_1
X_22899_ _22898_/X _32020_/Q _22908_/S VGND VGND VPWR VPWR _22900_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27426_ _27426_/A _30735_/B VGND VGND VPWR VPWR _27559_/S sky130_fd_sc_hd__nand2_8
X_24638_ _22960_/X _32808_/Q _24644_/S VGND VGND VPWR VPWR _24639_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24569_ _23062_/X _32777_/Q _24569_/S VGND VGND VPWR VPWR _24570_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_385_CLK clkbuf_6_41__f_CLK/X VGND VGND VPWR VPWR _35954_/CLK sky130_fd_sc_hd__clkbuf_16
X_27357_ _27357_/A VGND VGND VPWR VPWR _34028_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17110_ _17106_/X _17109_/X _16794_/X VGND VGND VPWR VPWR _17118_/C sky130_fd_sc_hd__o21ba_1
X_18090_ _35079_/Q _35015_/Q _34951_/Q _34887_/Q _17862_/X _17863_/X VGND VGND VPWR
+ VPWR _18090_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26308_ _25032_/X _33563_/Q _26320_/S VGND VGND VPWR VPWR _26309_/A sky130_fd_sc_hd__mux2_1
X_27288_ _27288_/A VGND VGND VPWR VPWR _33996_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17041_ _16796_/X _17039_/X _17040_/X _16799_/X VGND VGND VPWR VPWR _17041_/X sky130_fd_sc_hd__a22o_1
X_29027_ _29027_/A VGND VGND VPWR VPWR _34819_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_239_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26239_ _26239_/A VGND VGND VPWR VPWR _33530_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_137_CLK clkbuf_6_22__f_CLK/X VGND VGND VPWR VPWR _35791_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_144_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18992_ _18988_/X _18991_/X _18755_/X VGND VGND VPWR VPWR _18993_/D sky130_fd_sc_hd__o21ba_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _34051_/Q _33987_/Q _33923_/Q _32259_/Q _17726_/X _17727_/X VGND VGND VPWR
+ VPWR _17943_/X sky130_fd_sc_hd__mux4_1
X_29929_ _29929_/A VGND VGND VPWR VPWR _35215_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_1215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32940_ _36080_/CLK _32940_/D VGND VGND VPWR VPWR _32940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1075 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17874_ _33537_/Q _33473_/Q _33409_/Q _33345_/Q _17829_/X _17830_/X VGND VGND VPWR
+ VPWR _17874_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19613_ _20095_/A VGND VGND VPWR VPWR _19613_/X sky130_fd_sc_hd__buf_6
X_16825_ _16821_/X _16824_/X _16783_/X _16784_/X VGND VGND VPWR VPWR _16840_/B sky130_fd_sc_hd__o211a_1
X_32871_ _36007_/CLK _32871_/D VGND VGND VPWR VPWR _32871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34610_ _34932_/CLK _34610_/D VGND VGND VPWR VPWR _34610_/Q sky130_fd_sc_hd__dfxtp_1
X_31822_ _31822_/A VGND VGND VPWR VPWR _36112_/D sky130_fd_sc_hd__clkbuf_1
X_19544_ _33007_/Q _32943_/Q _32879_/Q _32815_/Q _19289_/X _19290_/X VGND VGND VPWR
+ VPWR _19544_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35590_ _35590_/CLK _35590_/D VGND VGND VPWR VPWR _35590_/Q sky130_fd_sc_hd__dfxtp_1
X_16756_ _16646_/X _16754_/X _16755_/X _16649_/X VGND VGND VPWR VPWR _16756_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34541_ _35307_/CLK _34541_/D VGND VGND VPWR VPWR _34541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31753_ _36080_/Q input28/X _31763_/S VGND VGND VPWR VPWR _31754_/A sky130_fd_sc_hd__mux2_1
X_19475_ _32493_/Q _32365_/Q _32045_/Q _36013_/Q _19223_/X _19364_/X VGND VGND VPWR
+ VPWR _19475_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16687_ _35295_/Q _35231_/Q _35167_/Q _32287_/Q _16653_/X _16654_/X VGND VGND VPWR
+ VPWR _16687_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18426_ _18422_/X _18425_/X _18371_/X VGND VGND VPWR VPWR _18434_/C sky130_fd_sc_hd__o21ba_1
XFILLER_185_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30704_ _35583_/Q _29203_/X _30704_/S VGND VGND VPWR VPWR _30705_/A sky130_fd_sc_hd__mux2_1
X_34472_ _35879_/CLK _34472_/D VGND VGND VPWR VPWR _34472_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31684_ _36047_/Q input12/X _31700_/S VGND VGND VPWR VPWR _31685_/A sky130_fd_sc_hd__mux2_1
X_36211_ _36211_/CLK _36211_/D VGND VGND VPWR VPWR _36211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33423_ _33490_/CLK _33423_/D VGND VGND VPWR VPWR _33423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18357_ _18357_/A VGND VGND VPWR VPWR _20146_/A sky130_fd_sc_hd__buf_12
X_30635_ _35550_/Q _29101_/X _30641_/S VGND VGND VPWR VPWR _30636_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_376_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _36077_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36142_ _36146_/CLK _36142_/D VGND VGND VPWR VPWR _36142_/Q sky130_fd_sc_hd__dfxtp_1
X_17308_ _17055_/X _17306_/X _17307_/X _17061_/X VGND VGND VPWR VPWR _17308_/X sky130_fd_sc_hd__a22o_1
X_33354_ _33548_/CLK _33354_/D VGND VGND VPWR VPWR _33354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18288_ _18357_/A VGND VGND VPWR VPWR _20095_/A sky130_fd_sc_hd__buf_12
X_30566_ _30566_/A VGND VGND VPWR VPWR _35517_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_8__f_CLK clkbuf_5_4_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_8__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_163_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32305_ _35052_/CLK _32305_/D VGND VGND VPWR VPWR _32305_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_128_CLK clkbuf_6_23__f_CLK/X VGND VGND VPWR VPWR _33685_/CLK sky130_fd_sc_hd__clkbuf_16
X_17239_ _17235_/X _17238_/X _17128_/X VGND VGND VPWR VPWR _17263_/A sky130_fd_sc_hd__o21ba_1
X_36073_ _36137_/CLK _36073_/D VGND VGND VPWR VPWR _36073_/Q sky130_fd_sc_hd__dfxtp_1
X_33285_ _33922_/CLK _33285_/D VGND VGND VPWR VPWR _33285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30497_ _30497_/A VGND VGND VPWR VPWR _35484_/D sky130_fd_sc_hd__clkbuf_1
X_35024_ _35282_/CLK _35024_/D VGND VGND VPWR VPWR _35024_/Q sky130_fd_sc_hd__dfxtp_1
X_20250_ _33027_/Q _32963_/Q _32899_/Q _32835_/Q _19995_/X _19996_/X VGND VGND VPWR
+ VPWR _20250_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32236_ _36018_/CLK _32236_/D VGND VGND VPWR VPWR _32236_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_196_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20181_ _32513_/Q _32385_/Q _32065_/Q _36033_/Q _19929_/X _20070_/X VGND VGND VPWR
+ VPWR _20181_/X sky130_fd_sc_hd__mux4_1
X_32167_ _35666_/CLK _32167_/D VGND VGND VPWR VPWR _32167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31118_ _35779_/Q _29216_/X _31130_/S VGND VGND VPWR VPWR _31119_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32098_ _35808_/CLK _32098_/D VGND VGND VPWR VPWR _32098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23940_ _23940_/A VGND VGND VPWR VPWR _32510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_233_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35926_ _36117_/CLK _35926_/D VGND VGND VPWR VPWR _35926_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_300_CLK clkbuf_6_50__f_CLK/X VGND VGND VPWR VPWR _35963_/CLK sky130_fd_sc_hd__clkbuf_16
X_31049_ _35746_/Q _29113_/X _31067_/S VGND VGND VPWR VPWR _31050_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35857_ _35921_/CLK _35857_/D VGND VGND VPWR VPWR _35857_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23871_ _23871_/A VGND VGND VPWR VPWR _32477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25610_ _33233_/Q _24255_/X _25622_/S VGND VGND VPWR VPWR _25611_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22822_ _32780_/Q _32716_/Q _32652_/Q _36108_/Q _22578_/X _21473_/A VGND VGND VPWR
+ VPWR _22822_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34808_ _34809_/CLK _34808_/D VGND VGND VPWR VPWR _34808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26590_ _26590_/A VGND VGND VPWR VPWR _33696_/D sky130_fd_sc_hd__clkbuf_1
X_35788_ _35788_/CLK _35788_/D VGND VGND VPWR VPWR _35788_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_808 _22904_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_819 _22991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25541_ _33202_/Q _24357_/X _25547_/S VGND VGND VPWR VPWR _25542_/A sky130_fd_sc_hd__mux2_1
X_22753_ _22753_/A _22753_/B _22753_/C _22753_/D VGND VGND VPWR VPWR _22754_/A sky130_fd_sc_hd__or4_4
X_34739_ _34739_/CLK _34739_/D VGND VGND VPWR VPWR _34739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21704_ _35819_/Q _32196_/Q _35691_/Q _35627_/Q _21560_/X _21561_/X VGND VGND VPWR
+ VPWR _21704_/X sky130_fd_sc_hd__mux4_1
X_28260_ _28371_/S VGND VGND VPWR VPWR _28279_/S sky130_fd_sc_hd__buf_4
X_25472_ _33169_/Q _24255_/X _25484_/S VGND VGND VPWR VPWR _25473_/A sky130_fd_sc_hd__mux2_1
X_22684_ _20597_/X _22682_/X _22683_/X _20603_/X VGND VGND VPWR VPWR _22684_/X sky130_fd_sc_hd__a22o_1
XFILLER_201_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24423_ _32711_/Q _24422_/X _24429_/S VGND VGND VPWR VPWR _24424_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27211_ _27211_/A VGND VGND VPWR VPWR _33959_/D sky130_fd_sc_hd__clkbuf_1
X_28191_ _26950_/X _34423_/Q _28207_/S VGND VGND VPWR VPWR _28192_/A sky130_fd_sc_hd__mux2_1
X_21635_ _35561_/Q _35497_/Q _35433_/Q _35369_/Q _21497_/X _21498_/X VGND VGND VPWR
+ VPWR _21635_/X sky130_fd_sc_hd__mux4_1
XFILLER_233_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_367_CLK clkbuf_6_42__f_CLK/X VGND VGND VPWR VPWR _36146_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27142_ _26999_/X _33927_/Q _27146_/S VGND VGND VPWR VPWR _27143_/A sky130_fd_sc_hd__mux2_1
X_24354_ input29/X VGND VGND VPWR VPWR _24354_/X sky130_fd_sc_hd__buf_4
XFILLER_51_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21566_ _33191_/Q _32551_/Q _35943_/Q _35879_/Q _21321_/X _21322_/X VGND VGND VPWR
+ VPWR _21566_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23305_ _32219_/Q _23303_/X _23334_/S VGND VGND VPWR VPWR _23306_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_119_CLK clkbuf_6_21__f_CLK/X VGND VGND VPWR VPWR _34001_/CLK sky130_fd_sc_hd__clkbuf_16
X_20517_ _18314_/X _20515_/X _20516_/X _18323_/X VGND VGND VPWR VPWR _20517_/X sky130_fd_sc_hd__a22o_1
XFILLER_126_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27073_ _26897_/X _33894_/Q _27083_/S VGND VGND VPWR VPWR _27074_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24285_ _24285_/A VGND VGND VPWR VPWR _32666_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21497_ _22556_/A VGND VGND VPWR VPWR _21497_/X sky130_fd_sc_hd__buf_4
XFILLER_165_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26024_ _26024_/A VGND VGND VPWR VPWR _33428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23236_ _23236_/A VGND VGND VPWR VPWR _32196_/D sky130_fd_sc_hd__clkbuf_1
X_20448_ _20155_/X _20446_/X _20447_/X _20158_/X VGND VGND VPWR VPWR _20448_/X sky130_fd_sc_hd__a22o_1
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23167_ _32167_/Q _23096_/X _23182_/S VGND VGND VPWR VPWR _23168_/A sky130_fd_sc_hd__mux2_1
XTAP_7146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20379_ _35847_/Q _32227_/Q _35719_/Q _35655_/Q _18289_/X _18291_/X VGND VGND VPWR
+ VPWR _20379_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1207 _23142_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22118_ _33783_/Q _33719_/Q _33655_/Q _33591_/Q _21796_/X _21797_/X VGND VGND VPWR
+ VPWR _22118_/X sky130_fd_sc_hd__mux4_1
XTAP_6434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1218 _24264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1229 _24416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23098_ _23098_/A VGND VGND VPWR VPWR _32145_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27975_ _27975_/A VGND VGND VPWR VPWR _34320_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29714_ _35114_/Q _29138_/X _29716_/S VGND VGND VPWR VPWR _29715_/A sky130_fd_sc_hd__mux2_1
XTAP_6478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26926_ _26925_/X _33839_/Q _26944_/S VGND VGND VPWR VPWR _26927_/A sky130_fd_sc_hd__mux2_1
X_22049_ _22045_/X _22048_/X _21728_/X VGND VGND VPWR VPWR _22071_/A sky130_fd_sc_hd__o21ba_1
XFILLER_94_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29645_ _29645_/A VGND VGND VPWR VPWR _35081_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26857_ input3/X VGND VGND VPWR VPWR _26857_/X sky130_fd_sc_hd__buf_4
XTAP_5799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16610_ _35741_/Q _35101_/Q _34461_/Q _33821_/Q _16434_/X _16435_/X VGND VGND VPWR
+ VPWR _16610_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25808_ _25091_/X _33326_/Q _25822_/S VGND VGND VPWR VPWR _25809_/A sky130_fd_sc_hd__mux2_1
X_17590_ _34041_/Q _33977_/Q _33913_/Q _32249_/Q _17373_/X _17374_/X VGND VGND VPWR
+ VPWR _17590_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29576_ _29576_/A VGND VGND VPWR VPWR _35048_/D sky130_fd_sc_hd__clkbuf_1
X_26788_ _33790_/Q _24394_/X _26790_/S VGND VGND VPWR VPWR _26789_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28527_ _28527_/A VGND VGND VPWR VPWR _34582_/D sky130_fd_sc_hd__clkbuf_1
X_16541_ _35803_/Q _32178_/Q _35675_/Q _35611_/Q _16254_/X _16255_/X VGND VGND VPWR
+ VPWR _16541_/X sky130_fd_sc_hd__mux4_1
X_25739_ _27968_/A _26685_/B VGND VGND VPWR VPWR _25872_/S sky130_fd_sc_hd__nand2_8
XFILLER_56_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19260_ _20095_/A VGND VGND VPWR VPWR _19260_/X sky130_fd_sc_hd__buf_4
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28458_ _28506_/S VGND VGND VPWR VPWR _28477_/S sky130_fd_sc_hd__buf_4
X_16472_ _16468_/X _16471_/X _16430_/X _16431_/X VGND VGND VPWR VPWR _16487_/B sky130_fd_sc_hd__o211a_2
XFILLER_108_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18211_ _16056_/X _18209_/X _18210_/X _16068_/X VGND VGND VPWR VPWR _18211_/X sky130_fd_sc_hd__a22o_1
X_27409_ _27409_/A VGND VGND VPWR VPWR _34053_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_358_CLK clkbuf_6_43__f_CLK/X VGND VGND VPWR VPWR _34222_/CLK sky130_fd_sc_hd__clkbuf_16
X_19191_ _32997_/Q _32933_/Q _32869_/Q _32805_/Q _18936_/X _18937_/X VGND VGND VPWR
+ VPWR _19191_/X sky130_fd_sc_hd__mux4_1
X_28389_ _26844_/X _34517_/Q _28393_/S VGND VGND VPWR VPWR _28390_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18142_ _35593_/Q _35529_/Q _35465_/Q _35401_/Q _17956_/X _17957_/X VGND VGND VPWR
+ VPWR _18142_/X sky130_fd_sc_hd__mux4_1
X_30420_ _23277_/X _35448_/Q _30434_/S VGND VGND VPWR VPWR _30421_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_917 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18073_ _33287_/Q _36167_/Q _33159_/Q _33095_/Q _17764_/X _17765_/X VGND VGND VPWR
+ VPWR _18073_/X sky130_fd_sc_hd__mux4_1
X_30351_ _30351_/A VGND VGND VPWR VPWR _35415_/D sky130_fd_sc_hd__clkbuf_1
X_17024_ _17018_/X _17023_/X _16775_/X VGND VGND VPWR VPWR _17046_/A sky130_fd_sc_hd__o21ba_1
X_33070_ _36081_/CLK _33070_/D VGND VGND VPWR VPWR _33070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30282_ _35383_/Q _29179_/X _30298_/S VGND VGND VPWR VPWR _30283_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32021_ _36052_/CLK _32021_/D VGND VGND VPWR VPWR _32021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18975_ _32479_/Q _32351_/Q _32031_/Q _35999_/Q _18870_/X _18658_/X VGND VGND VPWR
+ VPWR _18975_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ _17705_/X _17924_/X _17925_/X _17708_/X VGND VGND VPWR VPWR _17926_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33972_ _34228_/CLK _33972_/D VGND VGND VPWR VPWR _33972_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35711_ _35711_/CLK _35711_/D VGND VGND VPWR VPWR _35711_/Q sky130_fd_sc_hd__dfxtp_1
X_32923_ _36118_/CLK _32923_/D VGND VGND VPWR VPWR _32923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17857_ _35328_/Q _35264_/Q _35200_/Q _32320_/Q _17712_/X _17713_/X VGND VGND VPWR
+ VPWR _17857_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35642_ _35834_/CLK _35642_/D VGND VGND VPWR VPWR _35642_/Q sky130_fd_sc_hd__dfxtp_1
X_16808_ _17867_/A VGND VGND VPWR VPWR _16808_/X sky130_fd_sc_hd__buf_2
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32854_ _36116_/CLK _32854_/D VGND VGND VPWR VPWR _32854_/Q sky130_fd_sc_hd__dfxtp_1
X_17788_ _34558_/Q _32446_/Q _34430_/Q _34366_/Q _17578_/X _17579_/X VGND VGND VPWR
+ VPWR _17788_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31805_ _36105_/Q input55/X _31805_/S VGND VGND VPWR VPWR _31806_/A sky130_fd_sc_hd__mux2_1
X_19527_ _34542_/Q _32430_/Q _34414_/Q _34350_/Q _19525_/X _19526_/X VGND VGND VPWR
+ VPWR _19527_/X sky130_fd_sc_hd__mux4_1
XFILLER_223_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35573_ _36021_/CLK _35573_/D VGND VGND VPWR VPWR _35573_/Q sky130_fd_sc_hd__dfxtp_1
X_16739_ _16489_/X _16735_/X _16738_/X _16494_/X VGND VGND VPWR VPWR _16739_/X sky130_fd_sc_hd__a22o_1
XFILLER_235_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32785_ _35982_/CLK _32785_/D VGND VGND VPWR VPWR _32785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34524_ _35166_/CLK _34524_/D VGND VGND VPWR VPWR _34524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19458_ _35052_/Q _34988_/Q _34924_/Q _34860_/Q _19456_/X _19457_/X VGND VGND VPWR
+ VPWR _19458_/X sky130_fd_sc_hd__mux4_1
X_31736_ _36072_/Q input19/X _31742_/S VGND VGND VPWR VPWR _31737_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18409_ _20147_/A VGND VGND VPWR VPWR _18409_/X sky130_fd_sc_hd__buf_4
XFILLER_22_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34455_ _35667_/CLK _34455_/D VGND VGND VPWR VPWR _34455_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_349_CLK clkbuf_6_46__f_CLK/X VGND VGND VPWR VPWR _34227_/CLK sky130_fd_sc_hd__clkbuf_16
X_31667_ _31667_/A VGND VGND VPWR VPWR _36039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19389_ _20256_/A VGND VGND VPWR VPWR _19389_/X sky130_fd_sc_hd__buf_6
XFILLER_241_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33406_ _34302_/CLK _33406_/D VGND VGND VPWR VPWR _33406_/Q sky130_fd_sc_hd__dfxtp_1
X_21420_ _33251_/Q _36131_/Q _33123_/Q _33059_/Q _21305_/X _21306_/X VGND VGND VPWR
+ VPWR _21420_/X sky130_fd_sc_hd__mux4_1
X_30618_ _35542_/Q _29076_/X _30620_/S VGND VGND VPWR VPWR _30619_/A sky130_fd_sc_hd__mux2_1
X_34386_ _35028_/CLK _34386_/D VGND VGND VPWR VPWR _34386_/Q sky130_fd_sc_hd__dfxtp_1
X_31598_ _31598_/A VGND VGND VPWR VPWR _36006_/D sky130_fd_sc_hd__clkbuf_1
X_36125_ _36125_/CLK _36125_/D VGND VGND VPWR VPWR _36125_/Q sky130_fd_sc_hd__dfxtp_1
X_33337_ _34298_/CLK _33337_/D VGND VGND VPWR VPWR _33337_/Q sky130_fd_sc_hd__dfxtp_1
X_21351_ _35809_/Q _32185_/Q _35681_/Q _35617_/Q _21207_/X _21208_/X VGND VGND VPWR
+ VPWR _21351_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30549_ _30549_/A VGND VGND VPWR VPWR _35509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20302_ _20298_/X _20301_/X _20167_/X VGND VGND VPWR VPWR _20303_/D sky130_fd_sc_hd__o21ba_1
XFILLER_50_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24070_ _24070_/A VGND VGND VPWR VPWR _32571_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36056_ _36123_/CLK _36056_/D VGND VGND VPWR VPWR _36056_/Q sky130_fd_sc_hd__dfxtp_1
X_21282_ _35551_/Q _35487_/Q _35423_/Q _35359_/Q _21144_/X _21145_/X VGND VGND VPWR
+ VPWR _21282_/X sky130_fd_sc_hd__mux4_1
X_33268_ _34229_/CLK _33268_/D VGND VGND VPWR VPWR _33268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35007_ _35989_/CLK _35007_/D VGND VGND VPWR VPWR _35007_/Q sky130_fd_sc_hd__dfxtp_1
X_23021_ _23021_/A VGND VGND VPWR VPWR _32059_/D sky130_fd_sc_hd__clkbuf_1
X_20233_ _34562_/Q _32450_/Q _34434_/Q _34370_/Q _20231_/X _20232_/X VGND VGND VPWR
+ VPWR _20233_/X sky130_fd_sc_hd__mux4_1
X_32219_ _35715_/CLK _32219_/D VGND VGND VPWR VPWR _32219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33199_ _35952_/CLK _33199_/D VGND VGND VPWR VPWR _33199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20164_ _35072_/Q _35008_/Q _34944_/Q _34880_/Q _20162_/X _20163_/X VGND VGND VPWR
+ VPWR _20164_/X sky130_fd_sc_hd__mux4_1
XTAP_5007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27760_ _34219_/Q _24335_/X _27760_/S VGND VGND VPWR VPWR _27761_/A sky130_fd_sc_hd__mux2_1
X_20095_ _20095_/A VGND VGND VPWR VPWR _20095_/X sky130_fd_sc_hd__buf_6
X_24972_ _24972_/A VGND VGND VPWR VPWR _32965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26711_ _33753_/Q _24280_/X _26727_/S VGND VGND VPWR VPWR _26712_/A sky130_fd_sc_hd__mux2_1
X_35909_ _35909_/CLK _35909_/D VGND VGND VPWR VPWR _35909_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23923_ _23003_/X _32502_/Q _23941_/S VGND VGND VPWR VPWR _23924_/A sky130_fd_sc_hd__mux2_1
X_27691_ _27691_/A VGND VGND VPWR VPWR _34186_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29430_ _23152_/X _34979_/Q _29446_/S VGND VGND VPWR VPWR _29431_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23854_ _23854_/A VGND VGND VPWR VPWR _32469_/D sky130_fd_sc_hd__clkbuf_1
X_26642_ _25125_/X _33721_/Q _26654_/S VGND VGND VPWR VPWR _26643_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_605 _18435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_616 _18505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22805_ _22801_/X _22804_/X _22453_/A VGND VGND VPWR VPWR _22813_/C sky130_fd_sc_hd__o21ba_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29361_ _29361_/A VGND VGND VPWR VPWR _34946_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_627 _18712_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26573_ _25022_/X _33688_/Q _26591_/S VGND VGND VPWR VPWR _26574_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_638 _19245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23785_ _23785_/A VGND VGND VPWR VPWR _32437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1041 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_649 _20202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20997_ _20993_/X _20996_/X _20640_/X _20642_/X VGND VGND VPWR VPWR _21012_/B sky130_fd_sc_hd__o211a_1
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28312_ _28312_/A VGND VGND VPWR VPWR _34480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22736_ _33033_/Q _32969_/Q _32905_/Q _32841_/Q _20580_/X _20583_/X VGND VGND VPWR
+ VPWR _22736_/X sky130_fd_sc_hd__mux4_1
X_25524_ _33194_/Q _24332_/X _25526_/S VGND VGND VPWR VPWR _25525_/A sky130_fd_sc_hd__mux2_1
X_29292_ _29382_/S VGND VGND VPWR VPWR _29311_/S sky130_fd_sc_hd__buf_4
XFILLER_81_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28243_ _28243_/A VGND VGND VPWR VPWR _34447_/D sky130_fd_sc_hd__clkbuf_1
X_25455_ _25455_/A VGND VGND VPWR VPWR _33163_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22667_ _22501_/X _22665_/X _22666_/X _22506_/X VGND VGND VPWR VPWR _22667_/X sky130_fd_sc_hd__a22o_1
XFILLER_71_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24406_ _24406_/A VGND VGND VPWR VPWR _32705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21618_ _21442_/X _21616_/X _21617_/X _21447_/X VGND VGND VPWR VPWR _21618_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28174_ _26925_/X _34415_/Q _28186_/S VGND VGND VPWR VPWR _28175_/A sky130_fd_sc_hd__mux2_1
X_25386_ _25386_/A VGND VGND VPWR VPWR _33130_/D sky130_fd_sc_hd__clkbuf_1
X_22598_ _22455_/X _22596_/X _22597_/X _22458_/X VGND VGND VPWR VPWR _22598_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27125_ _26974_/X _33919_/Q _27125_/S VGND VGND VPWR VPWR _27126_/A sky130_fd_sc_hd__mux2_1
X_24337_ _24337_/A VGND VGND VPWR VPWR _32683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21549_ _33511_/Q _33447_/Q _33383_/Q _33319_/Q _21370_/X _21371_/X VGND VGND VPWR
+ VPWR _21549_/X sky130_fd_sc_hd__mux4_1
XFILLER_126_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1080 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27056_ _26872_/X _33886_/Q _27062_/S VGND VGND VPWR VPWR _27057_/A sky130_fd_sc_hd__mux2_1
X_24268_ _32661_/Q _24267_/X _24274_/S VGND VGND VPWR VPWR _24269_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26007_ _25186_/X _33421_/Q _26007_/S VGND VGND VPWR VPWR _26008_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23219_ _23219_/A VGND VGND VPWR VPWR _32190_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_1083 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24199_ _23010_/X _32632_/Q _24213_/S VGND VGND VPWR VPWR _24200_/A sky130_fd_sc_hd__mux2_1
XTAP_6220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1004 _17901_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1015 _17995_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1026 _17865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1037 _17152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1048 _17867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18760_ _34265_/Q _34201_/Q _34137_/Q _34073_/Q _18683_/X _18684_/X VGND VGND VPWR
+ VPWR _18760_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27958_ _34313_/Q _24428_/X _27958_/S VGND VGND VPWR VPWR _27959_/A sky130_fd_sc_hd__mux2_1
XTAP_5530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1059 _16592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17711_ _34812_/Q _34748_/Q _34684_/Q _34620_/Q _17641_/X _17642_/X VGND VGND VPWR
+ VPWR _17711_/X sky130_fd_sc_hd__mux4_1
XTAP_5563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26909_ input21/X VGND VGND VPWR VPWR _26909_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18691_ _32727_/Q _32663_/Q _32599_/Q _36055_/Q _18513_/X _18650_/X VGND VGND VPWR
+ VPWR _18691_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_5_18_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_18_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XTAP_5585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27889_ _34280_/Q _24326_/X _27895_/S VGND VGND VPWR VPWR _27890_/A sky130_fd_sc_hd__mux2_1
XTAP_5596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29628_ _35073_/Q _29210_/X _29644_/S VGND VGND VPWR VPWR _29629_/A sky130_fd_sc_hd__mux2_1
X_17642_ _17995_/A VGND VGND VPWR VPWR _17642_/X sky130_fd_sc_hd__buf_6
XTAP_4873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17573_ _17352_/X _17571_/X _17572_/X _17355_/X VGND VGND VPWR VPWR _17573_/X sky130_fd_sc_hd__a22o_1
X_29559_ _29559_/A VGND VGND VPWR VPWR _35040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_232_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19312_ _19101_/X _19310_/X _19311_/X _19106_/X VGND VGND VPWR VPWR _19312_/X sky130_fd_sc_hd__a22o_1
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16524_ _16518_/X _16523_/X _16455_/X VGND VGND VPWR VPWR _16525_/D sky130_fd_sc_hd__o21ba_1
X_32570_ _36027_/CLK _32570_/D VGND VGND VPWR VPWR _32570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31521_ _23310_/X _35970_/Q _31535_/S VGND VGND VPWR VPWR _31522_/A sky130_fd_sc_hd__mux2_1
X_19243_ _19239_/X _19242_/X _19108_/X VGND VGND VPWR VPWR _19244_/D sky130_fd_sc_hd__o21ba_1
XFILLER_108_1248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16455_ _17867_/A VGND VGND VPWR VPWR _16455_/X sky130_fd_sc_hd__buf_2
XFILLER_176_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34240_ _36165_/CLK _34240_/D VGND VGND VPWR VPWR _34240_/Q sky130_fd_sc_hd__dfxtp_1
X_31452_ _31452_/A VGND VGND VPWR VPWR _35937_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19174_ _34532_/Q _32420_/Q _34404_/Q _34340_/Q _19172_/X _19173_/X VGND VGND VPWR
+ VPWR _19174_/X sky130_fd_sc_hd__mux4_1
X_16386_ _16136_/X _16382_/X _16385_/X _16141_/X VGND VGND VPWR VPWR _16386_/X sky130_fd_sc_hd__a22o_1
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18125_ _33801_/Q _33737_/Q _33673_/Q _33609_/Q _17902_/X _17903_/X VGND VGND VPWR
+ VPWR _18125_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30403_ _23250_/X _35440_/Q _30413_/S VGND VGND VPWR VPWR _30404_/A sky130_fd_sc_hd__mux2_1
X_34171_ _34171_/CLK _34171_/D VGND VGND VPWR VPWR _34171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31383_ _31383_/A VGND VGND VPWR VPWR _35904_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33122_ _36130_/CLK _33122_/D VGND VGND VPWR VPWR _33122_/Q sky130_fd_sc_hd__dfxtp_1
X_18056_ _34822_/Q _34758_/Q _34694_/Q _34630_/Q _17994_/X _17995_/X VGND VGND VPWR
+ VPWR _18056_/X sky130_fd_sc_hd__mux4_1
X_30334_ _23090_/X _35407_/Q _30350_/S VGND VGND VPWR VPWR _30335_/A sky130_fd_sc_hd__mux2_1
XANTENNA_1 CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17007_ _17007_/A VGND VGND VPWR VPWR _17007_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33053_ _33244_/CLK _33053_/D VGND VGND VPWR VPWR _33053_/Q sky130_fd_sc_hd__dfxtp_1
X_30265_ _35375_/Q _29154_/X _30277_/S VGND VGND VPWR VPWR _30266_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32004_ _36194_/CLK _32004_/D VGND VGND VPWR VPWR _32004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30196_ _35342_/Q _29048_/X _30214_/S VGND VGND VPWR VPWR _30197_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18958_ _35038_/Q _34974_/Q _34910_/Q _34846_/Q _18750_/X _18751_/X VGND VGND VPWR
+ VPWR _18958_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17909_ _33538_/Q _33474_/Q _33410_/Q _33346_/Q _17829_/X _17830_/X VGND VGND VPWR
+ VPWR _17909_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33955_ _36130_/CLK _33955_/D VGND VGND VPWR VPWR _33955_/Q sky130_fd_sc_hd__dfxtp_1
X_18889_ _18748_/X _18887_/X _18888_/X _18753_/X VGND VGND VPWR VPWR _18889_/X sky130_fd_sc_hd__a22o_1
XFILLER_227_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32906_ _35978_/CLK _32906_/D VGND VGND VPWR VPWR _32906_/Q sky130_fd_sc_hd__dfxtp_1
X_20920_ _33237_/Q _36117_/Q _33109_/Q _33045_/Q _20620_/X _20621_/X VGND VGND VPWR
+ VPWR _20920_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33886_ _36200_/CLK _33886_/D VGND VGND VPWR VPWR _33886_/Q sky130_fd_sc_hd__dfxtp_1
X_32837_ _32965_/CLK _32837_/D VGND VGND VPWR VPWR _32837_/Q sky130_fd_sc_hd__dfxtp_1
X_20851_ _32979_/Q _32915_/Q _32851_/Q _32787_/Q _20633_/X _20635_/X VGND VGND VPWR
+ VPWR _20851_/X sky130_fd_sc_hd__mux4_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35625_ _35815_/CLK _35625_/D VGND VGND VPWR VPWR _35625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23570_ _23570_/A VGND VGND VPWR VPWR _32336_/D sky130_fd_sc_hd__clkbuf_1
X_35556_ _35811_/CLK _35556_/D VGND VGND VPWR VPWR _35556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32768_ _36098_/CLK _32768_/D VGND VGND VPWR VPWR _32768_/Q sky130_fd_sc_hd__dfxtp_1
X_20782_ _33233_/Q _36113_/Q _33105_/Q _33041_/Q _20620_/X _20621_/X VGND VGND VPWR
+ VPWR _20782_/X sky130_fd_sc_hd__mux4_1
XFILLER_126_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34507_ _35787_/CLK _34507_/D VGND VGND VPWR VPWR _34507_/Q sky130_fd_sc_hd__dfxtp_1
X_22521_ _35842_/Q _32221_/Q _35714_/Q _35650_/Q _22266_/X _22267_/X VGND VGND VPWR
+ VPWR _22521_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31719_ _36064_/Q input10/X _31721_/S VGND VGND VPWR VPWR _31720_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35487_ _35744_/CLK _35487_/D VGND VGND VPWR VPWR _35487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32699_ _33083_/CLK _32699_/D VGND VGND VPWR VPWR _32699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25240_ _25240_/A VGND VGND VPWR VPWR _33061_/D sky130_fd_sc_hd__clkbuf_1
X_34438_ _35078_/CLK _34438_/D VGND VGND VPWR VPWR _34438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22452_ _22305_/X _22450_/X _22451_/X _22308_/X VGND VGND VPWR VPWR _22452_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21403_ _22462_/A VGND VGND VPWR VPWR _21403_/X sky130_fd_sc_hd__clkbuf_8
X_25171_ input54/X VGND VGND VPWR VPWR _25171_/X sky130_fd_sc_hd__buf_4
X_34369_ _36038_/CLK _34369_/D VGND VGND VPWR VPWR _34369_/Q sky130_fd_sc_hd__dfxtp_1
X_22383_ _22305_/X _22379_/X _22382_/X _22308_/X VGND VGND VPWR VPWR _22383_/X sky130_fd_sc_hd__a22o_1
XFILLER_202_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36108_ _36109_/CLK _36108_/D VGND VGND VPWR VPWR _36108_/Q sky130_fd_sc_hd__dfxtp_1
X_24122_ _24122_/A VGND VGND VPWR VPWR _32595_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21334_ _21334_/A VGND VGND VPWR VPWR _36192_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36039_ _36039_/CLK _36039_/D VGND VGND VPWR VPWR _36039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28930_ _28930_/A VGND VGND VPWR VPWR _34773_/D sky130_fd_sc_hd__clkbuf_1
X_24053_ _24053_/A VGND VGND VPWR VPWR _32563_/D sky130_fd_sc_hd__clkbuf_1
X_21265_ _21089_/X _21263_/X _21264_/X _21094_/X VGND VGND VPWR VPWR _21265_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_50_CLK clkbuf_leaf_50_CLK/A VGND VGND VPWR VPWR _36130_/CLK sky130_fd_sc_hd__clkbuf_16
X_23004_ _23075_/S VGND VGND VPWR VPWR _23032_/S sky130_fd_sc_hd__buf_4
X_20216_ _20061_/X _20214_/X _20215_/X _20067_/X VGND VGND VPWR VPWR _20216_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28861_ _26943_/X _34741_/Q _28861_/S VGND VGND VPWR VPWR _28862_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21196_ _33501_/Q _33437_/Q _33373_/Q _33309_/Q _21017_/X _21018_/X VGND VGND VPWR
+ VPWR _21196_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27812_ _27812_/A VGND VGND VPWR VPWR _34243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20147_ _20147_/A VGND VGND VPWR VPWR _20147_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_89_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28792_ _26841_/X _34708_/Q _28798_/S VGND VGND VPWR VPWR _28793_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27743_ _27743_/A VGND VGND VPWR VPWR _34210_/D sky130_fd_sc_hd__clkbuf_1
X_20078_ _20000_/X _20076_/X _20077_/X _20003_/X VGND VGND VPWR VPWR _20078_/X sky130_fd_sc_hd__a22o_1
X_24955_ _24955_/A VGND VGND VPWR VPWR _32957_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23906_ _22979_/X _32494_/Q _23920_/S VGND VGND VPWR VPWR _23907_/A sky130_fd_sc_hd__mux2_1
X_27674_ _34178_/Q _24407_/X _27688_/S VGND VGND VPWR VPWR _27675_/A sky130_fd_sc_hd__mux2_1
XTAP_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24886_ _24886_/A VGND VGND VPWR VPWR _32924_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_218_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_402 _36210_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29413_ _23127_/X _34971_/Q _29425_/S VGND VGND VPWR VPWR _29414_/A sky130_fd_sc_hd__mux2_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_413 _36212_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26625_ _25100_/X _33713_/Q _26633_/S VGND VGND VPWR VPWR _26626_/A sky130_fd_sc_hd__mux2_1
X_23837_ _23837_/A VGND VGND VPWR VPWR _23970_/S sky130_fd_sc_hd__buf_12
XTAP_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_424 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_435 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_446 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29344_ _29344_/A VGND VGND VPWR VPWR _34938_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_457 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26556_ _24998_/X _33680_/Q _26570_/S VGND VGND VPWR VPWR _26557_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23768_ _22976_/X _32429_/Q _23784_/S VGND VGND VPWR VPWR _23769_/A sky130_fd_sc_hd__mux2_1
XANTENNA_468 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_479 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25507_ _25597_/S VGND VGND VPWR VPWR _25526_/S sky130_fd_sc_hd__buf_4
X_22719_ _34568_/Q _32456_/Q _34440_/Q _34376_/Q _22531_/X _22532_/X VGND VGND VPWR
+ VPWR _22719_/X sky130_fd_sc_hd__mux4_1
X_29275_ _29275_/A VGND VGND VPWR VPWR _34905_/D sky130_fd_sc_hd__clkbuf_1
X_23699_ _30329_/A _28913_/B VGND VGND VPWR VPWR _28778_/B sky130_fd_sc_hd__nor2_8
XFILLER_198_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26487_ _25097_/X _33648_/Q _26497_/S VGND VGND VPWR VPWR _26488_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28226_ _27002_/X _34440_/Q _28228_/S VGND VGND VPWR VPWR _28227_/A sky130_fd_sc_hd__mux2_1
X_16240_ _33747_/Q _33683_/Q _33619_/Q _33555_/Q _16137_/X _16138_/X VGND VGND VPWR
+ VPWR _16240_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25438_ _25156_/X _33155_/Q _25450_/S VGND VGND VPWR VPWR _25439_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16171_ _16165_/X _16170_/X _16100_/X VGND VGND VPWR VPWR _16172_/D sky130_fd_sc_hd__o21ba_1
X_28157_ _26900_/X _34407_/Q _28165_/S VGND VGND VPWR VPWR _28158_/A sky130_fd_sc_hd__mux2_1
X_25369_ _25053_/X _33122_/Q _25387_/S VGND VGND VPWR VPWR _25370_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27108_ _27108_/A VGND VGND VPWR VPWR _33910_/D sky130_fd_sc_hd__clkbuf_1
X_28088_ _28088_/A VGND VGND VPWR VPWR _34374_/D sky130_fd_sc_hd__clkbuf_1
X_19930_ _32506_/Q _32378_/Q _32058_/Q _36026_/Q _19929_/X _19717_/X VGND VGND VPWR
+ VPWR _19930_/X sky130_fd_sc_hd__mux4_1
X_27039_ _26847_/X _33878_/Q _27041_/S VGND VGND VPWR VPWR _27040_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_41_CLK clkbuf_6_7__f_CLK/X VGND VGND VPWR VPWR _36124_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_107_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30050_ _30050_/A VGND VGND VPWR VPWR _35273_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19861_ _32760_/Q _32696_/Q _32632_/Q _36088_/Q _19572_/X _19709_/X VGND VGND VPWR
+ VPWR _19861_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_1_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_1_0_CLK/X sky130_fd_sc_hd__clkbuf_8
X_18812_ _35546_/Q _35482_/Q _35418_/Q _35354_/Q _18491_/X _18492_/X VGND VGND VPWR
+ VPWR _18812_/X sky130_fd_sc_hd__mux4_1
XTAP_6050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput93 _31962_/Q VGND VGND VPWR VPWR D1[12] sky130_fd_sc_hd__buf_2
XFILLER_7_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19792_ _35830_/Q _32208_/Q _35702_/Q _35638_/Q _19613_/X _19614_/X VGND VGND VPWR
+ VPWR _19792_/X sky130_fd_sc_hd__mux4_1
XTAP_6061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18743_ _19449_/A VGND VGND VPWR VPWR _18743_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33740_ _34124_/CLK _33740_/D VGND VGND VPWR VPWR _33740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18674_ _35286_/Q _35222_/Q _35158_/Q _32278_/Q _18600_/X _18601_/X VGND VGND VPWR
+ VPWR _18674_/X sky130_fd_sc_hd__mux4_1
X_30952_ _30952_/A VGND VGND VPWR VPWR _35700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17625_ _17978_/A VGND VGND VPWR VPWR _17625_/X sky130_fd_sc_hd__buf_6
XTAP_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33671_ _34819_/CLK _33671_/D VGND VGND VPWR VPWR _33671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30883_ _30883_/A VGND VGND VPWR VPWR _35667_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35410_ _35922_/CLK _35410_/D VGND VGND VPWR VPWR _35410_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32622_ _36078_/CLK _32622_/D VGND VGND VPWR VPWR _32622_/Q sky130_fd_sc_hd__dfxtp_1
X_17556_ _33528_/Q _33464_/Q _33400_/Q _33336_/Q _17476_/X _17477_/X VGND VGND VPWR
+ VPWR _17556_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_980 _17855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35341_ _35341_/CLK _35341_/D VGND VGND VPWR VPWR _35341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16507_ _16357_/X _16505_/X _16506_/X _16361_/X VGND VGND VPWR VPWR _16507_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_991 _17860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32553_ _35944_/CLK _32553_/D VGND VGND VPWR VPWR _32553_/Q sky130_fd_sc_hd__dfxtp_1
X_17487_ _33014_/Q _32950_/Q _32886_/Q _32822_/Q _17342_/X _17343_/X VGND VGND VPWR
+ VPWR _17487_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31504_ _23283_/X _35962_/Q _31514_/S VGND VGND VPWR VPWR _31505_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19226_ _19010_/X _19224_/X _19225_/X _19014_/X VGND VGND VPWR VPWR _19226_/X sky130_fd_sc_hd__a22o_1
X_35272_ _35334_/CLK _35272_/D VGND VGND VPWR VPWR _35272_/Q sky130_fd_sc_hd__dfxtp_1
X_16438_ _35544_/Q _35480_/Q _35416_/Q _35352_/Q _16191_/X _16192_/X VGND VGND VPWR
+ VPWR _16438_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32484_ _36005_/CLK _32484_/D VGND VGND VPWR VPWR _32484_/Q sky130_fd_sc_hd__dfxtp_1
X_34223_ _34286_/CLK _34223_/D VGND VGND VPWR VPWR _34223_/Q sky130_fd_sc_hd__dfxtp_1
X_31435_ _23121_/X _35929_/Q _31451_/S VGND VGND VPWR VPWR _31436_/A sky130_fd_sc_hd__mux2_1
X_19157_ _19002_/X _19155_/X _19156_/X _19008_/X VGND VGND VPWR VPWR _19157_/X sky130_fd_sc_hd__a22o_1
X_16369_ _17932_/A VGND VGND VPWR VPWR _16369_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_145_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18108_ _18104_/X _18107_/X _17842_/X _17843_/X VGND VGND VPWR VPWR _18123_/B sky130_fd_sc_hd__o211a_1
X_34154_ _34154_/CLK _34154_/D VGND VGND VPWR VPWR _34154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31366_ _31366_/A VGND VGND VPWR VPWR _35896_/D sky130_fd_sc_hd__clkbuf_1
X_19088_ _20295_/A VGND VGND VPWR VPWR _19088_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_219_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33105_ _36114_/CLK _33105_/D VGND VGND VPWR VPWR _33105_/Q sky130_fd_sc_hd__dfxtp_1
X_18039_ _34054_/Q _33990_/Q _33926_/Q _32262_/Q _17726_/X _17727_/X VGND VGND VPWR
+ VPWR _18039_/X sky130_fd_sc_hd__mux4_1
X_30317_ _35400_/Q _29231_/X _30319_/S VGND VGND VPWR VPWR _30318_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34085_ _34149_/CLK _34085_/D VGND VGND VPWR VPWR _34085_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_32_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _34266_/CLK sky130_fd_sc_hd__clkbuf_16
X_31297_ _31408_/S VGND VGND VPWR VPWR _31316_/S sky130_fd_sc_hd__buf_4
X_33036_ _36045_/CLK _33036_/D VGND VGND VPWR VPWR _33036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21050_ _22462_/A VGND VGND VPWR VPWR _21050_/X sky130_fd_sc_hd__buf_4
XFILLER_67_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30248_ _35367_/Q _29129_/X _30256_/S VGND VGND VPWR VPWR _30249_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20001_ _35836_/Q _32214_/Q _35708_/Q _35644_/Q _19966_/X _19967_/X VGND VGND VPWR
+ VPWR _20001_/X sky130_fd_sc_hd__mux4_1
XFILLER_59_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30179_ _30179_/A VGND VGND VPWR VPWR _35334_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1038 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34987_ _34987_/CLK _34987_/D VGND VGND VPWR VPWR _34987_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1390 _17843_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24740_ _24740_/A VGND VGND VPWR VPWR _32855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21952_ _22460_/A VGND VGND VPWR VPWR _21952_/X sky130_fd_sc_hd__buf_4
X_33938_ _34197_/CLK _33938_/D VGND VGND VPWR VPWR _33938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20903_ _20674_/X _20899_/X _20902_/X _20684_/X VGND VGND VPWR VPWR _20903_/X sky130_fd_sc_hd__a22o_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24671_ _24671_/A VGND VGND VPWR VPWR _32823_/D sky130_fd_sc_hd__clkbuf_1
X_33869_ _35277_/CLK _33869_/D VGND VGND VPWR VPWR _33869_/Q sky130_fd_sc_hd__dfxtp_1
X_21883_ _21594_/X _21881_/X _21882_/X _21597_/X VGND VGND VPWR VPWR _21883_/X sky130_fd_sc_hd__a22o_1
XFILLER_242_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_99_CLK clkbuf_leaf_99_CLK/A VGND VGND VPWR VPWR _34967_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26410_ _25183_/X _33612_/Q _26412_/S VGND VGND VPWR VPWR _26411_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23622_ _23622_/A VGND VGND VPWR VPWR _32361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20834_ _34514_/Q _32402_/Q _34386_/Q _34322_/Q _20766_/X _20767_/X VGND VGND VPWR
+ VPWR _20834_/X sky130_fd_sc_hd__mux4_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35608_ _35675_/CLK _35608_/D VGND VGND VPWR VPWR _35608_/Q sky130_fd_sc_hd__dfxtp_1
X_27390_ _27390_/A VGND VGND VPWR VPWR _34044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23553_ _23065_/X _32330_/Q _23559_/S VGND VGND VPWR VPWR _23554_/A sky130_fd_sc_hd__mux2_1
X_26341_ _25081_/X _33579_/Q _26341_/S VGND VGND VPWR VPWR _26342_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20765_ _20674_/X _20763_/X _20764_/X _20684_/X VGND VGND VPWR VPWR _20765_/X sky130_fd_sc_hd__a22o_1
X_35539_ _35922_/CLK _35539_/D VGND VGND VPWR VPWR _35539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22504_ _33794_/Q _33730_/Q _33666_/Q _33602_/Q _22502_/X _22503_/X VGND VGND VPWR
+ VPWR _22504_/X sky130_fd_sc_hd__mux4_1
X_29060_ _29060_/A VGND VGND VPWR VPWR _34832_/D sky130_fd_sc_hd__clkbuf_1
X_26272_ _26272_/A VGND VGND VPWR VPWR _33546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23484_ _22963_/X _32297_/Q _23488_/S VGND VGND VPWR VPWR _23485_/A sky130_fd_sc_hd__mux2_1
X_20696_ _22373_/A VGND VGND VPWR VPWR _21759_/A sky130_fd_sc_hd__buf_12
XFILLER_149_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28011_ _28101_/S VGND VGND VPWR VPWR _28030_/S sky130_fd_sc_hd__buf_6
X_25223_ _25223_/A VGND VGND VPWR VPWR _33053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22435_ _22428_/X _22433_/X _22434_/X VGND VGND VPWR VPWR _22469_/A sky130_fd_sc_hd__o21ba_1
XFILLER_167_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25154_ _25153_/X _33026_/Q _25175_/S VGND VGND VPWR VPWR _25155_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22366_ _33278_/Q _36158_/Q _33150_/Q _33086_/Q _22364_/X _22365_/X VGND VGND VPWR
+ VPWR _22366_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24105_ _24105_/A VGND VGND VPWR VPWR _32588_/D sky130_fd_sc_hd__clkbuf_1
X_21317_ _35808_/Q _32184_/Q _35680_/Q _35616_/Q _21207_/X _21208_/X VGND VGND VPWR
+ VPWR _21317_/X sky130_fd_sc_hd__mux4_1
XFILLER_237_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29962_ _29962_/A VGND VGND VPWR VPWR _35231_/D sky130_fd_sc_hd__clkbuf_1
X_25085_ _25187_/S VGND VGND VPWR VPWR _25113_/S sky130_fd_sc_hd__buf_4
X_22297_ _33020_/Q _32956_/Q _32892_/Q _32828_/Q _22295_/X _22296_/X VGND VGND VPWR
+ VPWR _22297_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_CLK clkbuf_6_4__f_CLK/X VGND VGND VPWR VPWR _36200_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_190_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28913_ _30329_/A _28913_/B _31140_/B VGND VGND VPWR VPWR _29046_/S sky130_fd_sc_hd__nor3_4
X_24036_ _24036_/A VGND VGND VPWR VPWR _32555_/D sky130_fd_sc_hd__clkbuf_1
X_21248_ _33182_/Q _32542_/Q _35934_/Q _35870_/Q _20968_/X _20969_/X VGND VGND VPWR
+ VPWR _21248_/X sky130_fd_sc_hd__mux4_1
X_29893_ _35199_/Q _29203_/X _29893_/S VGND VGND VPWR VPWR _29894_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28844_ _28844_/A VGND VGND VPWR VPWR _34732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21179_ _33180_/Q _32540_/Q _35932_/Q _35868_/Q _20968_/X _20969_/X VGND VGND VPWR
+ VPWR _21179_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_1048 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28775_ _28775_/A VGND VGND VPWR VPWR _34700_/D sky130_fd_sc_hd__clkbuf_1
X_25987_ _25156_/X _33411_/Q _25999_/S VGND VGND VPWR VPWR _25988_/A sky130_fd_sc_hd__mux2_1
X_27726_ _27726_/A VGND VGND VPWR VPWR _34202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24938_ _24938_/A VGND VGND VPWR VPWR _32949_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27657_ _34170_/Q _24382_/X _27667_/S VGND VGND VPWR VPWR _27658_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24869_ _24869_/A VGND VGND VPWR VPWR _32916_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_221 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_232 _32136_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17410_ _32756_/Q _32692_/Q _32628_/Q _36084_/Q _17272_/X _17409_/X VGND VGND VPWR
+ VPWR _17410_/X sky130_fd_sc_hd__mux4_1
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_243 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26608_ _25075_/X _33705_/Q _26612_/S VGND VGND VPWR VPWR _26609_/A sky130_fd_sc_hd__mux2_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _19173_/A VGND VGND VPWR VPWR _18390_/X sky130_fd_sc_hd__buf_4
XANTENNA_254 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27588_ _34137_/Q _24280_/X _27604_/S VGND VGND VPWR VPWR _27589_/A sky130_fd_sc_hd__mux2_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_276 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_287 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29327_ _29327_/A VGND VGND VPWR VPWR _34930_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _32498_/Q _32370_/Q _32050_/Q _36018_/Q _17276_/X _17064_/X VGND VGND VPWR
+ VPWR _17341_/X sky130_fd_sc_hd__mux4_1
X_26539_ _25174_/X _33673_/Q _26539_/S VGND VGND VPWR VPWR _26540_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_298 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29258_ _29258_/A VGND VGND VPWR VPWR _34897_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17272_ _17978_/A VGND VGND VPWR VPWR _17272_/X sky130_fd_sc_hd__buf_6
XFILLER_186_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19011_ _20070_/A VGND VGND VPWR VPWR _19011_/X sky130_fd_sc_hd__clkbuf_4
X_28209_ _28236_/S VGND VGND VPWR VPWR _28228_/S sky130_fd_sc_hd__buf_6
X_16223_ _35730_/Q _35090_/Q _34450_/Q _33810_/Q _16049_/X _16051_/X VGND VGND VPWR
+ VPWR _16223_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29189_ _34874_/Q _29188_/X _29204_/S VGND VGND VPWR VPWR _29190_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31220_ _31220_/A VGND VGND VPWR VPWR _35827_/D sky130_fd_sc_hd__clkbuf_1
X_16154_ _16026_/X _16152_/X _16153_/X _16037_/X VGND VGND VPWR VPWR _16154_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31151_ _31151_/A VGND VGND VPWR VPWR _35794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16085_ _16074_/X _16077_/X _16082_/X _16084_/X VGND VGND VPWR VPWR _16085_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_14_CLK clkbuf_6_6__f_CLK/X VGND VGND VPWR VPWR _35801_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_154_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30102_ _30192_/S VGND VGND VPWR VPWR _30121_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_170_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19913_ _35065_/Q _35001_/Q _34937_/Q _34873_/Q _19809_/X _19810_/X VGND VGND VPWR
+ VPWR _19913_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31082_ _35762_/Q _29163_/X _31088_/S VGND VGND VPWR VPWR _31083_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30033_ _35265_/Q _29210_/X _30049_/S VGND VGND VPWR VPWR _30034_/A sky130_fd_sc_hd__mux2_1
X_19844_ _19807_/X _19842_/X _19843_/X _19812_/X VGND VGND VPWR VPWR _19844_/X sky130_fd_sc_hd__a22o_1
X_34910_ _34973_/CLK _34910_/D VGND VGND VPWR VPWR _34910_/Q sky130_fd_sc_hd__dfxtp_1
X_35890_ _35955_/CLK _35890_/D VGND VGND VPWR VPWR _35890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34841_ _35034_/CLK _34841_/D VGND VGND VPWR VPWR _34841_/Q sky130_fd_sc_hd__dfxtp_1
X_19775_ _19495_/X _19773_/X _19774_/X _19500_/X VGND VGND VPWR VPWR _19775_/X sky130_fd_sc_hd__a22o_1
X_16987_ _16702_/X _16985_/X _16986_/X _16708_/X VGND VGND VPWR VPWR _16987_/X sky130_fd_sc_hd__a22o_1
XFILLER_37_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18726_ _18649_/X _18724_/X _18725_/X _18655_/X VGND VGND VPWR VPWR _18726_/X sky130_fd_sc_hd__a22o_1
XFILLER_110_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34772_ _34775_/CLK _34772_/D VGND VGND VPWR VPWR _34772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31984_ _36201_/CLK _31984_/D VGND VGND VPWR VPWR _31984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33723_ _33723_/CLK _33723_/D VGND VGND VPWR VPWR _33723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18657_ _20208_/A VGND VGND VPWR VPWR _18657_/X sky130_fd_sc_hd__clkbuf_4
X_30935_ _35692_/Q _29144_/X _30953_/S VGND VGND VPWR VPWR _30936_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17608_ _17602_/X _17607_/X _17500_/X VGND VGND VPWR VPWR _17616_/C sky130_fd_sc_hd__o21ba_1
XFILLER_91_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33654_ _34295_/CLK _33654_/D VGND VGND VPWR VPWR _33654_/Q sky130_fd_sc_hd__dfxtp_1
X_30866_ _23342_/X _35660_/Q _30868_/S VGND VGND VPWR VPWR _30867_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18588_ _20155_/A VGND VGND VPWR VPWR _18588_/X sky130_fd_sc_hd__buf_4
XFILLER_127_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32605_ _36062_/CLK _32605_/D VGND VGND VPWR VPWR _32605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17539_ _34807_/Q _34743_/Q _34679_/Q _34615_/Q _17288_/X _17289_/X VGND VGND VPWR
+ VPWR _17539_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33585_ _33779_/CLK _33585_/D VGND VGND VPWR VPWR _33585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30797_ _23234_/X _35627_/Q _30797_/S VGND VGND VPWR VPWR _30798_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35324_ _35326_/CLK _35324_/D VGND VGND VPWR VPWR _35324_/Q sky130_fd_sc_hd__dfxtp_1
X_20550_ _18326_/X _20548_/X _20549_/X _18337_/X VGND VGND VPWR VPWR _20550_/X sky130_fd_sc_hd__a22o_1
X_32536_ _36001_/CLK _32536_/D VGND VGND VPWR VPWR _32536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19209_ _19205_/X _19208_/X _19108_/X VGND VGND VPWR VPWR _19210_/D sky130_fd_sc_hd__o21ba_1
X_35255_ _35319_/CLK _35255_/D VGND VGND VPWR VPWR _35255_/Q sky130_fd_sc_hd__dfxtp_1
X_20481_ _18356_/X _20479_/X _20480_/X _18368_/X VGND VGND VPWR VPWR _20481_/X sky130_fd_sc_hd__a22o_1
X_32467_ _35986_/CLK _32467_/D VGND VGND VPWR VPWR _32467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22220_ _22148_/X _22218_/X _22219_/X _22153_/X VGND VGND VPWR VPWR _22220_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34206_ _36200_/CLK _34206_/D VGND VGND VPWR VPWR _34206_/Q sky130_fd_sc_hd__dfxtp_1
X_31418_ _23096_/X _35921_/Q _31430_/S VGND VGND VPWR VPWR _31419_/A sky130_fd_sc_hd__mux2_1
X_35186_ _35250_/CLK _35186_/D VGND VGND VPWR VPWR _35186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32398_ _35282_/CLK _32398_/D VGND VGND VPWR VPWR _32398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22151_ _33784_/Q _33720_/Q _33656_/Q _33592_/Q _22149_/X _22150_/X VGND VGND VPWR
+ VPWR _22151_/X sky130_fd_sc_hd__mux4_1
X_34137_ _34265_/CLK _34137_/D VGND VGND VPWR VPWR _34137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31349_ _31349_/A VGND VGND VPWR VPWR _35888_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21102_ _32730_/Q _32666_/Q _32602_/Q _36058_/Q _20813_/X _20950_/X VGND VGND VPWR
+ VPWR _21102_/X sky130_fd_sc_hd__mux4_1
XTAP_6808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34068_ _34197_/CLK _34068_/D VGND VGND VPWR VPWR _34068_/Q sky130_fd_sc_hd__dfxtp_1
X_22082_ _22075_/X _22080_/X _22081_/X VGND VGND VPWR VPWR _22116_/A sky130_fd_sc_hd__o21ba_1
XTAP_6819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33019_ _33083_/CLK _33019_/D VGND VGND VPWR VPWR _33019_/Q sky130_fd_sc_hd__dfxtp_1
X_21033_ _35800_/Q _32175_/Q _35672_/Q _35608_/Q _20854_/X _20855_/X VGND VGND VPWR
+ VPWR _21033_/X sky130_fd_sc_hd__mux4_1
X_25910_ _25910_/A VGND VGND VPWR VPWR _33374_/D sky130_fd_sc_hd__clkbuf_1
X_26890_ _26890_/A VGND VGND VPWR VPWR _33827_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25841_ _25140_/X _33342_/Q _25843_/S VGND VGND VPWR VPWR _25842_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28560_ _26897_/X _34598_/Q _28570_/S VGND VGND VPWR VPWR _28561_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22984_ _22984_/A VGND VGND VPWR VPWR _32047_/D sky130_fd_sc_hd__clkbuf_1
X_25772_ _25038_/X _33309_/Q _25780_/S VGND VGND VPWR VPWR _25773_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27511_ _27559_/S VGND VGND VPWR VPWR _27530_/S sky130_fd_sc_hd__buf_4
X_24723_ _22883_/X _32847_/Q _24739_/S VGND VGND VPWR VPWR _24724_/A sky130_fd_sc_hd__mux2_1
X_28491_ _28491_/A VGND VGND VPWR VPWR _34565_/D sky130_fd_sc_hd__clkbuf_1
X_21935_ _34034_/Q _33970_/Q _33906_/Q _32242_/Q _21620_/X _21621_/X VGND VGND VPWR
+ VPWR _21935_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27442_ _26844_/X _34069_/Q _27446_/S VGND VGND VPWR VPWR _27443_/A sky130_fd_sc_hd__mux2_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24654_ _24654_/A VGND VGND VPWR VPWR _32815_/D sky130_fd_sc_hd__clkbuf_1
X_21866_ _34288_/Q _34224_/Q _34160_/Q _34096_/Q _21689_/X _21690_/X VGND VGND VPWR
+ VPWR _21866_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20817_ _22582_/A VGND VGND VPWR VPWR _20817_/X sky130_fd_sc_hd__clkbuf_8
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23605_ _23605_/A VGND VGND VPWR VPWR _32353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_242_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27373_ _27373_/A VGND VGND VPWR VPWR _34036_/D sky130_fd_sc_hd__clkbuf_1
X_24585_ _24585_/A VGND VGND VPWR VPWR _32782_/D sky130_fd_sc_hd__clkbuf_1
X_21797_ _22503_/A VGND VGND VPWR VPWR _21797_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_243_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29112_ _29112_/A VGND VGND VPWR VPWR _34849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26324_ _26324_/A VGND VGND VPWR VPWR _33570_/D sky130_fd_sc_hd__clkbuf_1
X_20748_ _20742_/X _20747_/X _20611_/X VGND VGND VPWR VPWR _20772_/A sky130_fd_sc_hd__o21ba_1
X_23536_ _23536_/A VGND VGND VPWR VPWR _32321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29043_ _29043_/A VGND VGND VPWR VPWR _34827_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26255_ _25153_/X _33538_/Q _26269_/S VGND VGND VPWR VPWR _26256_/A sky130_fd_sc_hd__mux2_1
X_23467_ _22938_/X _32289_/Q _23467_/S VGND VGND VPWR VPWR _23468_/A sky130_fd_sc_hd__mux2_1
X_20679_ _22312_/A VGND VGND VPWR VPWR _20679_/X sky130_fd_sc_hd__buf_6
XFILLER_109_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22418_ _35327_/Q _35263_/Q _35199_/Q _32319_/Q _22312_/X _22313_/X VGND VGND VPWR
+ VPWR _22418_/X sky130_fd_sc_hd__mux4_1
X_25206_ _25206_/A VGND VGND VPWR VPWR _33045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23398_ _23398_/A VGND VGND VPWR VPWR _32257_/D sky130_fd_sc_hd__clkbuf_1
X_26186_ _26186_/A VGND VGND VPWR VPWR _33505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25137_ input42/X VGND VGND VPWR VPWR _25137_/X sky130_fd_sc_hd__buf_2
X_22349_ _35069_/Q _35005_/Q _34941_/Q _34877_/Q _22109_/X _22110_/X VGND VGND VPWR
+ VPWR _22349_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29945_ _29945_/A VGND VGND VPWR VPWR _35223_/D sky130_fd_sc_hd__clkbuf_1
X_25068_ _25068_/A VGND VGND VPWR VPWR _32998_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24019_ _22945_/X _32547_/Q _24035_/S VGND VGND VPWR VPWR _24020_/A sky130_fd_sc_hd__mux2_1
X_16910_ _16910_/A _16910_/B _16910_/C _16910_/D VGND VGND VPWR VPWR _16911_/A sky130_fd_sc_hd__or4_4
XFILLER_219_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17890_ _17705_/X _17888_/X _17889_/X _17708_/X VGND VGND VPWR VPWR _17890_/X sky130_fd_sc_hd__a22o_1
X_29876_ _29876_/A VGND VGND VPWR VPWR _35190_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16841_ _16841_/A VGND VGND VPWR VPWR _31971_/D sky130_fd_sc_hd__clkbuf_1
X_28827_ _28827_/A VGND VGND VPWR VPWR _34724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19560_ _35055_/Q _34991_/Q _34927_/Q _34863_/Q _19456_/X _19457_/X VGND VGND VPWR
+ VPWR _19560_/X sky130_fd_sc_hd__mux4_1
X_28758_ _26990_/X _34692_/Q _28768_/S VGND VGND VPWR VPWR _28759_/A sky130_fd_sc_hd__mux2_1
X_16772_ _33506_/Q _33442_/Q _33378_/Q _33314_/Q _16770_/X _16771_/X VGND VGND VPWR
+ VPWR _16772_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18511_ _18443_/X _18509_/X _18510_/X _18446_/X VGND VGND VPWR VPWR _18511_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27709_ _27709_/A VGND VGND VPWR VPWR _34194_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19491_ _19454_/X _19489_/X _19490_/X _19459_/X VGND VGND VPWR VPWR _19491_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28689_ _26888_/X _34659_/Q _28705_/S VGND VGND VPWR VPWR _28690_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ _18436_/X _18439_/X _18440_/X _18441_/X VGND VGND VPWR VPWR _18442_/X sky130_fd_sc_hd__a22o_1
X_30720_ _30720_/A VGND VGND VPWR VPWR _35590_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_3_CLK clkbuf_leaf_9_CLK/A VGND VGND VPWR VPWR _34782_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18373_ _20061_/A VGND VGND VPWR VPWR _19449_/A sky130_fd_sc_hd__buf_12
X_30651_ _30651_/A VGND VGND VPWR VPWR _35557_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _17149_/X _17322_/X _17323_/X _17152_/X VGND VGND VPWR VPWR _17324_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33370_ _33946_/CLK _33370_/D VGND VGND VPWR VPWR _33370_/Q sky130_fd_sc_hd__dfxtp_1
X_30582_ _23319_/X _35525_/Q _30590_/S VGND VGND VPWR VPWR _30583_/A sky130_fd_sc_hd__mux2_1
X_32321_ _32967_/CLK _32321_/D VGND VGND VPWR VPWR _32321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17255_ _17249_/X _17254_/X _17147_/X VGND VGND VPWR VPWR _17263_/C sky130_fd_sc_hd__o21ba_1
XFILLER_70_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16206_ _33746_/Q _33682_/Q _33618_/Q _33554_/Q _16137_/X _16138_/X VGND VGND VPWR
+ VPWR _16206_/X sky130_fd_sc_hd__mux4_1
X_35040_ _35040_/CLK _35040_/D VGND VGND VPWR VPWR _35040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32252_ _34171_/CLK _32252_/D VGND VGND VPWR VPWR _32252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17186_ _34797_/Q _34733_/Q _34669_/Q _34605_/Q _16935_/X _16936_/X VGND VGND VPWR
+ VPWR _17186_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_6_50__f_CLK clkbuf_5_25_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_50__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_31_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31203_ _31203_/A VGND VGND VPWR VPWR _35819_/D sky130_fd_sc_hd__clkbuf_1
X_16137_ _17902_/A VGND VGND VPWR VPWR _16137_/X sky130_fd_sc_hd__buf_6
XFILLER_196_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32183_ _35807_/CLK _32183_/D VGND VGND VPWR VPWR _32183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31134_ _35787_/Q _29240_/X _31138_/S VGND VGND VPWR VPWR _31135_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16068_ _17865_/A VGND VGND VPWR VPWR _16068_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_233_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35942_ _35942_/CLK _35942_/D VGND VGND VPWR VPWR _35942_/Q sky130_fd_sc_hd__dfxtp_1
X_31065_ _35754_/Q _29138_/X _31067_/S VGND VGND VPWR VPWR _31066_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30016_ _35257_/Q _29185_/X _30028_/S VGND VGND VPWR VPWR _30017_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19827_ _19708_/X _19825_/X _19826_/X _19714_/X VGND VGND VPWR VPWR _19827_/X sky130_fd_sc_hd__a22o_1
X_35873_ _35940_/CLK _35873_/D VGND VGND VPWR VPWR _35873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_919 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34824_ _35337_/CLK _34824_/D VGND VGND VPWR VPWR _34824_/Q sky130_fd_sc_hd__dfxtp_1
X_19758_ _35765_/Q _35125_/Q _34485_/Q _33845_/Q _19440_/X _19441_/X VGND VGND VPWR
+ VPWR _19758_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18709_ _35031_/Q _34967_/Q _34903_/Q _34839_/Q _18392_/X _18394_/X VGND VGND VPWR
+ VPWR _18709_/X sky130_fd_sc_hd__mux4_1
X_34755_ _34819_/CLK _34755_/D VGND VGND VPWR VPWR _34755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31967_ _34970_/CLK _31967_/D VGND VGND VPWR VPWR _31967_/Q sky130_fd_sc_hd__dfxtp_1
X_19689_ _33203_/Q _32563_/Q _35955_/Q _35891_/Q _19374_/X _19375_/X VGND VGND VPWR
+ VPWR _19689_/X sky130_fd_sc_hd__mux4_1
X_21720_ _33772_/Q _33708_/Q _33644_/Q _33580_/Q _21443_/X _21444_/X VGND VGND VPWR
+ VPWR _21720_/X sky130_fd_sc_hd__mux4_1
X_33706_ _34281_/CLK _33706_/D VGND VGND VPWR VPWR _33706_/Q sky130_fd_sc_hd__dfxtp_1
X_30918_ _35684_/Q _29120_/X _30932_/S VGND VGND VPWR VPWR _30919_/A sky130_fd_sc_hd__mux2_1
X_34686_ _35837_/CLK _34686_/D VGND VGND VPWR VPWR _34686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31898_ _23267_/X _36149_/Q _31898_/S VGND VGND VPWR VPWR _31899_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21651_ _33514_/Q _33450_/Q _33386_/Q _33322_/Q _21370_/X _21371_/X VGND VGND VPWR
+ VPWR _21651_/X sky130_fd_sc_hd__mux4_1
X_33637_ _33702_/CLK _33637_/D VGND VGND VPWR VPWR _33637_/Q sky130_fd_sc_hd__dfxtp_1
X_30849_ _30849_/A VGND VGND VPWR VPWR _35651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20602_ _22373_/A VGND VGND VPWR VPWR _22511_/A sky130_fd_sc_hd__buf_12
X_24370_ _24401_/A VGND VGND VPWR VPWR _24398_/S sky130_fd_sc_hd__buf_4
XFILLER_240_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33568_ _34010_/CLK _33568_/D VGND VGND VPWR VPWR _33568_/Q sky130_fd_sc_hd__dfxtp_1
X_21582_ _34024_/Q _33960_/Q _33896_/Q _32215_/Q _21267_/X _21268_/X VGND VGND VPWR
+ VPWR _21582_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23321_ _23321_/A VGND VGND VPWR VPWR _32224_/D sky130_fd_sc_hd__clkbuf_1
X_32519_ _36039_/CLK _32519_/D VGND VGND VPWR VPWR _32519_/Q sky130_fd_sc_hd__dfxtp_1
X_20533_ _33228_/Q _32588_/Q _35980_/Q _35916_/Q _18375_/X _18376_/X VGND VGND VPWR
+ VPWR _20533_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_976 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35307_ _35307_/CLK _35307_/D VGND VGND VPWR VPWR _35307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33499_ _36194_/CLK _33499_/D VGND VGND VPWR VPWR _33499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23252_ _23252_/A VGND VGND VPWR VPWR _32201_/D sky130_fd_sc_hd__clkbuf_1
X_26040_ _25035_/X _33436_/Q _26050_/S VGND VGND VPWR VPWR _26041_/A sky130_fd_sc_hd__mux2_1
X_20464_ _19449_/A _20462_/X _20463_/X _19452_/A VGND VGND VPWR VPWR _20464_/X sky130_fd_sc_hd__a22o_1
XFILLER_165_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35238_ _35239_/CLK _35238_/D VGND VGND VPWR VPWR _35238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22203_ _22556_/A VGND VGND VPWR VPWR _22203_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_10_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23183_ _23183_/A VGND VGND VPWR VPWR _32174_/D sky130_fd_sc_hd__clkbuf_1
X_35169_ _35296_/CLK _35169_/D VGND VGND VPWR VPWR _35169_/Q sky130_fd_sc_hd__dfxtp_1
X_20395_ _33800_/Q _33736_/Q _33672_/Q _33608_/Q _20202_/X _20203_/X VGND VGND VPWR
+ VPWR _20395_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22134_ _21947_/X _22132_/X _22133_/X _21950_/X VGND VGND VPWR VPWR _22134_/X sky130_fd_sc_hd__a22o_1
XTAP_6605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27991_ _26853_/X _34328_/Q _28009_/S VGND VGND VPWR VPWR _27992_/A sky130_fd_sc_hd__mux2_1
XTAP_6616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput250 _32117_/Q VGND VGND VPWR VPWR D3[39] sky130_fd_sc_hd__buf_2
Xoutput261 _32127_/Q VGND VGND VPWR VPWR D3[49] sky130_fd_sc_hd__buf_2
XFILLER_47_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput272 _32137_/Q VGND VGND VPWR VPWR D3[59] sky130_fd_sc_hd__buf_2
X_29730_ _29730_/A VGND VGND VPWR VPWR _35121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26942_ _26942_/A VGND VGND VPWR VPWR _33844_/D sky130_fd_sc_hd__clkbuf_1
X_22065_ _35317_/Q _35253_/Q _35189_/Q _32309_/Q _21959_/X _21960_/X VGND VGND VPWR
+ VPWR _22065_/X sky130_fd_sc_hd__mux4_1
XTAP_6649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21016_ _20736_/X _21014_/X _21015_/X _20741_/X VGND VGND VPWR VPWR _21016_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29661_ _29661_/A VGND VGND VPWR VPWR _35088_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26873_ _26872_/X _33822_/Q _26882_/S VGND VGND VPWR VPWR _26874_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28612_ _26974_/X _34623_/Q _28612_/S VGND VGND VPWR VPWR _28613_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25824_ _25872_/S VGND VGND VPWR VPWR _25843_/S sky130_fd_sc_hd__buf_4
X_29592_ _35056_/Q _29157_/X _29602_/S VGND VGND VPWR VPWR _29593_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28543_ _26872_/X _34590_/Q _28549_/S VGND VGND VPWR VPWR _28544_/A sky130_fd_sc_hd__mux2_1
X_25755_ _25013_/X _33301_/Q _25759_/S VGND VGND VPWR VPWR _25756_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22967_ _22966_/X _32042_/Q _22970_/S VGND VGND VPWR VPWR _22968_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24706_ _24706_/A VGND VGND VPWR VPWR _32840_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28474_ _28474_/A VGND VGND VPWR VPWR _34557_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21918_ _35569_/Q _35505_/Q _35441_/Q _35377_/Q _21850_/X _21851_/X VGND VGND VPWR
+ VPWR _21918_/X sky130_fd_sc_hd__mux4_1
XFILLER_243_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25686_ _25686_/A VGND VGND VPWR VPWR _33269_/D sky130_fd_sc_hd__clkbuf_1
X_22898_ input61/X VGND VGND VPWR VPWR _22898_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_230_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27425_ _27425_/A VGND VGND VPWR VPWR _34061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24637_ _24637_/A VGND VGND VPWR VPWR _32807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21849_ _21594_/X _21847_/X _21848_/X _21597_/X VGND VGND VPWR VPWR _21849_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27356_ _34028_/Q _24338_/X _27374_/S VGND VGND VPWR VPWR _27357_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24568_ _24568_/A VGND VGND VPWR VPWR _32776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26307_ _26307_/A VGND VGND VPWR VPWR _33562_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23519_ _23519_/A VGND VGND VPWR VPWR _32313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27287_ _27014_/X _33996_/Q _27289_/S VGND VGND VPWR VPWR _27288_/A sky130_fd_sc_hd__mux2_1
X_24499_ _24499_/A VGND VGND VPWR VPWR _32743_/D sky130_fd_sc_hd__clkbuf_1
X_29026_ _34819_/Q _24410_/X _29038_/S VGND VGND VPWR VPWR _29027_/A sky130_fd_sc_hd__mux2_1
X_17040_ _35305_/Q _35241_/Q _35177_/Q _32297_/Q _17006_/X _17007_/X VGND VGND VPWR
+ VPWR _17040_/X sky130_fd_sc_hd__mux4_1
X_26238_ _25128_/X _33530_/Q _26248_/S VGND VGND VPWR VPWR _26239_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26169_ _25026_/X _33497_/Q _26185_/S VGND VGND VPWR VPWR _26170_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18991_ _18748_/X _18989_/X _18990_/X _18753_/X VGND VGND VPWR VPWR _18991_/X sky130_fd_sc_hd__a22o_1
XFILLER_152_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17942_ _33539_/Q _33475_/Q _33411_/Q _33347_/Q _17829_/X _17830_/X VGND VGND VPWR
+ VPWR _17942_/X sky130_fd_sc_hd__mux4_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29928_ _35215_/Q _29055_/X _29944_/S VGND VGND VPWR VPWR _29929_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17873_ _17548_/X _17871_/X _17872_/X _17553_/X VGND VGND VPWR VPWR _17873_/X sky130_fd_sc_hd__a22o_1
X_29859_ _29859_/A VGND VGND VPWR VPWR _35182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19612_ _19608_/X _19611_/X _19436_/X _19437_/X VGND VGND VPWR VPWR _19629_/B sky130_fd_sc_hd__o211a_1
X_16824_ _16710_/X _16822_/X _16823_/X _16714_/X VGND VGND VPWR VPWR _16824_/X sky130_fd_sc_hd__a22o_1
X_32870_ _36007_/CLK _32870_/D VGND VGND VPWR VPWR _32870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31821_ _23093_/X _36112_/Q _31835_/S VGND VGND VPWR VPWR _31822_/A sky130_fd_sc_hd__mux2_1
X_19543_ _32495_/Q _32367_/Q _32047_/Q _36015_/Q _19223_/X _19364_/X VGND VGND VPWR
+ VPWR _19543_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_1041 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16755_ _33185_/Q _32545_/Q _35937_/Q _35873_/Q _16721_/X _16722_/X VGND VGND VPWR
+ VPWR _16755_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34540_ _35304_/CLK _34540_/D VGND VGND VPWR VPWR _34540_/Q sky130_fd_sc_hd__dfxtp_1
X_19474_ _19355_/X _19472_/X _19473_/X _19361_/X VGND VGND VPWR VPWR _19474_/X sky130_fd_sc_hd__a22o_1
X_31752_ _31752_/A VGND VGND VPWR VPWR _36079_/D sky130_fd_sc_hd__clkbuf_1
X_16686_ _34783_/Q _34719_/Q _34655_/Q _34591_/Q _16582_/X _16583_/X VGND VGND VPWR
+ VPWR _16686_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18425_ _18356_/X _18423_/X _18424_/X _18368_/X VGND VGND VPWR VPWR _18425_/X sky130_fd_sc_hd__a22o_1
X_30703_ _30703_/A VGND VGND VPWR VPWR _35582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34471_ _34859_/CLK _34471_/D VGND VGND VPWR VPWR _34471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31683_ _31683_/A VGND VGND VPWR VPWR _36046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33422_ _33490_/CLK _33422_/D VGND VGND VPWR VPWR _33422_/Q sky130_fd_sc_hd__dfxtp_1
X_36210_ _36211_/CLK _36210_/D VGND VGND VPWR VPWR _36210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18356_ _20160_/A VGND VGND VPWR VPWR _18356_/X sky130_fd_sc_hd__buf_4
XFILLER_194_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30634_ _30634_/A VGND VGND VPWR VPWR _35549_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_221_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_36141_ _36141_/CLK _36141_/D VGND VGND VPWR VPWR _36141_/Q sky130_fd_sc_hd__dfxtp_1
X_17307_ _33265_/Q _36145_/Q _33137_/Q _33073_/Q _17058_/X _17059_/X VGND VGND VPWR
+ VPWR _17307_/X sky130_fd_sc_hd__mux4_1
X_33353_ _33545_/CLK _33353_/D VGND VGND VPWR VPWR _33353_/Q sky130_fd_sc_hd__dfxtp_1
X_18287_ _20206_/A VGND VGND VPWR VPWR _18287_/X sky130_fd_sc_hd__buf_4
X_30565_ _23294_/X _35517_/Q _30569_/S VGND VGND VPWR VPWR _30566_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32304_ _35758_/CLK _32304_/D VGND VGND VPWR VPWR _32304_/Q sky130_fd_sc_hd__dfxtp_1
X_17238_ _17202_/X _17236_/X _17237_/X _17205_/X VGND VGND VPWR VPWR _17238_/X sky130_fd_sc_hd__a22o_1
X_36072_ _36072_/CLK _36072_/D VGND VGND VPWR VPWR _36072_/Q sky130_fd_sc_hd__dfxtp_1
X_33284_ _33922_/CLK _33284_/D VGND VGND VPWR VPWR _33284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30496_ _23130_/X _35484_/Q _30506_/S VGND VGND VPWR VPWR _30497_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35023_ _35282_/CLK _35023_/D VGND VGND VPWR VPWR _35023_/Q sky130_fd_sc_hd__dfxtp_1
X_32235_ _36136_/CLK _32235_/D VGND VGND VPWR VPWR _32235_/Q sky130_fd_sc_hd__dfxtp_1
X_17169_ _34029_/Q _33965_/Q _33901_/Q _32237_/Q _17020_/X _17021_/X VGND VGND VPWR
+ VPWR _17169_/X sky130_fd_sc_hd__mux4_1
XFILLER_235_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32166_ _35664_/CLK _32166_/D VGND VGND VPWR VPWR _32166_/Q sky130_fd_sc_hd__dfxtp_1
X_20180_ _20061_/X _20178_/X _20179_/X _20067_/X VGND VGND VPWR VPWR _20180_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31117_ _31117_/A VGND VGND VPWR VPWR _35778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32097_ _35807_/CLK _32097_/D VGND VGND VPWR VPWR _32097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35925_ _35925_/CLK _35925_/D VGND VGND VPWR VPWR _35925_/Q sky130_fd_sc_hd__dfxtp_1
X_31048_ _31138_/S VGND VGND VPWR VPWR _31067_/S sky130_fd_sc_hd__buf_4
XFILLER_9_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35856_ _35921_/CLK _35856_/D VGND VGND VPWR VPWR _35856_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23870_ _22926_/X _32477_/Q _23878_/S VGND VGND VPWR VPWR _23871_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22821_ _22817_/X _22820_/X _22434_/A VGND VGND VPWR VPWR _22843_/A sky130_fd_sc_hd__o21ba_1
X_34807_ _35638_/CLK _34807_/D VGND VGND VPWR VPWR _34807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35787_ _35787_/CLK _35787_/D VGND VGND VPWR VPWR _35787_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_809 _22904_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32999_ _36072_/CLK _32999_/D VGND VGND VPWR VPWR _32999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25540_ _25540_/A VGND VGND VPWR VPWR _33201_/D sky130_fd_sc_hd__clkbuf_1
X_22752_ _22748_/X _22751_/X _22467_/X VGND VGND VPWR VPWR _22753_/D sky130_fd_sc_hd__o21ba_1
X_34738_ _34932_/CLK _34738_/D VGND VGND VPWR VPWR _34738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21703_ _21699_/X _21702_/X _21383_/X _21384_/X VGND VGND VPWR VPWR _21718_/B sky130_fd_sc_hd__o211a_1
X_22683_ _33223_/Q _32583_/Q _35975_/Q _35911_/Q _22380_/X _22381_/X VGND VGND VPWR
+ VPWR _22683_/X sky130_fd_sc_hd__mux4_1
X_25471_ _25471_/A VGND VGND VPWR VPWR _33168_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34669_ _35304_/CLK _34669_/D VGND VGND VPWR VPWR _34669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27210_ _26900_/X _33959_/Q _27218_/S VGND VGND VPWR VPWR _27211_/A sky130_fd_sc_hd__mux2_1
X_24422_ input53/X VGND VGND VPWR VPWR _24422_/X sky130_fd_sc_hd__buf_6
X_21634_ _21594_/X _21632_/X _21633_/X _21597_/X VGND VGND VPWR VPWR _21634_/X sky130_fd_sc_hd__a22o_1
X_28190_ _28190_/A VGND VGND VPWR VPWR _34422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27141_ _27141_/A VGND VGND VPWR VPWR _33926_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_240_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24353_ _24353_/A VGND VGND VPWR VPWR _32688_/D sky130_fd_sc_hd__clkbuf_1
X_21565_ _35559_/Q _35495_/Q _35431_/Q _35367_/Q _21497_/X _21498_/X VGND VGND VPWR
+ VPWR _21565_/X sky130_fd_sc_hd__mux4_1
XFILLER_205_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23304_ _23346_/S VGND VGND VPWR VPWR _23334_/S sky130_fd_sc_hd__buf_4
X_20516_ _34316_/Q _34252_/Q _34188_/Q _34124_/Q _18345_/X _18346_/X VGND VGND VPWR
+ VPWR _20516_/X sky130_fd_sc_hd__mux4_1
X_24284_ _32666_/Q _24283_/X _24305_/S VGND VGND VPWR VPWR _24285_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27072_ _27072_/A VGND VGND VPWR VPWR _33893_/D sky130_fd_sc_hd__clkbuf_1
X_21496_ _21241_/X _21494_/X _21495_/X _21244_/X VGND VGND VPWR VPWR _21496_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26023_ _25010_/X _33428_/Q _26029_/S VGND VGND VPWR VPWR _26024_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_1019 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23235_ _32196_/Q _23234_/X _23235_/S VGND VGND VPWR VPWR _23236_/A sky130_fd_sc_hd__mux2_1
X_20447_ _35337_/Q _35273_/Q _35209_/Q _32329_/Q _18388_/X _18390_/X VGND VGND VPWR
+ VPWR _20447_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23166_ _23166_/A VGND VGND VPWR VPWR _32166_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20378_ _20374_/X _20377_/X _20142_/X _20143_/X VGND VGND VPWR VPWR _20393_/B sky130_fd_sc_hd__o211a_1
XFILLER_162_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1076 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22117_ _22117_/A VGND VGND VPWR VPWR _36214_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1208 _23145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23097_ _32145_/Q _23096_/X _23115_/S VGND VGND VPWR VPWR _23098_/A sky130_fd_sc_hd__mux2_1
XTAP_6435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27974_ _26829_/X _34320_/Q _27988_/S VGND VGND VPWR VPWR _27975_/A sky130_fd_sc_hd__mux2_1
XANTENNA_1219 _24267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29713_ _29713_/A VGND VGND VPWR VPWR _35113_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26925_ input27/X VGND VGND VPWR VPWR _26925_/X sky130_fd_sc_hd__buf_4
XFILLER_0_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22048_ _21802_/X _22046_/X _22047_/X _21805_/X VGND VGND VPWR VPWR _22048_/X sky130_fd_sc_hd__a22o_1
XTAP_6479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29644_ _35081_/Q _29234_/X _29644_/S VGND VGND VPWR VPWR _29645_/A sky130_fd_sc_hd__mux2_1
XTAP_5767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26856_ _26856_/A VGND VGND VPWR VPWR _33816_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25807_ _25807_/A VGND VGND VPWR VPWR _33325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29575_ _35048_/Q _29132_/X _29581_/S VGND VGND VPWR VPWR _29576_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26787_ _26787_/A VGND VGND VPWR VPWR _33789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23999_ _23999_/A VGND VGND VPWR VPWR _32537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28526_ _26847_/X _34582_/Q _28528_/S VGND VGND VPWR VPWR _28527_/A sky130_fd_sc_hd__mux2_1
X_16540_ _16536_/X _16539_/X _16430_/X _16431_/X VGND VGND VPWR VPWR _16557_/B sky130_fd_sc_hd__o211a_2
XFILLER_21_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25738_ _25738_/A VGND VGND VPWR VPWR _26685_/B sky130_fd_sc_hd__buf_12
XFILLER_147_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16471_ _16357_/X _16469_/X _16470_/X _16361_/X VGND VGND VPWR VPWR _16471_/X sky130_fd_sc_hd__a22o_1
X_28457_ _28457_/A VGND VGND VPWR VPWR _34549_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25669_ _33261_/Q _24342_/X _25685_/S VGND VGND VPWR VPWR _25670_/A sky130_fd_sc_hd__mux2_1
X_18210_ _35083_/Q _35019_/Q _34955_/Q _34891_/Q _16079_/X _16081_/X VGND VGND VPWR
+ VPWR _18210_/X sky130_fd_sc_hd__mux4_1
X_27408_ _34053_/Q _24416_/X _27416_/S VGND VGND VPWR VPWR _27409_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19190_ _32485_/Q _32357_/Q _32037_/Q _36005_/Q _18870_/X _19011_/X VGND VGND VPWR
+ VPWR _19190_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28388_ _28388_/A VGND VGND VPWR VPWR _34516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18141_ _15977_/X _18139_/X _18140_/X _15987_/X VGND VGND VPWR VPWR _18141_/X sky130_fd_sc_hd__a22o_1
XFILLER_212_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27339_ _34020_/Q _24314_/X _27353_/S VGND VGND VPWR VPWR _27340_/A sky130_fd_sc_hd__mux2_1
X_18072_ _32775_/Q _32711_/Q _32647_/Q _36103_/Q _17978_/X _17762_/X VGND VGND VPWR
+ VPWR _18072_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30350_ _23114_/X _35415_/Q _30350_/S VGND VGND VPWR VPWR _30351_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_929 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29009_ _34811_/Q _24385_/X _29017_/S VGND VGND VPWR VPWR _29010_/A sky130_fd_sc_hd__mux2_1
X_17023_ _16849_/X _17019_/X _17022_/X _16852_/X VGND VGND VPWR VPWR _17023_/X sky130_fd_sc_hd__a22o_1
X_30281_ _30281_/A VGND VGND VPWR VPWR _35382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32020_ _35986_/CLK _32020_/D VGND VGND VPWR VPWR _32020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18974_ _18649_/X _18972_/X _18973_/X _18655_/X VGND VGND VPWR VPWR _18974_/X sky130_fd_sc_hd__a22o_1
XFILLER_234_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17925_ _33218_/Q _32578_/Q _35970_/Q _35906_/Q _17780_/X _17781_/X VGND VGND VPWR
+ VPWR _17925_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33971_ _34228_/CLK _33971_/D VGND VGND VPWR VPWR _33971_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_294_CLK clkbuf_6_51__f_CLK/X VGND VGND VPWR VPWR _35903_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35710_ _35710_/CLK _35710_/D VGND VGND VPWR VPWR _35710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17856_ _34816_/Q _34752_/Q _34688_/Q _34624_/Q _17641_/X _17642_/X VGND VGND VPWR
+ VPWR _17856_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32922_ _34146_/CLK _32922_/D VGND VGND VPWR VPWR _32922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16807_ _16801_/X _16802_/X _16805_/X _16806_/X VGND VGND VPWR VPWR _16807_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35641_ _35834_/CLK _35641_/D VGND VGND VPWR VPWR _35641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17787_ _17502_/X _17785_/X _17786_/X _17505_/X VGND VGND VPWR VPWR _17787_/X sky130_fd_sc_hd__a22o_1
X_32853_ _32983_/CLK _32853_/D VGND VGND VPWR VPWR _32853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31804_ _31804_/A VGND VGND VPWR VPWR _36104_/D sky130_fd_sc_hd__clkbuf_1
X_19526_ _20232_/A VGND VGND VPWR VPWR _19526_/X sky130_fd_sc_hd__buf_4
XFILLER_53_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16738_ _34273_/Q _34209_/Q _34145_/Q _34081_/Q _16736_/X _16737_/X VGND VGND VPWR
+ VPWR _16738_/X sky130_fd_sc_hd__mux4_1
X_32784_ _36049_/CLK _32784_/D VGND VGND VPWR VPWR _32784_/Q sky130_fd_sc_hd__dfxtp_1
X_35572_ _36021_/CLK _35572_/D VGND VGND VPWR VPWR _35572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34523_ _34970_/CLK _34523_/D VGND VGND VPWR VPWR _34523_/Q sky130_fd_sc_hd__dfxtp_1
X_19457_ _19457_/A VGND VGND VPWR VPWR _19457_/X sky130_fd_sc_hd__clkbuf_4
X_31735_ _31735_/A VGND VGND VPWR VPWR _36071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16669_ _34015_/Q _33951_/Q _33887_/Q _32159_/Q _16667_/X _16668_/X VGND VGND VPWR
+ VPWR _16669_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18408_ _20146_/A VGND VGND VPWR VPWR _18408_/X sky130_fd_sc_hd__buf_6
X_31666_ _36039_/Q input53/X _31670_/S VGND VGND VPWR VPWR _31667_/A sky130_fd_sc_hd__mux2_1
X_34454_ _35667_/CLK _34454_/D VGND VGND VPWR VPWR _34454_/Q sky130_fd_sc_hd__dfxtp_1
X_19388_ _33771_/Q _33707_/Q _33643_/Q _33579_/Q _19143_/X _19144_/X VGND VGND VPWR
+ VPWR _19388_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18339_ input81/X VGND VGND VPWR VPWR _20142_/A sky130_fd_sc_hd__buf_12
X_33405_ _33789_/CLK _33405_/D VGND VGND VPWR VPWR _33405_/Q sky130_fd_sc_hd__dfxtp_1
X_30617_ _30617_/A VGND VGND VPWR VPWR _35541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34385_ _36204_/CLK _34385_/D VGND VGND VPWR VPWR _34385_/Q sky130_fd_sc_hd__dfxtp_1
X_31597_ _36006_/Q input17/X _31607_/S VGND VGND VPWR VPWR _31598_/A sky130_fd_sc_hd__mux2_1
XFILLER_198_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33336_ _34297_/CLK _33336_/D VGND VGND VPWR VPWR _33336_/Q sky130_fd_sc_hd__dfxtp_1
X_21350_ _21346_/X _21349_/X _21030_/X _21031_/X VGND VGND VPWR VPWR _21365_/B sky130_fd_sc_hd__o211a_1
X_36124_ _36124_/CLK _36124_/D VGND VGND VPWR VPWR _36124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30548_ _23267_/X _35509_/Q _30548_/S VGND VGND VPWR VPWR _30549_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20301_ _20160_/X _20299_/X _20300_/X _20165_/X VGND VGND VPWR VPWR _20301_/X sky130_fd_sc_hd__a22o_1
X_36055_ _36055_/CLK _36055_/D VGND VGND VPWR VPWR _36055_/Q sky130_fd_sc_hd__dfxtp_1
X_21281_ _21241_/X _21279_/X _21280_/X _21244_/X VGND VGND VPWR VPWR _21281_/X sky130_fd_sc_hd__a22o_1
X_33267_ _36147_/CLK _33267_/D VGND VGND VPWR VPWR _33267_/Q sky130_fd_sc_hd__dfxtp_1
X_30479_ _23105_/X _35476_/Q _30485_/S VGND VGND VPWR VPWR _30480_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23020_ _23019_/X _32059_/Q _23032_/S VGND VGND VPWR VPWR _23021_/A sky130_fd_sc_hd__mux2_1
X_20232_ _20232_/A VGND VGND VPWR VPWR _20232_/X sky130_fd_sc_hd__buf_4
X_32218_ _35903_/CLK _32218_/D VGND VGND VPWR VPWR _32218_/Q sky130_fd_sc_hd__dfxtp_1
X_35006_ _35517_/CLK _35006_/D VGND VGND VPWR VPWR _35006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33198_ _35822_/CLK _33198_/D VGND VGND VPWR VPWR _33198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32149_ _35280_/CLK _32149_/D VGND VGND VPWR VPWR _32149_/Q sky130_fd_sc_hd__dfxtp_1
X_20163_ _20163_/A VGND VGND VPWR VPWR _20163_/X sky130_fd_sc_hd__buf_4
XFILLER_115_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24971_ _23050_/X _32965_/Q _24979_/S VGND VGND VPWR VPWR _24972_/A sky130_fd_sc_hd__mux2_1
X_20094_ _33791_/Q _33727_/Q _33663_/Q _33599_/Q _19849_/X _19850_/X VGND VGND VPWR
+ VPWR _20094_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_285_CLK clkbuf_6_56__f_CLK/X VGND VGND VPWR VPWR _36027_/CLK sky130_fd_sc_hd__clkbuf_16
X_26710_ _26710_/A VGND VGND VPWR VPWR _33752_/D sky130_fd_sc_hd__clkbuf_1
X_35908_ _35970_/CLK _35908_/D VGND VGND VPWR VPWR _35908_/Q sky130_fd_sc_hd__dfxtp_1
X_23922_ _23970_/S VGND VGND VPWR VPWR _23941_/S sky130_fd_sc_hd__buf_4
XTAP_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27690_ _34186_/Q _24431_/X _27696_/S VGND VGND VPWR VPWR _27691_/A sky130_fd_sc_hd__mux2_1
XTAP_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26641_ _26641_/A VGND VGND VPWR VPWR _33720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35839_ _35903_/CLK _35839_/D VGND VGND VPWR VPWR _35839_/Q sky130_fd_sc_hd__dfxtp_1
X_23853_ _22901_/X _32469_/Q _23857_/S VGND VGND VPWR VPWR _23854_/A sky130_fd_sc_hd__mux2_1
XTAP_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_606 _18435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29360_ _23310_/X _34946_/Q _29374_/S VGND VGND VPWR VPWR _29361_/A sky130_fd_sc_hd__mux2_1
X_22804_ _20597_/X _22802_/X _22803_/X _20603_/X VGND VGND VPWR VPWR _22804_/X sky130_fd_sc_hd__a22o_1
XANTENNA_617 _18539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26572_ _26683_/S VGND VGND VPWR VPWR _26591_/S sky130_fd_sc_hd__buf_4
XANTENNA_628 _18757_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20996_ _20957_/X _20994_/X _20995_/X _20961_/X VGND VGND VPWR VPWR _20996_/X sky130_fd_sc_hd__a22o_1
X_23784_ _23000_/X _32437_/Q _23784_/S VGND VGND VPWR VPWR _23785_/A sky130_fd_sc_hd__mux2_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_639 _19315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_1001 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28311_ _34480_/Q _24351_/X _28321_/S VGND VGND VPWR VPWR _28312_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25523_ _25523_/A VGND VGND VPWR VPWR _33193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22735_ _32521_/Q _32393_/Q _32073_/Q _36041_/Q _22582_/X _21607_/A VGND VGND VPWR
+ VPWR _22735_/X sky130_fd_sc_hd__mux4_1
X_29291_ _29291_/A VGND VGND VPWR VPWR _34913_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28242_ _34447_/Q _24249_/X _28258_/S VGND VGND VPWR VPWR _28243_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25454_ _25180_/X _33163_/Q _25458_/S VGND VGND VPWR VPWR _25455_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22666_ _34311_/Q _34247_/Q _34183_/Q _34119_/Q _22395_/X _22396_/X VGND VGND VPWR
+ VPWR _22666_/X sky130_fd_sc_hd__mux4_1
XFILLER_213_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24405_ _32705_/Q _24404_/X _24429_/S VGND VGND VPWR VPWR _24406_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28173_ _28173_/A VGND VGND VPWR VPWR _34414_/D sky130_fd_sc_hd__clkbuf_1
X_21617_ _34281_/Q _34217_/Q _34153_/Q _34089_/Q _21336_/X _21337_/X VGND VGND VPWR
+ VPWR _21617_/X sky130_fd_sc_hd__mux4_1
X_25385_ _25078_/X _33130_/Q _25387_/S VGND VGND VPWR VPWR _25386_/A sky130_fd_sc_hd__mux2_1
X_22597_ _35332_/Q _35268_/Q _35204_/Q _32324_/Q _22312_/X _22313_/X VGND VGND VPWR
+ VPWR _22597_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27124_ _27124_/A VGND VGND VPWR VPWR _33918_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24336_ _32683_/Q _24335_/X _24336_/S VGND VGND VPWR VPWR _24337_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21548_ _21442_/X _21546_/X _21547_/X _21447_/X VGND VGND VPWR VPWR _21548_/X sky130_fd_sc_hd__a22o_1
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27055_ _27055_/A VGND VGND VPWR VPWR _33885_/D sky130_fd_sc_hd__clkbuf_1
X_21479_ _21479_/A VGND VGND VPWR VPWR _36196_/D sky130_fd_sc_hd__clkbuf_1
X_24267_ input62/X VGND VGND VPWR VPWR _24267_/X sky130_fd_sc_hd__buf_6
XFILLER_119_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26006_ _26006_/A VGND VGND VPWR VPWR _33420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23218_ _32190_/Q _23217_/X _23235_/S VGND VGND VPWR VPWR _23219_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24198_ _24198_/A VGND VGND VPWR VPWR _32631_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1095 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23149_ _23421_/S VGND VGND VPWR VPWR _23350_/S sky130_fd_sc_hd__buf_4
XTAP_6221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1005 _17901_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1016 _17995_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1027 _17865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1038 _17152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27957_ _27957_/A VGND VGND VPWR VPWR _34312_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1049 _17867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17710_ _17704_/X _17709_/X _17500_/X VGND VGND VPWR VPWR _17720_/C sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_276_CLK clkbuf_6_58__f_CLK/X VGND VGND VPWR VPWR _33787_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26908_ _26908_/A VGND VGND VPWR VPWR _33833_/D sky130_fd_sc_hd__clkbuf_1
X_18690_ _18686_/X _18689_/X _18311_/X VGND VGND VPWR VPWR _18712_/A sky130_fd_sc_hd__o21ba_1
XTAP_5564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27888_ _27888_/A VGND VGND VPWR VPWR _34279_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_208_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17641_ _17994_/A VGND VGND VPWR VPWR _17641_/X sky130_fd_sc_hd__buf_6
XTAP_5597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29627_ _29627_/A VGND VGND VPWR VPWR _35072_/D sky130_fd_sc_hd__clkbuf_1
X_26839_ _26838_/X _33811_/Q _26851_/S VGND VGND VPWR VPWR _26840_/A sky130_fd_sc_hd__mux2_1
XTAP_4863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1041 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17572_ _33208_/Q _32568_/Q _35960_/Q _35896_/Q _17427_/X _17428_/X VGND VGND VPWR
+ VPWR _17572_/X sky130_fd_sc_hd__mux4_1
X_29558_ _35040_/Q _29107_/X _29560_/S VGND VGND VPWR VPWR _29559_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19311_ _35048_/Q _34984_/Q _34920_/Q _34856_/Q _19103_/X _19104_/X VGND VGND VPWR
+ VPWR _19311_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28509_ _28641_/S VGND VGND VPWR VPWR _28528_/S sky130_fd_sc_hd__buf_6
XFILLER_204_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16523_ _16448_/X _16521_/X _16522_/X _16453_/X VGND VGND VPWR VPWR _16523_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29489_ _29489_/A VGND VGND VPWR VPWR _35007_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31520_ _31520_/A VGND VGND VPWR VPWR _35969_/D sky130_fd_sc_hd__clkbuf_1
X_19242_ _19101_/X _19240_/X _19241_/X _19106_/X VGND VGND VPWR VPWR _19242_/X sky130_fd_sc_hd__a22o_1
XFILLER_220_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16454_ _16448_/X _16449_/X _16452_/X _16453_/X VGND VGND VPWR VPWR _16454_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31451_ _23145_/X _35937_/Q _31451_/S VGND VGND VPWR VPWR _31452_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19173_ _19173_/A VGND VGND VPWR VPWR _19173_/X sky130_fd_sc_hd__buf_4
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16385_ _34263_/Q _34199_/Q _34135_/Q _34071_/Q _16383_/X _16384_/X VGND VGND VPWR
+ VPWR _16385_/X sky130_fd_sc_hd__mux4_2
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_200_CLK clkbuf_6_51__f_CLK/X VGND VGND VPWR VPWR _35906_/CLK sky130_fd_sc_hd__clkbuf_16
X_18124_ _18124_/A VGND VGND VPWR VPWR _32008_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_185_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30402_ _30402_/A VGND VGND VPWR VPWR _35439_/D sky130_fd_sc_hd__clkbuf_1
X_34170_ _34299_/CLK _34170_/D VGND VGND VPWR VPWR _34170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31382_ _35904_/Q input46/X _31400_/S VGND VGND VPWR VPWR _31383_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33121_ _36128_/CLK _33121_/D VGND VGND VPWR VPWR _33121_/Q sky130_fd_sc_hd__dfxtp_1
X_18055_ _18051_/X _18054_/X _17853_/X VGND VGND VPWR VPWR _18063_/C sky130_fd_sc_hd__o21ba_1
X_30333_ _30333_/A VGND VGND VPWR VPWR _35406_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_2 _32114_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17006_ _17712_/A VGND VGND VPWR VPWR _17006_/X sky130_fd_sc_hd__buf_4
X_33052_ _36124_/CLK _33052_/D VGND VGND VPWR VPWR _33052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30264_ _30264_/A VGND VGND VPWR VPWR _35374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32003_ _34202_/CLK _32003_/D VGND VGND VPWR VPWR _32003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30195_ _30327_/S VGND VGND VPWR VPWR _30214_/S sky130_fd_sc_hd__buf_4
X_18957_ _34526_/Q _32414_/Q _34398_/Q _34334_/Q _18819_/X _18820_/X VGND VGND VPWR
+ VPWR _18957_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_267_CLK clkbuf_6_59__f_CLK/X VGND VGND VPWR VPWR _36160_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_239_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17908_ _17908_/A VGND VGND VPWR VPWR _17908_/X sky130_fd_sc_hd__clkbuf_8
X_33954_ _34146_/CLK _33954_/D VGND VGND VPWR VPWR _33954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18888_ _35036_/Q _34972_/Q _34908_/Q _34844_/Q _18750_/X _18751_/X VGND VGND VPWR
+ VPWR _18888_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32905_ _36107_/CLK _32905_/D VGND VGND VPWR VPWR _32905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17839_ _32512_/Q _32384_/Q _32064_/Q _36032_/Q _17629_/X _17770_/X VGND VGND VPWR
+ VPWR _17839_/X sky130_fd_sc_hd__mux4_1
X_33885_ _34205_/CLK _33885_/D VGND VGND VPWR VPWR _33885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20850_ _32467_/Q _32339_/Q _32019_/Q _35987_/Q _20817_/X _22463_/A VGND VGND VPWR
+ VPWR _20850_/X sky130_fd_sc_hd__mux4_1
X_35624_ _35879_/CLK _35624_/D VGND VGND VPWR VPWR _35624_/Q sky130_fd_sc_hd__dfxtp_1
X_32836_ _32901_/CLK _32836_/D VGND VGND VPWR VPWR _32836_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19509_ _33262_/Q _36142_/Q _33134_/Q _33070_/Q _19358_/X _19359_/X VGND VGND VPWR
+ VPWR _19509_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20781_ _32721_/Q _32657_/Q _32593_/Q _36049_/Q _22462_/A _22313_/A VGND VGND VPWR
+ VPWR _20781_/X sky130_fd_sc_hd__mux4_1
X_35555_ _35555_/CLK _35555_/D VGND VGND VPWR VPWR _35555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32767_ _36097_/CLK _32767_/D VGND VGND VPWR VPWR _32767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34506_ _35788_/CLK _34506_/D VGND VGND VPWR VPWR _34506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22520_ _22516_/X _22519_/X _22442_/X _22443_/X VGND VGND VPWR VPWR _22537_/B sky130_fd_sc_hd__o211a_1
XFILLER_74_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31718_ _31718_/A VGND VGND VPWR VPWR _36063_/D sky130_fd_sc_hd__clkbuf_1
X_32698_ _36090_/CLK _32698_/D VGND VGND VPWR VPWR _32698_/Q sky130_fd_sc_hd__dfxtp_1
X_35486_ _35808_/CLK _35486_/D VGND VGND VPWR VPWR _35486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34437_ _35781_/CLK _34437_/D VGND VGND VPWR VPWR _34437_/Q sky130_fd_sc_hd__dfxtp_1
X_22451_ _33216_/Q _32576_/Q _35968_/Q _35904_/Q _22380_/X _22381_/X VGND VGND VPWR
+ VPWR _22451_/X sky130_fd_sc_hd__mux4_1
X_31649_ _36031_/Q input44/X _31649_/S VGND VGND VPWR VPWR _31650_/A sky130_fd_sc_hd__mux2_1
XFILLER_206_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21402_ _34530_/Q _32418_/Q _34402_/Q _34338_/Q _21119_/X _21120_/X VGND VGND VPWR
+ VPWR _21402_/X sky130_fd_sc_hd__mux4_1
X_25170_ _25170_/A VGND VGND VPWR VPWR _33031_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22382_ _33214_/Q _32574_/Q _35966_/Q _35902_/Q _22380_/X _22381_/X VGND VGND VPWR
+ VPWR _22382_/X sky130_fd_sc_hd__mux4_1
X_34368_ _36038_/CLK _34368_/D VGND VGND VPWR VPWR _34368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36107_ _36107_/CLK _36107_/D VGND VGND VPWR VPWR _36107_/Q sky130_fd_sc_hd__dfxtp_1
X_24121_ _22895_/X _32595_/Q _24129_/S VGND VGND VPWR VPWR _24122_/A sky130_fd_sc_hd__mux2_1
X_21333_ _21333_/A _21333_/B _21333_/C _21333_/D VGND VGND VPWR VPWR _21334_/A sky130_fd_sc_hd__or4_1
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33319_ _35991_/CLK _33319_/D VGND VGND VPWR VPWR _33319_/Q sky130_fd_sc_hd__dfxtp_1
X_34299_ _34299_/CLK _34299_/D VGND VGND VPWR VPWR _34299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36038_ _36038_/CLK _36038_/D VGND VGND VPWR VPWR _36038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24052_ _22994_/X _32563_/Q _24056_/S VGND VGND VPWR VPWR _24053_/A sky130_fd_sc_hd__mux2_1
X_21264_ _34271_/Q _34207_/Q _34143_/Q _34079_/Q _20983_/X _20984_/X VGND VGND VPWR
+ VPWR _21264_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20215_ _33282_/Q _36162_/Q _33154_/Q _33090_/Q _20064_/X _20065_/X VGND VGND VPWR
+ VPWR _20215_/X sky130_fd_sc_hd__mux4_1
X_23003_ input35/X VGND VGND VPWR VPWR _23003_/X sky130_fd_sc_hd__clkbuf_4
Xmax_cap282 _29046_/S VGND VGND VPWR VPWR _28998_/A sky130_fd_sc_hd__buf_12
XFILLER_176_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28860_ _28860_/A VGND VGND VPWR VPWR _34740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21195_ _21089_/X _21193_/X _21194_/X _21094_/X VGND VGND VPWR VPWR _21195_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27811_ _34243_/Q _24410_/X _27823_/S VGND VGND VPWR VPWR _27812_/A sky130_fd_sc_hd__mux2_1
X_20146_ _20146_/A VGND VGND VPWR VPWR _20146_/X sky130_fd_sc_hd__buf_4
X_28791_ _28791_/A VGND VGND VPWR VPWR _34707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_258_CLK clkbuf_6_60__f_CLK/X VGND VGND VPWR VPWR _36100_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27742_ _34210_/Q _24307_/X _27760_/S VGND VGND VPWR VPWR _27743_/A sky130_fd_sc_hd__mux2_1
X_20077_ _35774_/Q _35134_/Q _34494_/Q _33854_/Q _19793_/X _19794_/X VGND VGND VPWR
+ VPWR _20077_/X sky130_fd_sc_hd__mux4_1
X_24954_ _23025_/X _32957_/Q _24958_/S VGND VGND VPWR VPWR _24955_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_27__f_CLK clkbuf_5_13_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_27__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XTAP_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23905_ _23905_/A VGND VGND VPWR VPWR _32493_/D sky130_fd_sc_hd__clkbuf_1
X_27673_ _27673_/A VGND VGND VPWR VPWR _34177_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24885_ _22923_/X _32924_/Q _24895_/S VGND VGND VPWR VPWR _24886_/A sky130_fd_sc_hd__mux2_1
XTAP_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29412_ _29412_/A VGND VGND VPWR VPWR _34970_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_403 _36210_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26624_ _26624_/A VGND VGND VPWR VPWR _33712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23836_ _25462_/A input83/X _23561_/B VGND VGND VPWR VPWR _23837_/A sky130_fd_sc_hd__or3b_1
XFILLER_122_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_414 _36212_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_425 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_436 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29343_ _23283_/X _34938_/Q _29353_/S VGND VGND VPWR VPWR _29344_/A sky130_fd_sc_hd__mux2_1
XANTENNA_447 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26555_ _26555_/A VGND VGND VPWR VPWR _33679_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_458 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23767_ _23767_/A VGND VGND VPWR VPWR _32428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20979_ _20975_/X _20978_/X _20700_/X VGND VGND VPWR VPWR _20980_/D sky130_fd_sc_hd__o21ba_1
XANTENNA_469 _31992_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_430_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _34283_/CLK sky130_fd_sc_hd__clkbuf_16
X_25506_ _25506_/A VGND VGND VPWR VPWR _33185_/D sky130_fd_sc_hd__clkbuf_1
X_22718_ _22455_/X _22716_/X _22717_/X _22458_/X VGND VGND VPWR VPWR _22718_/X sky130_fd_sc_hd__a22o_1
XFILLER_159_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29274_ _23121_/X _34905_/Q _29290_/S VGND VGND VPWR VPWR _29275_/A sky130_fd_sc_hd__mux2_1
XFILLER_214_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26486_ _26486_/A VGND VGND VPWR VPWR _33647_/D sky130_fd_sc_hd__clkbuf_1
X_23698_ _30329_/B _29049_/B VGND VGND VPWR VPWR _28913_/B sky130_fd_sc_hd__nand2_2
X_28225_ _28225_/A VGND VGND VPWR VPWR _34439_/D sky130_fd_sc_hd__clkbuf_1
X_25437_ _25437_/A VGND VGND VPWR VPWR _33154_/D sky130_fd_sc_hd__clkbuf_1
X_22649_ _35846_/Q _32225_/Q _35718_/Q _35654_/Q _20589_/X _20591_/X VGND VGND VPWR
+ VPWR _22649_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_1072 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16170_ _16087_/X _16168_/X _16169_/X _16097_/X VGND VGND VPWR VPWR _16170_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28156_ _28156_/A VGND VGND VPWR VPWR _34406_/D sky130_fd_sc_hd__clkbuf_1
X_25368_ _25458_/S VGND VGND VPWR VPWR _25387_/S sky130_fd_sc_hd__buf_4
XFILLER_166_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27107_ _26946_/X _33910_/Q _27125_/S VGND VGND VPWR VPWR _27108_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24319_ _24319_/A VGND VGND VPWR VPWR _32677_/D sky130_fd_sc_hd__clkbuf_1
X_28087_ _26996_/X _34374_/Q _28093_/S VGND VGND VPWR VPWR _28088_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25299_ _25299_/A VGND VGND VPWR VPWR _33089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27038_ _27038_/A VGND VGND VPWR VPWR _33877_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19860_ _19854_/X _19859_/X _19781_/X VGND VGND VPWR VPWR _19884_/A sky130_fd_sc_hd__o21ba_1
XFILLER_134_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18811_ _18588_/X _18809_/X _18810_/X _18591_/X VGND VGND VPWR VPWR _18811_/X sky130_fd_sc_hd__a22o_1
XTAP_6040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput94 _31963_/Q VGND VGND VPWR VPWR D1[13] sky130_fd_sc_hd__buf_2
X_19791_ _19785_/X _19788_/X _19789_/X _19790_/X VGND VGND VPWR VPWR _19816_/B sky130_fd_sc_hd__o211a_1
XTAP_6062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28989_ _28989_/A VGND VGND VPWR VPWR _34801_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_249_CLK clkbuf_6_63__f_CLK/X VGND VGND VPWR VPWR _34057_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18742_ _18737_/X _18740_/X _18741_/X VGND VGND VPWR VPWR _18757_/C sky130_fd_sc_hd__o21ba_1
XFILLER_231_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18673_ _34774_/Q _34710_/Q _34646_/Q _34582_/Q _18529_/X _18530_/X VGND VGND VPWR
+ VPWR _18673_/X sky130_fd_sc_hd__mux4_1
X_30951_ _35700_/Q _29169_/X _30953_/S VGND VGND VPWR VPWR _30952_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17624_ _17620_/X _17623_/X _17481_/X VGND VGND VPWR VPWR _17650_/A sky130_fd_sc_hd__o21ba_1
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33670_ _34312_/CLK _33670_/D VGND VGND VPWR VPWR _33670_/Q sky130_fd_sc_hd__dfxtp_1
X_30882_ _35667_/Q _29067_/X _30890_/S VGND VGND VPWR VPWR _30883_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _17908_/A VGND VGND VPWR VPWR _17555_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32621_ _36077_/CLK _32621_/D VGND VGND VPWR VPWR _32621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_970 _31678_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_421_CLK clkbuf_6_38__f_CLK/X VGND VGND VPWR VPWR _35315_/CLK sky130_fd_sc_hd__clkbuf_16
X_16506_ _32986_/Q _32922_/Q _32858_/Q _32794_/Q _16283_/X _16284_/X VGND VGND VPWR
+ VPWR _16506_/X sky130_fd_sc_hd__mux4_1
X_35340_ _35340_/CLK _35340_/D VGND VGND VPWR VPWR _35340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32552_ _35947_/CLK _32552_/D VGND VGND VPWR VPWR _32552_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_981 _17902_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_992 _17860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17486_ _32502_/Q _32374_/Q _32054_/Q _36022_/Q _17276_/X _17417_/X VGND VGND VPWR
+ VPWR _17486_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31503_ _31503_/A VGND VGND VPWR VPWR _35961_/D sky130_fd_sc_hd__clkbuf_1
X_16437_ _16288_/X _16433_/X _16436_/X _16291_/X VGND VGND VPWR VPWR _16437_/X sky130_fd_sc_hd__a22o_1
X_19225_ _32998_/Q _32934_/Q _32870_/Q _32806_/Q _18936_/X _18937_/X VGND VGND VPWR
+ VPWR _19225_/X sky130_fd_sc_hd__mux4_1
X_35271_ _35339_/CLK _35271_/D VGND VGND VPWR VPWR _35271_/Q sky130_fd_sc_hd__dfxtp_1
X_32483_ _36003_/CLK _32483_/D VGND VGND VPWR VPWR _32483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31434_ _31434_/A VGND VGND VPWR VPWR _35928_/D sky130_fd_sc_hd__clkbuf_1
X_34222_ _34222_/CLK _34222_/D VGND VGND VPWR VPWR _34222_/Q sky130_fd_sc_hd__dfxtp_1
X_19156_ _33252_/Q _36132_/Q _33124_/Q _33060_/Q _19005_/X _19006_/X VGND VGND VPWR
+ VPWR _19156_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16368_ _17931_/A VGND VGND VPWR VPWR _16368_/X sky130_fd_sc_hd__buf_6
XFILLER_199_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18107_ _17154_/A _18105_/X _18106_/X _17159_/A VGND VGND VPWR VPWR _18107_/X sky130_fd_sc_hd__a22o_1
XFILLER_160_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34153_ _34153_/CLK _34153_/D VGND VGND VPWR VPWR _34153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31365_ _35896_/Q input37/X _31379_/S VGND VGND VPWR VPWR _31366_/A sky130_fd_sc_hd__mux2_1
X_19087_ _20294_/A VGND VGND VPWR VPWR _19087_/X sky130_fd_sc_hd__buf_6
XFILLER_173_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16299_ _34772_/Q _34708_/Q _34644_/Q _34580_/Q _16229_/X _16230_/X VGND VGND VPWR
+ VPWR _16299_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18038_ _33542_/Q _33478_/Q _33414_/Q _33350_/Q _17829_/X _17830_/X VGND VGND VPWR
+ VPWR _18038_/X sky130_fd_sc_hd__mux4_1
X_30316_ _30316_/A VGND VGND VPWR VPWR _35399_/D sky130_fd_sc_hd__clkbuf_1
X_33104_ _36114_/CLK _33104_/D VGND VGND VPWR VPWR _33104_/Q sky130_fd_sc_hd__dfxtp_1
X_34084_ _34149_/CLK _34084_/D VGND VGND VPWR VPWR _34084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31296_ _31296_/A VGND VGND VPWR VPWR _35863_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_488_CLK clkbuf_6_2__f_CLK/X VGND VGND VPWR VPWR _35808_/CLK sky130_fd_sc_hd__clkbuf_16
X_33035_ _35977_/CLK _33035_/D VGND VGND VPWR VPWR _33035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30247_ _30247_/A VGND VGND VPWR VPWR _35366_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20000_ _20155_/A VGND VGND VPWR VPWR _20000_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_154_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30178_ _35334_/Q _29225_/X _30184_/S VGND VGND VPWR VPWR _30179_/A sky130_fd_sc_hd__mux2_1
X_19989_ _19855_/X _19987_/X _19988_/X _19858_/X VGND VGND VPWR VPWR _19989_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34986_ _34986_/CLK _34986_/D VGND VGND VPWR VPWR _34986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1380 _28506_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1391 _17932_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33937_ _36228_/CLK _33937_/D VGND VGND VPWR VPWR _33937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21951_ _21947_/X _21948_/X _21949_/X _21950_/X VGND VGND VPWR VPWR _21951_/X sky130_fd_sc_hd__a22o_1
XFILLER_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20902_ _35284_/Q _35220_/Q _35156_/Q _32276_/Q _20900_/X _20901_/X VGND VGND VPWR
+ VPWR _20902_/X sky130_fd_sc_hd__mux4_1
XFILLER_227_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24670_ _23007_/X _32823_/Q _24686_/S VGND VGND VPWR VPWR _24671_/A sky130_fd_sc_hd__mux2_1
X_33868_ _35853_/CLK _33868_/D VGND VGND VPWR VPWR _33868_/Q sky130_fd_sc_hd__dfxtp_1
X_21882_ _35760_/Q _35120_/Q _34480_/Q _33840_/Q _21740_/X _21741_/X VGND VGND VPWR
+ VPWR _21882_/X sky130_fd_sc_hd__mux4_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35607_ _35671_/CLK _35607_/D VGND VGND VPWR VPWR _35607_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23621_ _32361_/Q _23228_/X _23625_/S VGND VGND VPWR VPWR _23622_/A sky130_fd_sc_hd__mux2_1
X_20833_ _20674_/X _20831_/X _20832_/X _20684_/X VGND VGND VPWR VPWR _20833_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32819_ _35765_/CLK _32819_/D VGND VGND VPWR VPWR _32819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33799_ _34819_/CLK _33799_/D VGND VGND VPWR VPWR _33799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_412_CLK clkbuf_6_33__f_CLK/X VGND VGND VPWR VPWR _36011_/CLK sky130_fd_sc_hd__clkbuf_16
X_26340_ _26340_/A VGND VGND VPWR VPWR _33578_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23552_ _23552_/A VGND VGND VPWR VPWR _32329_/D sky130_fd_sc_hd__clkbuf_1
X_35538_ _35922_/CLK _35538_/D VGND VGND VPWR VPWR _35538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20764_ _35280_/Q _35216_/Q _35152_/Q _32272_/Q _20679_/X _20681_/X VGND VGND VPWR
+ VPWR _20764_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_946 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22503_ _22503_/A VGND VGND VPWR VPWR _22503_/X sky130_fd_sc_hd__buf_6
XFILLER_17_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26271_ _25177_/X _33546_/Q _26277_/S VGND VGND VPWR VPWR _26272_/A sky130_fd_sc_hd__mux2_1
X_35469_ _35792_/CLK _35469_/D VGND VGND VPWR VPWR _35469_/Q sky130_fd_sc_hd__dfxtp_1
X_20695_ _35022_/Q _34958_/Q _34894_/Q _34830_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _20695_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23483_ _23483_/A VGND VGND VPWR VPWR _32296_/D sky130_fd_sc_hd__clkbuf_1
X_28010_ _28010_/A VGND VGND VPWR VPWR _34337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25222_ _25038_/X _33053_/Q _25230_/S VGND VGND VPWR VPWR _25223_/A sky130_fd_sc_hd__mux2_1
X_22434_ _22434_/A VGND VGND VPWR VPWR _22434_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_17_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_17_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_104_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25153_ input48/X VGND VGND VPWR VPWR _25153_/X sky130_fd_sc_hd__buf_2
XFILLER_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22365_ _22370_/A VGND VGND VPWR VPWR _22365_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_164_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24104_ _23071_/X _32588_/Q _24106_/S VGND VGND VPWR VPWR _24105_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21316_ _21309_/X _21315_/X _21030_/X _21031_/X VGND VGND VPWR VPWR _21333_/B sky130_fd_sc_hd__o211a_1
X_22296_ _22430_/A VGND VGND VPWR VPWR _22296_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29961_ _35231_/Q _29104_/X _29965_/S VGND VGND VPWR VPWR _29962_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25084_ input24/X VGND VGND VPWR VPWR _25084_/X sky130_fd_sc_hd__buf_6
XFILLER_117_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_479_CLK clkbuf_6_9__f_CLK/X VGND VGND VPWR VPWR _35928_/CLK sky130_fd_sc_hd__clkbuf_16
X_28912_ _28912_/A VGND VGND VPWR VPWR _34765_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21247_ _35550_/Q _35486_/Q _35422_/Q _35358_/Q _21144_/X _21145_/X VGND VGND VPWR
+ VPWR _21247_/X sky130_fd_sc_hd__mux4_1
X_24035_ _22969_/X _32555_/Q _24035_/S VGND VGND VPWR VPWR _24036_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29892_ _29892_/A VGND VGND VPWR VPWR _35198_/D sky130_fd_sc_hd__clkbuf_1
X_21178_ _35548_/Q _35484_/Q _35420_/Q _35356_/Q _21144_/X _21145_/X VGND VGND VPWR
+ VPWR _21178_/X sky130_fd_sc_hd__mux4_1
X_28843_ _26915_/X _34732_/Q _28861_/S VGND VGND VPWR VPWR _28844_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20129_ _20129_/A VGND VGND VPWR VPWR _20129_/X sky130_fd_sc_hd__buf_4
X_28774_ _27014_/X _34700_/Q _28776_/S VGND VGND VPWR VPWR _28775_/A sky130_fd_sc_hd__mux2_1
XFILLER_213_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25986_ _25986_/A VGND VGND VPWR VPWR _33410_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_219_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27725_ _34202_/Q _24283_/X _27739_/S VGND VGND VPWR VPWR _27726_/A sky130_fd_sc_hd__mux2_1
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24937_ _23000_/X _32949_/Q _24937_/S VGND VGND VPWR VPWR _24938_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27656_ _27656_/A VGND VGND VPWR VPWR _34169_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_200 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24868_ _22898_/X _32916_/Q _24874_/S VGND VGND VPWR VPWR _24869_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_211 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_222 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26607_ _26607_/A VGND VGND VPWR VPWR _33704_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23819_ _23819_/A VGND VGND VPWR VPWR _32453_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_233 _32136_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27587_ _27587_/A VGND VGND VPWR VPWR _34136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24799_ _24799_/A VGND VGND VPWR VPWR _32883_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_266 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_403_CLK clkbuf_6_32__f_CLK/X VGND VGND VPWR VPWR _35818_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_277 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17340_ _17055_/X _17338_/X _17339_/X _17061_/X VGND VGND VPWR VPWR _17340_/X sky130_fd_sc_hd__a22o_1
X_29326_ _23256_/X _34930_/Q _29332_/S VGND VGND VPWR VPWR _29327_/A sky130_fd_sc_hd__mux2_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26538_ _26538_/A VGND VGND VPWR VPWR _33672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_288 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_299 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29257_ _23096_/X _34897_/Q _29269_/S VGND VGND VPWR VPWR _29258_/A sky130_fd_sc_hd__mux2_1
X_17271_ _17267_/X _17270_/X _17128_/X VGND VGND VPWR VPWR _17297_/A sky130_fd_sc_hd__o21ba_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26469_ _26469_/A VGND VGND VPWR VPWR _33639_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19010_ _20208_/A VGND VGND VPWR VPWR _19010_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_70_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16222_ _35794_/Q _32168_/Q _35666_/Q _35602_/Q _16045_/X _16046_/X VGND VGND VPWR
+ VPWR _16222_/X sky130_fd_sc_hd__mux4_1
X_28208_ _28208_/A VGND VGND VPWR VPWR _34431_/D sky130_fd_sc_hd__clkbuf_1
X_29188_ input39/X VGND VGND VPWR VPWR _29188_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_195_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16153_ _32976_/Q _32912_/Q _32848_/Q _32784_/Q _16033_/X _16035_/X VGND VGND VPWR
+ VPWR _16153_/X sky130_fd_sc_hd__mux4_1
X_28139_ _28139_/A VGND VGND VPWR VPWR _34398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31150_ _35794_/Q input45/X _31160_/S VGND VGND VPWR VPWR _31151_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16084_ _17152_/A VGND VGND VPWR VPWR _16084_/X sky130_fd_sc_hd__buf_4
XFILLER_181_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30101_ _30101_/A VGND VGND VPWR VPWR _35297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1088 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19912_ _34553_/Q _32441_/Q _34425_/Q _34361_/Q _19878_/X _19879_/X VGND VGND VPWR
+ VPWR _19912_/X sky130_fd_sc_hd__mux4_1
X_31081_ _31081_/A VGND VGND VPWR VPWR _35761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30032_ _30032_/A VGND VGND VPWR VPWR _35264_/D sky130_fd_sc_hd__clkbuf_1
X_19843_ _35063_/Q _34999_/Q _34935_/Q _34871_/Q _19809_/X _19810_/X VGND VGND VPWR
+ VPWR _19843_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34840_ _35292_/CLK _34840_/D VGND VGND VPWR VPWR _34840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19774_ _34294_/Q _34230_/Q _34166_/Q _34102_/Q _19742_/X _19743_/X VGND VGND VPWR
+ VPWR _19774_/X sky130_fd_sc_hd__mux4_1
XFILLER_209_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16986_ _33256_/Q _36136_/Q _33128_/Q _33064_/Q _16705_/X _16706_/X VGND VGND VPWR
+ VPWR _16986_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18725_ _33240_/Q _36120_/Q _33112_/Q _33048_/Q _18652_/X _18653_/X VGND VGND VPWR
+ VPWR _18725_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34771_ _34775_/CLK _34771_/D VGND VGND VPWR VPWR _34771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31983_ _36201_/CLK _31983_/D VGND VGND VPWR VPWR _31983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33722_ _33787_/CLK _33722_/D VGND VGND VPWR VPWR _33722_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_10__f_CLK clkbuf_5_5_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_10__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_224_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18656_ _18649_/X _18651_/X _18654_/X _18655_/X VGND VGND VPWR VPWR _18656_/X sky130_fd_sc_hd__a22o_1
X_30934_ _31003_/S VGND VGND VPWR VPWR _30953_/S sky130_fd_sc_hd__buf_4
XTAP_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17607_ _17352_/X _17605_/X _17606_/X _17355_/X VGND VGND VPWR VPWR _17607_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30865_ _30865_/A VGND VGND VPWR VPWR _35659_/D sky130_fd_sc_hd__clkbuf_1
X_33653_ _34292_/CLK _33653_/D VGND VGND VPWR VPWR _33653_/Q sky130_fd_sc_hd__dfxtp_1
X_18587_ _18581_/X _18586_/X _18340_/X _18342_/X VGND VGND VPWR VPWR _18608_/B sky130_fd_sc_hd__o211a_1
XFILLER_79_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32604_ _36127_/CLK _32604_/D VGND VGND VPWR VPWR _32604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17538_ _17534_/X _17537_/X _17500_/X VGND VGND VPWR VPWR _17546_/C sky130_fd_sc_hd__o21ba_1
X_30796_ _30796_/A VGND VGND VPWR VPWR _35626_/D sky130_fd_sc_hd__clkbuf_1
X_33584_ _33775_/CLK _33584_/D VGND VGND VPWR VPWR _33584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_946 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35323_ _35515_/CLK _35323_/D VGND VGND VPWR VPWR _35323_/Q sky130_fd_sc_hd__dfxtp_1
X_32535_ _35863_/CLK _32535_/D VGND VGND VPWR VPWR _32535_/Q sky130_fd_sc_hd__dfxtp_1
X_17469_ _17154_/X _17467_/X _17468_/X _17159_/X VGND VGND VPWR VPWR _17469_/X sky130_fd_sc_hd__a22o_1
XFILLER_242_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19208_ _19101_/X _19206_/X _19207_/X _19106_/X VGND VGND VPWR VPWR _19208_/X sky130_fd_sc_hd__a22o_1
X_20480_ _35082_/Q _35018_/Q _34954_/Q _34890_/Q _18379_/X _18381_/X VGND VGND VPWR
+ VPWR _20480_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35254_ _35319_/CLK _35254_/D VGND VGND VPWR VPWR _35254_/Q sky130_fd_sc_hd__dfxtp_1
X_32466_ _36052_/CLK _32466_/D VGND VGND VPWR VPWR _32466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34205_ _34205_/CLK _34205_/D VGND VGND VPWR VPWR _34205_/Q sky130_fd_sc_hd__dfxtp_1
X_31417_ _31417_/A VGND VGND VPWR VPWR _35920_/D sky130_fd_sc_hd__clkbuf_1
X_19139_ _19135_/X _19138_/X _19108_/X VGND VGND VPWR VPWR _19140_/D sky130_fd_sc_hd__o21ba_1
X_32397_ _34124_/CLK _32397_/D VGND VGND VPWR VPWR _32397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35185_ _35308_/CLK _35185_/D VGND VGND VPWR VPWR _35185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22150_ _22503_/A VGND VGND VPWR VPWR _22150_/X sky130_fd_sc_hd__clkbuf_4
X_34136_ _34266_/CLK _34136_/D VGND VGND VPWR VPWR _34136_/Q sky130_fd_sc_hd__dfxtp_1
X_31348_ _35888_/Q input28/X _31358_/S VGND VGND VPWR VPWR _31349_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_1155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21101_ _21095_/X _21100_/X _21022_/X VGND VGND VPWR VPWR _21125_/A sky130_fd_sc_hd__o21ba_1
XFILLER_218_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22081_ _22434_/A VGND VGND VPWR VPWR _22081_/X sky130_fd_sc_hd__buf_2
XTAP_6809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34067_ _34260_/CLK _34067_/D VGND VGND VPWR VPWR _34067_/Q sky130_fd_sc_hd__dfxtp_1
X_31279_ _35855_/Q input12/X _31295_/S VGND VGND VPWR VPWR _31280_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21032_ _21026_/X _21029_/X _21030_/X _21031_/X VGND VGND VPWR VPWR _21057_/B sky130_fd_sc_hd__o211a_1
XFILLER_173_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33018_ _36090_/CLK _33018_/D VGND VGND VPWR VPWR _33018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25840_ _25840_/A VGND VGND VPWR VPWR _33341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25771_ _25771_/A VGND VGND VPWR VPWR _33308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22983_ _22982_/X _32047_/Q _23001_/S VGND VGND VPWR VPWR _22984_/A sky130_fd_sc_hd__mux2_1
X_34969_ _35293_/CLK _34969_/D VGND VGND VPWR VPWR _34969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27510_ _27510_/A VGND VGND VPWR VPWR _34101_/D sky130_fd_sc_hd__clkbuf_1
X_24722_ _24722_/A VGND VGND VPWR VPWR _32846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28490_ _26993_/X _34565_/Q _28498_/S VGND VGND VPWR VPWR _28491_/A sky130_fd_sc_hd__mux2_1
X_21934_ _33522_/Q _33458_/Q _33394_/Q _33330_/Q _21723_/X _21724_/X VGND VGND VPWR
+ VPWR _21934_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27441_ _27441_/A VGND VGND VPWR VPWR _34068_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24653_ _22982_/X _32815_/Q _24665_/S VGND VGND VPWR VPWR _24654_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21865_ _33776_/Q _33712_/Q _33648_/Q _33584_/Q _21796_/X _21797_/X VGND VGND VPWR
+ VPWR _21865_/X sky130_fd_sc_hd__mux4_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23604_ _32353_/Q _23145_/X _23604_/S VGND VGND VPWR VPWR _23605_/A sky130_fd_sc_hd__mux2_1
X_20816_ _20614_/X _20814_/X _20815_/X _20623_/X VGND VGND VPWR VPWR _20816_/X sky130_fd_sc_hd__a22o_1
X_27372_ _34036_/Q _24363_/X _27374_/S VGND VGND VPWR VPWR _27373_/A sky130_fd_sc_hd__mux2_1
X_24584_ _22875_/X _32782_/Q _24602_/S VGND VGND VPWR VPWR _24585_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21796_ _22502_/A VGND VGND VPWR VPWR _21796_/X sky130_fd_sc_hd__buf_4
X_29111_ _34849_/Q _29110_/X _29111_/S VGND VGND VPWR VPWR _29112_/A sky130_fd_sc_hd__mux2_1
X_26323_ _25053_/X _33570_/Q _26341_/S VGND VGND VPWR VPWR _26324_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_5_0_0_CLK clkbuf_5_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_5_0_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_51_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23535_ _23038_/X _32321_/Q _23551_/S VGND VGND VPWR VPWR _23536_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20747_ _20743_/X _20744_/X _20745_/X _20746_/X VGND VGND VPWR VPWR _20747_/X sky130_fd_sc_hd__a22o_1
X_29042_ _34827_/Q _24434_/X _29046_/S VGND VGND VPWR VPWR _29043_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26254_ _26254_/A VGND VGND VPWR VPWR _33537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23466_ _23466_/A VGND VGND VPWR VPWR _32288_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20678_ _22578_/A VGND VGND VPWR VPWR _22312_/A sky130_fd_sc_hd__buf_12
X_25205_ _25013_/X _33045_/Q _25209_/S VGND VGND VPWR VPWR _25206_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22417_ _34815_/Q _34751_/Q _34687_/Q _34623_/Q _22241_/X _22242_/X VGND VGND VPWR
+ VPWR _22417_/X sky130_fd_sc_hd__mux4_1
X_26185_ _25050_/X _33505_/Q _26185_/S VGND VGND VPWR VPWR _26186_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23397_ _32257_/Q _23307_/X _23413_/S VGND VGND VPWR VPWR _23398_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25136_ _25136_/A VGND VGND VPWR VPWR _33020_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22348_ _34557_/Q _32445_/Q _34429_/Q _34365_/Q _22178_/X _22179_/X VGND VGND VPWR
+ VPWR _22348_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29944_ _35223_/Q _29079_/X _29944_/S VGND VGND VPWR VPWR _29945_/A sky130_fd_sc_hd__mux2_1
X_25067_ _25066_/X _32998_/Q _25082_/S VGND VGND VPWR VPWR _25068_/A sky130_fd_sc_hd__mux2_1
X_22279_ _35067_/Q _35003_/Q _34939_/Q _34875_/Q _22109_/X _22110_/X VGND VGND VPWR
+ VPWR _22279_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24018_ _24018_/A VGND VGND VPWR VPWR _32546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29875_ _35190_/Q _29175_/X _29893_/S VGND VGND VPWR VPWR _29876_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16840_ _16840_/A _16840_/B _16840_/C _16840_/D VGND VGND VPWR VPWR _16841_/A sky130_fd_sc_hd__or4_4
X_28826_ _26891_/X _34724_/Q _28840_/S VGND VGND VPWR VPWR _28827_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16771_ _17830_/A VGND VGND VPWR VPWR _16771_/X sky130_fd_sc_hd__clkbuf_4
X_28757_ _28757_/A VGND VGND VPWR VPWR _34691_/D sky130_fd_sc_hd__clkbuf_1
X_25969_ _25969_/A VGND VGND VPWR VPWR _33402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18510_ _34002_/Q _33938_/Q _33874_/Q _32146_/Q _18408_/X _18409_/X VGND VGND VPWR
+ VPWR _18510_/X sky130_fd_sc_hd__mux4_1
X_27708_ _34194_/Q _24258_/X _27718_/S VGND VGND VPWR VPWR _27709_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19490_ _35053_/Q _34989_/Q _34925_/Q _34861_/Q _19456_/X _19457_/X VGND VGND VPWR
+ VPWR _19490_/X sky130_fd_sc_hd__mux4_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28688_ _28688_/A VGND VGND VPWR VPWR _34658_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18441_ _20158_/A VGND VGND VPWR VPWR _18441_/X sky130_fd_sc_hd__buf_4
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27639_ _27639_/A VGND VGND VPWR VPWR _34161_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _18355_/X _18369_/X _18371_/X VGND VGND VPWR VPWR _18402_/C sky130_fd_sc_hd__o21ba_1
XFILLER_178_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30650_ _35557_/Q _29123_/X _30662_/S VGND VGND VPWR VPWR _30651_/A sky130_fd_sc_hd__mux2_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _35313_/Q _35249_/Q _35185_/Q _32305_/Q _17006_/X _17007_/X VGND VGND VPWR
+ VPWR _17323_/X sky130_fd_sc_hd__mux4_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29309_ _23231_/X _34922_/Q _29311_/S VGND VGND VPWR VPWR _29310_/A sky130_fd_sc_hd__mux2_1
X_30581_ _30581_/A VGND VGND VPWR VPWR _35524_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32320_ _32967_/CLK _32320_/D VGND VGND VPWR VPWR _32320_/Q sky130_fd_sc_hd__dfxtp_1
X_17254_ _16999_/X _17252_/X _17253_/X _17002_/X VGND VGND VPWR VPWR _17254_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16205_ _16205_/A VGND VGND VPWR VPWR _31953_/D sky130_fd_sc_hd__clkbuf_1
X_32251_ _34171_/CLK _32251_/D VGND VGND VPWR VPWR _32251_/Q sky130_fd_sc_hd__dfxtp_1
X_17185_ _17181_/X _17184_/X _17147_/X VGND VGND VPWR VPWR _17193_/C sky130_fd_sc_hd__o21ba_1
XFILLER_31_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31202_ _35819_/Q input22/X _31202_/S VGND VGND VPWR VPWR _31203_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16136_ _17855_/A VGND VGND VPWR VPWR _16136_/X sky130_fd_sc_hd__buf_4
XFILLER_31_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32182_ _36134_/CLK _32182_/D VGND VGND VPWR VPWR _32182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31133_ _31133_/A VGND VGND VPWR VPWR _35786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16067_ _17773_/A VGND VGND VPWR VPWR _17865_/A sky130_fd_sc_hd__buf_12
XFILLER_29_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31064_ _31064_/A VGND VGND VPWR VPWR _35753_/D sky130_fd_sc_hd__clkbuf_1
X_35941_ _35941_/CLK _35941_/D VGND VGND VPWR VPWR _35941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30015_ _30015_/A VGND VGND VPWR VPWR _35256_/D sky130_fd_sc_hd__clkbuf_1
X_19826_ _33271_/Q _36151_/Q _33143_/Q _33079_/Q _19711_/X _19712_/X VGND VGND VPWR
+ VPWR _19826_/X sky130_fd_sc_hd__mux4_1
XFILLER_233_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35872_ _35940_/CLK _35872_/D VGND VGND VPWR VPWR _35872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34823_ _35080_/CLK _34823_/D VGND VGND VPWR VPWR _34823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19757_ _35829_/Q _32207_/Q _35701_/Q _35637_/Q _19613_/X _19614_/X VGND VGND VPWR
+ VPWR _19757_/X sky130_fd_sc_hd__mux4_1
X_16969_ _34791_/Q _34727_/Q _34663_/Q _34599_/Q _16935_/X _16936_/X VGND VGND VPWR
+ VPWR _16969_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18708_ _34519_/Q _32407_/Q _34391_/Q _34327_/Q _18466_/X _18467_/X VGND VGND VPWR
+ VPWR _18708_/X sky130_fd_sc_hd__mux4_1
X_34754_ _34819_/CLK _34754_/D VGND VGND VPWR VPWR _34754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31966_ _35166_/CLK _31966_/D VGND VGND VPWR VPWR _31966_/Q sky130_fd_sc_hd__dfxtp_1
X_19688_ _35571_/Q _35507_/Q _35443_/Q _35379_/Q _19550_/X _19551_/X VGND VGND VPWR
+ VPWR _19688_/X sky130_fd_sc_hd__mux4_1
X_33705_ _34281_/CLK _33705_/D VGND VGND VPWR VPWR _33705_/Q sky130_fd_sc_hd__dfxtp_1
X_18639_ _18635_/X _18638_/X _18400_/X VGND VGND VPWR VPWR _18640_/D sky130_fd_sc_hd__o21ba_1
X_30917_ _30917_/A VGND VGND VPWR VPWR _35683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_227_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34685_ _35965_/CLK _34685_/D VGND VGND VPWR VPWR _34685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31897_ _31897_/A VGND VGND VPWR VPWR _36148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33636_ _34276_/CLK _33636_/D VGND VGND VPWR VPWR _33636_/Q sky130_fd_sc_hd__dfxtp_1
X_21650_ _21442_/X _21648_/X _21649_/X _21447_/X VGND VGND VPWR VPWR _21650_/X sky130_fd_sc_hd__a22o_1
X_30848_ _23313_/X _35651_/Q _30860_/S VGND VGND VPWR VPWR _30849_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20601_ input74/X input73/X VGND VGND VPWR VPWR _22373_/A sky130_fd_sc_hd__nor2b_4
XFILLER_33_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21581_ _33512_/Q _33448_/Q _33384_/Q _33320_/Q _21370_/X _21371_/X VGND VGND VPWR
+ VPWR _21581_/X sky130_fd_sc_hd__mux4_1
X_33567_ _34016_/CLK _33567_/D VGND VGND VPWR VPWR _33567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30779_ _23148_/X _35618_/Q _30797_/S VGND VGND VPWR VPWR _30780_/A sky130_fd_sc_hd__mux2_1
X_23320_ _32224_/Q _23319_/X _23334_/S VGND VGND VPWR VPWR _23321_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35306_ _36011_/CLK _35306_/D VGND VGND VPWR VPWR _35306_/Q sky130_fd_sc_hd__dfxtp_1
X_32518_ _32518_/CLK _32518_/D VGND VGND VPWR VPWR _32518_/Q sky130_fd_sc_hd__dfxtp_1
X_20532_ _35596_/Q _35532_/Q _35468_/Q _35404_/Q _20256_/X _20257_/X VGND VGND VPWR
+ VPWR _20532_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_1187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33498_ _34202_/CLK _33498_/D VGND VGND VPWR VPWR _33498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20463_ _33290_/Q _36170_/Q _33162_/Q _33098_/Q _18328_/X _19457_/A VGND VGND VPWR
+ VPWR _20463_/X sky130_fd_sc_hd__mux4_1
X_23251_ _32201_/Q _23250_/X _23268_/S VGND VGND VPWR VPWR _23252_/A sky130_fd_sc_hd__mux2_1
X_35237_ _36004_/CLK _35237_/D VGND VGND VPWR VPWR _35237_/Q sky130_fd_sc_hd__dfxtp_1
X_32449_ _32518_/CLK _32449_/D VGND VGND VPWR VPWR _32449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22202_ _21947_/X _22200_/X _22201_/X _21950_/X VGND VGND VPWR VPWR _22202_/X sky130_fd_sc_hd__a22o_1
X_20394_ _20394_/A VGND VGND VPWR VPWR _32135_/D sky130_fd_sc_hd__buf_4
XFILLER_174_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23182_ _32174_/Q _23114_/X _23182_/S VGND VGND VPWR VPWR _23183_/A sky130_fd_sc_hd__mux2_1
X_35168_ _35294_/CLK _35168_/D VGND VGND VPWR VPWR _35168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34119_ _34819_/CLK _34119_/D VGND VGND VPWR VPWR _34119_/Q sky130_fd_sc_hd__dfxtp_1
X_22133_ _35767_/Q _35127_/Q _34487_/Q _33847_/Q _22093_/X _22094_/X VGND VGND VPWR
+ VPWR _22133_/X sky130_fd_sc_hd__mux4_1
XFILLER_238_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27990_ _28101_/S VGND VGND VPWR VPWR _28009_/S sky130_fd_sc_hd__buf_6
Xoutput240 _32080_/Q VGND VGND VPWR VPWR D3[2] sky130_fd_sc_hd__buf_2
X_35099_ _35933_/CLK _35099_/D VGND VGND VPWR VPWR _35099_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput251 _32081_/Q VGND VGND VPWR VPWR D3[3] sky130_fd_sc_hd__buf_2
XTAP_6617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput262 _32082_/Q VGND VGND VPWR VPWR D3[4] sky130_fd_sc_hd__buf_2
XFILLER_47_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26941_ _26940_/X _33844_/Q _26944_/S VGND VGND VPWR VPWR _26942_/A sky130_fd_sc_hd__mux2_1
XTAP_6639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput273 _32083_/Q VGND VGND VPWR VPWR D3[5] sky130_fd_sc_hd__buf_2
X_22064_ _34805_/Q _34741_/Q _34677_/Q _34613_/Q _21888_/X _21889_/X VGND VGND VPWR
+ VPWR _22064_/X sky130_fd_sc_hd__mux4_1
XTAP_5905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21015_ _34264_/Q _34200_/Q _34136_/Q _34072_/Q _20983_/X _20984_/X VGND VGND VPWR
+ VPWR _21015_/X sky130_fd_sc_hd__mux4_1
XFILLER_87_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29660_ _35088_/Q _29058_/X _29674_/S VGND VGND VPWR VPWR _29661_/A sky130_fd_sc_hd__mux2_1
XTAP_5938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26872_ input8/X VGND VGND VPWR VPWR _26872_/X sky130_fd_sc_hd__buf_4
XTAP_5949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28611_ _28611_/A VGND VGND VPWR VPWR _34622_/D sky130_fd_sc_hd__clkbuf_1
X_25823_ _25823_/A VGND VGND VPWR VPWR _33333_/D sky130_fd_sc_hd__clkbuf_1
X_29591_ _29591_/A VGND VGND VPWR VPWR _35055_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_214_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25754_ _25754_/A VGND VGND VPWR VPWR _33300_/D sky130_fd_sc_hd__clkbuf_1
X_28542_ _28542_/A VGND VGND VPWR VPWR _34589_/D sky130_fd_sc_hd__clkbuf_1
X_22966_ input21/X VGND VGND VPWR VPWR _22966_/X sky130_fd_sc_hd__buf_2
XFILLER_28_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24705_ _23059_/X _32840_/Q _24707_/S VGND VGND VPWR VPWR _24706_/A sky130_fd_sc_hd__mux2_1
X_28473_ _26968_/X _34557_/Q _28477_/S VGND VGND VPWR VPWR _28474_/A sky130_fd_sc_hd__mux2_1
X_21917_ _21594_/X _21915_/X _21916_/X _21597_/X VGND VGND VPWR VPWR _21917_/X sky130_fd_sc_hd__a22o_1
X_25685_ _33269_/Q _24366_/X _25685_/S VGND VGND VPWR VPWR _25686_/A sky130_fd_sc_hd__mux2_1
X_22897_ _22897_/A VGND VGND VPWR VPWR _32019_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27424_ _34061_/Q _24440_/X _27424_/S VGND VGND VPWR VPWR _27425_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24636_ _22957_/X _32807_/Q _24644_/S VGND VGND VPWR VPWR _24637_/A sky130_fd_sc_hd__mux2_1
XFILLER_230_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21848_ _35759_/Q _35119_/Q _34479_/Q _33839_/Q _21740_/X _21741_/X VGND VGND VPWR
+ VPWR _21848_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27355_ _27424_/S VGND VGND VPWR VPWR _27374_/S sky130_fd_sc_hd__buf_4
X_24567_ _23059_/X _32776_/Q _24569_/S VGND VGND VPWR VPWR _24568_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21779_ _35821_/Q _32198_/Q _35693_/Q _35629_/Q _21560_/X _21561_/X VGND VGND VPWR
+ VPWR _21779_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26306_ _25029_/X _33562_/Q _26320_/S VGND VGND VPWR VPWR _26307_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23518_ _23013_/X _32313_/Q _23530_/S VGND VGND VPWR VPWR _23519_/A sky130_fd_sc_hd__mux2_1
X_27286_ _27286_/A VGND VGND VPWR VPWR _33995_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24498_ _22957_/X _32743_/Q _24506_/S VGND VGND VPWR VPWR _24499_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29025_ _29025_/A VGND VGND VPWR VPWR _34818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26237_ _26237_/A VGND VGND VPWR VPWR _33529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23449_ _22910_/X _32280_/Q _23467_/S VGND VGND VPWR VPWR _23450_/A sky130_fd_sc_hd__mux2_1
XFILLER_221_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26168_ _26168_/A VGND VGND VPWR VPWR _33496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25119_ input36/X VGND VGND VPWR VPWR _25119_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_152_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26099_ _25122_/X _33464_/Q _26113_/S VGND VGND VPWR VPWR _26100_/A sky130_fd_sc_hd__mux2_1
X_18990_ _35039_/Q _34975_/Q _34911_/Q _34847_/Q _18750_/X _18751_/X VGND VGND VPWR
+ VPWR _18990_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ _17901_/X _17939_/X _17940_/X _17906_/X VGND VGND VPWR VPWR _17941_/X sky130_fd_sc_hd__a22o_1
X_29927_ _29927_/A VGND VGND VPWR VPWR _35214_/D sky130_fd_sc_hd__clkbuf_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17872_ _34305_/Q _34241_/Q _34177_/Q _34113_/Q _17795_/X _17796_/X VGND VGND VPWR
+ VPWR _17872_/X sky130_fd_sc_hd__mux4_1
X_29858_ _35182_/Q _29151_/X _29872_/S VGND VGND VPWR VPWR _29859_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19611_ _19363_/X _19609_/X _19610_/X _19367_/X VGND VGND VPWR VPWR _19611_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28809_ _26866_/X _34716_/Q _28819_/S VGND VGND VPWR VPWR _28810_/A sky130_fd_sc_hd__mux2_1
X_16823_ _32995_/Q _32931_/Q _32867_/Q _32803_/Q _16636_/X _16637_/X VGND VGND VPWR
+ VPWR _16823_/X sky130_fd_sc_hd__mux4_1
X_29789_ _30059_/A _30870_/B VGND VGND VPWR VPWR _29922_/S sky130_fd_sc_hd__nor2_8
X_31820_ _31820_/A VGND VGND VPWR VPWR _36111_/D sky130_fd_sc_hd__clkbuf_1
X_19542_ _19355_/X _19540_/X _19541_/X _19361_/X VGND VGND VPWR VPWR _19542_/X sky130_fd_sc_hd__a22o_1
XFILLER_19_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16754_ _35553_/Q _35489_/Q _35425_/Q _35361_/Q _16544_/X _16545_/X VGND VGND VPWR
+ VPWR _16754_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19473_ _33261_/Q _36141_/Q _33133_/Q _33069_/Q _19358_/X _19359_/X VGND VGND VPWR
+ VPWR _19473_/X sky130_fd_sc_hd__mux4_1
X_16685_ _16681_/X _16684_/X _16441_/X VGND VGND VPWR VPWR _16693_/C sky130_fd_sc_hd__o21ba_1
X_31751_ _36079_/Q input27/X _31763_/S VGND VGND VPWR VPWR _31752_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18424_ _33167_/Q _32527_/Q _35919_/Q _35855_/Q _18363_/X _18365_/X VGND VGND VPWR
+ VPWR _18424_/X sky130_fd_sc_hd__mux4_1
X_30702_ _35582_/Q _29200_/X _30704_/S VGND VGND VPWR VPWR _30703_/A sky130_fd_sc_hd__mux2_1
XFILLER_234_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34470_ _35749_/CLK _34470_/D VGND VGND VPWR VPWR _34470_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31682_ _36046_/Q input1/X _31700_/S VGND VGND VPWR VPWR _31683_/A sky130_fd_sc_hd__mux2_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33421_ _34060_/CLK _33421_/D VGND VGND VPWR VPWR _33421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18355_ _18344_/X _18347_/X _18352_/X _18354_/X VGND VGND VPWR VPWR _18355_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30633_ _35549_/Q _29098_/X _30641_/S VGND VGND VPWR VPWR _30634_/A sky130_fd_sc_hd__mux2_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17306_ _32753_/Q _32689_/Q _32625_/Q _36081_/Q _17272_/X _17056_/X VGND VGND VPWR
+ VPWR _17306_/X sky130_fd_sc_hd__mux4_1
X_36140_ _36141_/CLK _36140_/D VGND VGND VPWR VPWR _36140_/Q sky130_fd_sc_hd__dfxtp_1
X_33352_ _34306_/CLK _33352_/D VGND VGND VPWR VPWR _33352_/Q sky130_fd_sc_hd__dfxtp_1
X_30564_ _30564_/A VGND VGND VPWR VPWR _35516_/D sky130_fd_sc_hd__clkbuf_1
X_18286_ _20067_/A VGND VGND VPWR VPWR _20206_/A sky130_fd_sc_hd__buf_12
XFILLER_174_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32303_ _35564_/CLK _32303_/D VGND VGND VPWR VPWR _32303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17237_ _34031_/Q _33967_/Q _33903_/Q _32239_/Q _17020_/X _17021_/X VGND VGND VPWR
+ VPWR _17237_/X sky130_fd_sc_hd__mux4_1
X_36071_ _36072_/CLK _36071_/D VGND VGND VPWR VPWR _36071_/Q sky130_fd_sc_hd__dfxtp_1
X_33283_ _36165_/CLK _33283_/D VGND VGND VPWR VPWR _33283_/Q sky130_fd_sc_hd__dfxtp_1
X_30495_ _30495_/A VGND VGND VPWR VPWR _35483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1043 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35022_ _35729_/CLK _35022_/D VGND VGND VPWR VPWR _35022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_970 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32234_ _36139_/CLK _32234_/D VGND VGND VPWR VPWR _32234_/Q sky130_fd_sc_hd__dfxtp_1
X_17168_ _33517_/Q _33453_/Q _33389_/Q _33325_/Q _17123_/X _17124_/X VGND VGND VPWR
+ VPWR _17168_/X sky130_fd_sc_hd__mux4_2
XFILLER_155_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16119_ _16115_/X _16118_/X _16040_/X _16042_/X VGND VGND VPWR VPWR _16134_/B sky130_fd_sc_hd__o211a_1
XFILLER_115_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32165_ _35792_/CLK _32165_/D VGND VGND VPWR VPWR _32165_/Q sky130_fd_sc_hd__dfxtp_1
X_17099_ _17055_/X _17097_/X _17098_/X _17061_/X VGND VGND VPWR VPWR _17099_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31116_ _35778_/Q _29213_/X _31130_/S VGND VGND VPWR VPWR _31117_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32096_ _35807_/CLK _32096_/D VGND VGND VPWR VPWR _32096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35924_ _35927_/CLK _35924_/D VGND VGND VPWR VPWR _35924_/Q sky130_fd_sc_hd__dfxtp_1
X_31047_ _31047_/A VGND VGND VPWR VPWR _35745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19809_ _20162_/A VGND VGND VPWR VPWR _19809_/X sky130_fd_sc_hd__buf_4
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35855_ _35917_/CLK _35855_/D VGND VGND VPWR VPWR _35855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22820_ _20626_/X _22818_/X _22819_/X _20637_/X VGND VGND VPWR VPWR _22820_/X sky130_fd_sc_hd__a22o_1
X_34806_ _35575_/CLK _34806_/D VGND VGND VPWR VPWR _34806_/Q sky130_fd_sc_hd__dfxtp_1
X_35786_ _35788_/CLK _35786_/D VGND VGND VPWR VPWR _35786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32998_ _36070_/CLK _32998_/D VGND VGND VPWR VPWR _32998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22751_ _22460_/X _22749_/X _22750_/X _22465_/X VGND VGND VPWR VPWR _22751_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34737_ _34932_/CLK _34737_/D VGND VGND VPWR VPWR _34737_/Q sky130_fd_sc_hd__dfxtp_1
X_31949_ _31949_/A VGND VGND VPWR VPWR _36173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21702_ _21663_/X _21700_/X _21701_/X _21667_/X VGND VGND VPWR VPWR _21702_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25470_ _33168_/Q _24252_/X _25484_/S VGND VGND VPWR VPWR _25471_/A sky130_fd_sc_hd__mux2_1
X_22682_ _35591_/Q _35527_/Q _35463_/Q _35399_/Q _22556_/X _22557_/X VGND VGND VPWR
+ VPWR _22682_/X sky130_fd_sc_hd__mux4_1
X_34668_ _35304_/CLK _34668_/D VGND VGND VPWR VPWR _34668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24421_ _24421_/A VGND VGND VPWR VPWR _32710_/D sky130_fd_sc_hd__clkbuf_1
X_33619_ _33685_/CLK _33619_/D VGND VGND VPWR VPWR _33619_/Q sky130_fd_sc_hd__dfxtp_1
X_21633_ _35753_/Q _35113_/Q _34473_/Q _33833_/Q _21387_/X _21388_/X VGND VGND VPWR
+ VPWR _21633_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34599_ _36005_/CLK _34599_/D VGND VGND VPWR VPWR _34599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27140_ _26996_/X _33926_/Q _27146_/S VGND VGND VPWR VPWR _27141_/A sky130_fd_sc_hd__mux2_1
X_24352_ _32688_/Q _24351_/X _24367_/S VGND VGND VPWR VPWR _24353_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21564_ _21241_/X _21562_/X _21563_/X _21244_/X VGND VGND VPWR VPWR _21564_/X sky130_fd_sc_hd__a22o_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23303_ input46/X VGND VGND VPWR VPWR _23303_/X sky130_fd_sc_hd__buf_4
X_20515_ _33804_/Q _33740_/Q _33676_/Q _33612_/Q _18320_/X _18321_/X VGND VGND VPWR
+ VPWR _20515_/X sky130_fd_sc_hd__mux4_1
X_27071_ _26894_/X _33893_/Q _27083_/S VGND VGND VPWR VPWR _27072_/A sky130_fd_sc_hd__mux2_1
X_24283_ input4/X VGND VGND VPWR VPWR _24283_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_165_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21495_ _35749_/Q _35109_/Q _34469_/Q _33829_/Q _21387_/X _21388_/X VGND VGND VPWR
+ VPWR _21495_/X sky130_fd_sc_hd__mux4_1
X_26022_ _26022_/A VGND VGND VPWR VPWR _33427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23234_ input22/X VGND VGND VPWR VPWR _23234_/X sky130_fd_sc_hd__buf_4
XFILLER_101_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20446_ _34825_/Q _34761_/Q _34697_/Q _34633_/Q _20294_/X _20295_/X VGND VGND VPWR
+ VPWR _20446_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1022 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23165_ _32166_/Q _23093_/X _23182_/S VGND VGND VPWR VPWR _23166_/A sky130_fd_sc_hd__mux2_1
XTAP_7126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20377_ _20069_/X _20375_/X _20376_/X _20073_/X VGND VGND VPWR VPWR _20377_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22116_ _22116_/A _22116_/B _22116_/C _22116_/D VGND VGND VPWR VPWR _22117_/A sky130_fd_sc_hd__or4_4
XTAP_6414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27973_ _27973_/A VGND VGND VPWR VPWR _34319_/D sky130_fd_sc_hd__clkbuf_1
X_23096_ input34/X VGND VGND VPWR VPWR _23096_/X sky130_fd_sc_hd__buf_4
XANTENNA_1209 _23274_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29712_ _35113_/Q _29135_/X _29716_/S VGND VGND VPWR VPWR _29713_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26924_ _26924_/A VGND VGND VPWR VPWR _33838_/D sky130_fd_sc_hd__clkbuf_1
X_22047_ _34037_/Q _33973_/Q _33909_/Q _32245_/Q _21973_/X _21974_/X VGND VGND VPWR
+ VPWR _22047_/X sky130_fd_sc_hd__mux4_1
XFILLER_248_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29643_ _29643_/A VGND VGND VPWR VPWR _35080_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26855_ _26853_/X _33816_/Q _26882_/S VGND VGND VPWR VPWR _26856_/A sky130_fd_sc_hd__mux2_1
XTAP_5779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25806_ _25088_/X _33325_/Q _25822_/S VGND VGND VPWR VPWR _25807_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26786_ _33789_/Q _24391_/X _26790_/S VGND VGND VPWR VPWR _26787_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29574_ _29574_/A VGND VGND VPWR VPWR _35047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_235_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23998_ _22914_/X _32537_/Q _24014_/S VGND VGND VPWR VPWR _23999_/A sky130_fd_sc_hd__mux2_1
XFILLER_217_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25737_ input87/X _29049_/B input88/X VGND VGND VPWR VPWR _25738_/A sky130_fd_sc_hd__and3b_1
X_28525_ _28525_/A VGND VGND VPWR VPWR _34581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22949_ _22948_/X _32036_/Q _22970_/S VGND VGND VPWR VPWR _22950_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16470_ _32985_/Q _32921_/Q _32857_/Q _32793_/Q _16283_/X _16284_/X VGND VGND VPWR
+ VPWR _16470_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25668_ _25668_/A VGND VGND VPWR VPWR _33260_/D sky130_fd_sc_hd__clkbuf_1
X_28456_ _26943_/X _34549_/Q _28456_/S VGND VGND VPWR VPWR _28457_/A sky130_fd_sc_hd__mux2_1
XFILLER_243_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27407_ _27407_/A VGND VGND VPWR VPWR _34052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24619_ _22932_/X _32799_/Q _24623_/S VGND VGND VPWR VPWR _24620_/A sky130_fd_sc_hd__mux2_1
X_28387_ _26841_/X _34516_/Q _28393_/S VGND VGND VPWR VPWR _28388_/A sky130_fd_sc_hd__mux2_1
X_25599_ _31815_/B VGND VGND VPWR VPWR _25602_/A sky130_fd_sc_hd__inv_2
XFILLER_106_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18140_ _35785_/Q _35145_/Q _34505_/Q _33865_/Q _17846_/X _17847_/X VGND VGND VPWR
+ VPWR _18140_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27338_ _27338_/A VGND VGND VPWR VPWR _34019_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18071_ _18067_/X _18070_/X _17834_/X VGND VGND VPWR VPWR _18093_/A sky130_fd_sc_hd__o21ba_2
XFILLER_12_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27269_ _26987_/X _33987_/Q _27281_/S VGND VGND VPWR VPWR _27270_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17022_ _34025_/Q _33961_/Q _33897_/Q _32226_/Q _17020_/X _17021_/X VGND VGND VPWR
+ VPWR _17022_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29008_ _29008_/A VGND VGND VPWR VPWR _34810_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30280_ _35382_/Q _29175_/X _30298_/S VGND VGND VPWR VPWR _30281_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18973_ _33247_/Q _36127_/Q _33119_/Q _33055_/Q _18652_/X _18653_/X VGND VGND VPWR
+ VPWR _18973_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17924_ _35586_/Q _35522_/Q _35458_/Q _35394_/Q _17603_/X _17604_/X VGND VGND VPWR
+ VPWR _17924_/X sky130_fd_sc_hd__mux4_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33970_ _34222_/CLK _33970_/D VGND VGND VPWR VPWR _33970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32921_ _36055_/CLK _32921_/D VGND VGND VPWR VPWR _32921_/Q sky130_fd_sc_hd__dfxtp_1
X_17855_ _17855_/A VGND VGND VPWR VPWR _17855_/X sky130_fd_sc_hd__buf_4
XFILLER_67_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35640_ _35766_/CLK _35640_/D VGND VGND VPWR VPWR _35640_/Q sky130_fd_sc_hd__dfxtp_1
X_16806_ _17159_/A VGND VGND VPWR VPWR _16806_/X sky130_fd_sc_hd__clkbuf_4
X_32852_ _35991_/CLK _32852_/D VGND VGND VPWR VPWR _32852_/Q sky130_fd_sc_hd__dfxtp_1
X_17786_ _35326_/Q _35262_/Q _35198_/Q _32318_/Q _17712_/X _17713_/X VGND VGND VPWR
+ VPWR _17786_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31803_ _36104_/Q input54/X _31805_/S VGND VGND VPWR VPWR _31804_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19525_ _20231_/A VGND VGND VPWR VPWR _19525_/X sky130_fd_sc_hd__buf_6
X_35571_ _36019_/CLK _35571_/D VGND VGND VPWR VPWR _35571_/Q sky130_fd_sc_hd__dfxtp_1
X_16737_ _17957_/A VGND VGND VPWR VPWR _16737_/X sky130_fd_sc_hd__buf_4
X_32783_ _35985_/CLK _32783_/D VGND VGND VPWR VPWR _32783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34522_ _34970_/CLK _34522_/D VGND VGND VPWR VPWR _34522_/Q sky130_fd_sc_hd__dfxtp_1
X_19456_ _20162_/A VGND VGND VPWR VPWR _19456_/X sky130_fd_sc_hd__buf_4
X_31734_ _36071_/Q input18/X _31742_/S VGND VGND VPWR VPWR _31735_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16668_ _17847_/A VGND VGND VPWR VPWR _16668_/X sky130_fd_sc_hd__buf_4
XFILLER_201_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18407_ _33487_/Q _33423_/Q _33359_/Q _33295_/Q _18298_/X _18299_/X VGND VGND VPWR
+ VPWR _18407_/X sky130_fd_sc_hd__mux4_2
X_34453_ _35730_/CLK _34453_/D VGND VGND VPWR VPWR _34453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31665_ _31665_/A VGND VGND VPWR VPWR _36038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19387_ _19387_/A VGND VGND VPWR VPWR _32106_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16599_ _16595_/X _16598_/X _16422_/X VGND VGND VPWR VPWR _16623_/A sky130_fd_sc_hd__o21ba_1
X_33404_ _33723_/CLK _33404_/D VGND VGND VPWR VPWR _33404_/Q sky130_fd_sc_hd__dfxtp_1
X_18338_ _18326_/X _18331_/X _18336_/X _18337_/X VGND VGND VPWR VPWR _18338_/X sky130_fd_sc_hd__a22o_1
X_30616_ _35541_/Q _29073_/X _30620_/S VGND VGND VPWR VPWR _30617_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34384_ _36211_/CLK _34384_/D VGND VGND VPWR VPWR _34384_/Q sky130_fd_sc_hd__dfxtp_1
X_31596_ _31596_/A VGND VGND VPWR VPWR _36005_/D sky130_fd_sc_hd__clkbuf_1
X_36123_ _36123_/CLK _36123_/D VGND VGND VPWR VPWR _36123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33335_ _34039_/CLK _33335_/D VGND VGND VPWR VPWR _33335_/Q sky130_fd_sc_hd__dfxtp_1
X_18269_ _34573_/Q _32461_/Q _34445_/Q _34381_/Q _16063_/X _16065_/X VGND VGND VPWR
+ VPWR _18269_/X sky130_fd_sc_hd__mux4_1
X_30547_ _30547_/A VGND VGND VPWR VPWR _35508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20300_ _35076_/Q _35012_/Q _34948_/Q _34884_/Q _20162_/X _20163_/X VGND VGND VPWR
+ VPWR _20300_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36054_ _36055_/CLK _36054_/D VGND VGND VPWR VPWR _36054_/Q sky130_fd_sc_hd__dfxtp_1
X_21280_ _35743_/Q _35103_/Q _34463_/Q _33823_/Q _21034_/X _21035_/X VGND VGND VPWR
+ VPWR _21280_/X sky130_fd_sc_hd__mux4_1
X_33266_ _33520_/CLK _33266_/D VGND VGND VPWR VPWR _33266_/Q sky130_fd_sc_hd__dfxtp_1
X_30478_ _30478_/A VGND VGND VPWR VPWR _35475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35005_ _35989_/CLK _35005_/D VGND VGND VPWR VPWR _35005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20231_ _20231_/A VGND VGND VPWR VPWR _20231_/X sky130_fd_sc_hd__buf_6
X_32217_ _35968_/CLK _32217_/D VGND VGND VPWR VPWR _32217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33197_ _35885_/CLK _33197_/D VGND VGND VPWR VPWR _33197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20162_ _20162_/A VGND VGND VPWR VPWR _20162_/X sky130_fd_sc_hd__buf_4
XFILLER_143_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32148_ _34001_/CLK _32148_/D VGND VGND VPWR VPWR _32148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24970_ _24970_/A VGND VGND VPWR VPWR _32964_/D sky130_fd_sc_hd__clkbuf_1
X_20093_ _20093_/A VGND VGND VPWR VPWR _32126_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_48_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32079_ _34973_/CLK _32079_/D VGND VGND VPWR VPWR _32079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23921_ _23921_/A VGND VGND VPWR VPWR _32501_/D sky130_fd_sc_hd__clkbuf_1
X_35907_ _35971_/CLK _35907_/D VGND VGND VPWR VPWR _35907_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26640_ _25122_/X _33720_/Q _26654_/S VGND VGND VPWR VPWR _26641_/A sky130_fd_sc_hd__mux2_1
X_35838_ _35903_/CLK _35838_/D VGND VGND VPWR VPWR _35838_/Q sky130_fd_sc_hd__dfxtp_1
X_23852_ _23852_/A VGND VGND VPWR VPWR _32468_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22803_ _33227_/Q _32587_/Q _35979_/Q _35915_/Q _20675_/X _20676_/X VGND VGND VPWR
+ VPWR _22803_/X sky130_fd_sc_hd__mux4_1
XANTENNA_607 _18435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26571_ _26571_/A VGND VGND VPWR VPWR _33687_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_618 _18571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35769_ _35771_/CLK _35769_/D VGND VGND VPWR VPWR _35769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23783_ _23783_/A VGND VGND VPWR VPWR _32436_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20995_ _32983_/Q _32919_/Q _32855_/Q _32791_/Q _20883_/X _20884_/X VGND VGND VPWR
+ VPWR _20995_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_629 _18787_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28310_ _28310_/A VGND VGND VPWR VPWR _34479_/D sky130_fd_sc_hd__clkbuf_1
X_25522_ _33193_/Q _24329_/X _25526_/S VGND VGND VPWR VPWR _25523_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22734_ _21749_/A _22732_/X _22733_/X _21752_/A VGND VGND VPWR VPWR _22734_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_1013 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29290_ _23145_/X _34913_/Q _29290_/S VGND VGND VPWR VPWR _29291_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28241_ _28241_/A VGND VGND VPWR VPWR _34446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25453_ _25453_/A VGND VGND VPWR VPWR _33162_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22665_ _33799_/Q _33735_/Q _33671_/Q _33607_/Q _22502_/X _22503_/X VGND VGND VPWR
+ VPWR _22665_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1079 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24404_ input47/X VGND VGND VPWR VPWR _24404_/X sky130_fd_sc_hd__buf_6
X_21616_ _33769_/Q _33705_/Q _33641_/Q _33577_/Q _21443_/X _21444_/X VGND VGND VPWR
+ VPWR _21616_/X sky130_fd_sc_hd__mux4_1
X_28172_ _26922_/X _34414_/Q _28186_/S VGND VGND VPWR VPWR _28173_/A sky130_fd_sc_hd__mux2_1
X_25384_ _25384_/A VGND VGND VPWR VPWR _33129_/D sky130_fd_sc_hd__clkbuf_1
X_22596_ _34820_/Q _34756_/Q _34692_/Q _34628_/Q _22594_/X _22595_/X VGND VGND VPWR
+ VPWR _22596_/X sky130_fd_sc_hd__mux4_1
XFILLER_205_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27123_ _26971_/X _33918_/Q _27125_/S VGND VGND VPWR VPWR _27124_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24335_ input22/X VGND VGND VPWR VPWR _24335_/X sky130_fd_sc_hd__buf_4
XFILLER_103_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21547_ _34279_/Q _34215_/Q _34151_/Q _34087_/Q _21336_/X _21337_/X VGND VGND VPWR
+ VPWR _21547_/X sky130_fd_sc_hd__mux4_1
X_27054_ _26869_/X _33885_/Q _27062_/S VGND VGND VPWR VPWR _27055_/A sky130_fd_sc_hd__mux2_1
X_24266_ _24266_/A VGND VGND VPWR VPWR _32660_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21478_ _21478_/A _21478_/B _21478_/C _21478_/D VGND VGND VPWR VPWR _21479_/A sky130_fd_sc_hd__or4_4
X_26005_ _25183_/X _33420_/Q _26007_/S VGND VGND VPWR VPWR _26006_/A sky130_fd_sc_hd__mux2_1
X_23217_ input17/X VGND VGND VPWR VPWR _23217_/X sky130_fd_sc_hd__clkbuf_4
X_20429_ _34057_/Q _33993_/Q _33929_/Q _32265_/Q _18358_/X _18360_/X VGND VGND VPWR
+ VPWR _20429_/X sky130_fd_sc_hd__mux4_1
X_24197_ _23007_/X _32631_/Q _24213_/S VGND VGND VPWR VPWR _24198_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23148_ input13/X VGND VGND VPWR VPWR _23148_/X sky130_fd_sc_hd__buf_4
XFILLER_107_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1006 _17862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1017 _17995_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1028 _17865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27956_ _34312_/Q _24425_/X _27958_/S VGND VGND VPWR VPWR _27957_/A sky130_fd_sc_hd__mux2_1
XTAP_6255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23079_ input86/X VGND VGND VPWR VPWR _29049_/B sky130_fd_sc_hd__buf_4
XTAP_5510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1039 _17152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26907_ _26906_/X _33833_/Q _26913_/S VGND VGND VPWR VPWR _26908_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27887_ _34279_/Q _24323_/X _27895_/S VGND VGND VPWR VPWR _27888_/A sky130_fd_sc_hd__mux2_1
XTAP_5576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29626_ _35072_/Q _29206_/X _29644_/S VGND VGND VPWR VPWR _29627_/A sky130_fd_sc_hd__mux2_1
XTAP_4853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ _17636_/X _17639_/X _17500_/X VGND VGND VPWR VPWR _17650_/C sky130_fd_sc_hd__o21ba_1
XTAP_5598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26838_ input56/X VGND VGND VPWR VPWR _26838_/X sky130_fd_sc_hd__buf_4
XFILLER_75_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29557_ _29557_/A VGND VGND VPWR VPWR _35039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17571_ _35576_/Q _35512_/Q _35448_/Q _35384_/Q _17250_/X _17251_/X VGND VGND VPWR
+ VPWR _17571_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26769_ _33781_/Q _24366_/X _26769_/S VGND VGND VPWR VPWR _26770_/A sky130_fd_sc_hd__mux2_1
X_19310_ _34536_/Q _32424_/Q _34408_/Q _34344_/Q _19172_/X _19173_/X VGND VGND VPWR
+ VPWR _19310_/X sky130_fd_sc_hd__mux4_1
X_28508_ _30735_/B _28778_/B VGND VGND VPWR VPWR _28641_/S sky130_fd_sc_hd__nand2_8
XFILLER_147_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16522_ _35034_/Q _34970_/Q _34906_/Q _34842_/Q _16450_/X _16451_/X VGND VGND VPWR
+ VPWR _16522_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29488_ _23300_/X _35007_/Q _29488_/S VGND VGND VPWR VPWR _29489_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19241_ _35046_/Q _34982_/Q _34918_/Q _34854_/Q _19103_/X _19104_/X VGND VGND VPWR
+ VPWR _19241_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28439_ _28439_/A VGND VGND VPWR VPWR _34540_/D sky130_fd_sc_hd__clkbuf_1
X_16453_ _17159_/A VGND VGND VPWR VPWR _16453_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16384_ _17957_/A VGND VGND VPWR VPWR _16384_/X sky130_fd_sc_hd__buf_4
X_31450_ _31450_/A VGND VGND VPWR VPWR _35936_/D sky130_fd_sc_hd__clkbuf_1
X_19172_ _20012_/A VGND VGND VPWR VPWR _19172_/X sky130_fd_sc_hd__clkbuf_8
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18123_ _18123_/A _18123_/B _18123_/C _18123_/D VGND VGND VPWR VPWR _18124_/A sky130_fd_sc_hd__or4_4
X_30401_ _23247_/X _35439_/Q _30413_/S VGND VGND VPWR VPWR _30402_/A sky130_fd_sc_hd__mux2_1
X_31381_ _31408_/S VGND VGND VPWR VPWR _31400_/S sky130_fd_sc_hd__buf_4
XFILLER_12_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33120_ _34146_/CLK _33120_/D VGND VGND VPWR VPWR _33120_/Q sky130_fd_sc_hd__dfxtp_1
X_18054_ _15997_/X _18052_/X _18053_/X _16003_/X VGND VGND VPWR VPWR _18054_/X sky130_fd_sc_hd__a22o_1
X_30332_ _23077_/X _35406_/Q _30350_/S VGND VGND VPWR VPWR _30333_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_3 _32114_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17005_ _34792_/Q _34728_/Q _34664_/Q _34600_/Q _16935_/X _16936_/X VGND VGND VPWR
+ VPWR _17005_/X sky130_fd_sc_hd__mux4_1
X_33051_ _36123_/CLK _33051_/D VGND VGND VPWR VPWR _33051_/Q sky130_fd_sc_hd__dfxtp_1
X_30263_ _35374_/Q _29151_/X _30277_/S VGND VGND VPWR VPWR _30264_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32002_ _36194_/CLK _32002_/D VGND VGND VPWR VPWR _32002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30194_ _31275_/A _31140_/A VGND VGND VPWR VPWR _30327_/S sky130_fd_sc_hd__nor2_8
XFILLER_112_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18956_ _18743_/X _18952_/X _18955_/X _18746_/X VGND VGND VPWR VPWR _18956_/X sky130_fd_sc_hd__a22o_1
XFILLER_234_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17907_ _17901_/X _17904_/X _17905_/X _17906_/X VGND VGND VPWR VPWR _17907_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33953_ _34145_/CLK _33953_/D VGND VGND VPWR VPWR _33953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18887_ _34524_/Q _32412_/Q _34396_/Q _34332_/Q _18819_/X _18820_/X VGND VGND VPWR
+ VPWR _18887_/X sky130_fd_sc_hd__mux4_1
X_32904_ _36171_/CLK _32904_/D VGND VGND VPWR VPWR _32904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17838_ _17761_/X _17836_/X _17837_/X _17767_/X VGND VGND VPWR VPWR _17838_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33884_ _34205_/CLK _33884_/D VGND VGND VPWR VPWR _33884_/Q sky130_fd_sc_hd__dfxtp_1
X_35623_ _35815_/CLK _35623_/D VGND VGND VPWR VPWR _35623_/Q sky130_fd_sc_hd__dfxtp_1
X_32835_ _32965_/CLK _32835_/D VGND VGND VPWR VPWR _32835_/Q sky130_fd_sc_hd__dfxtp_1
X_17769_ _17769_/A VGND VGND VPWR VPWR _17769_/X sky130_fd_sc_hd__clkbuf_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19508_ _32750_/Q _32686_/Q _32622_/Q _36078_/Q _19219_/X _19356_/X VGND VGND VPWR
+ VPWR _19508_/X sky130_fd_sc_hd__mux4_1
X_35554_ _35555_/CLK _35554_/D VGND VGND VPWR VPWR _35554_/Q sky130_fd_sc_hd__dfxtp_1
X_20780_ _20776_/X _20779_/X _20611_/X VGND VGND VPWR VPWR _20804_/A sky130_fd_sc_hd__o21ba_1
X_32766_ _36097_/CLK _32766_/D VGND VGND VPWR VPWR _32766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34505_ _35845_/CLK _34505_/D VGND VGND VPWR VPWR _34505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19439_ _35820_/Q _32197_/Q _35692_/Q _35628_/Q _19260_/X _19261_/X VGND VGND VPWR
+ VPWR _19439_/X sky130_fd_sc_hd__mux4_1
X_31717_ _36063_/Q input9/X _31721_/S VGND VGND VPWR VPWR _31718_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35485_ _35935_/CLK _35485_/D VGND VGND VPWR VPWR _35485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32697_ _36088_/CLK _32697_/D VGND VGND VPWR VPWR _32697_/Q sky130_fd_sc_hd__dfxtp_1
X_34436_ _35332_/CLK _34436_/D VGND VGND VPWR VPWR _34436_/Q sky130_fd_sc_hd__dfxtp_1
X_22450_ _35584_/Q _35520_/Q _35456_/Q _35392_/Q _22203_/X _22204_/X VGND VGND VPWR
+ VPWR _22450_/X sky130_fd_sc_hd__mux4_1
X_31648_ _31648_/A VGND VGND VPWR VPWR _36030_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21401_ _21754_/A VGND VGND VPWR VPWR _21401_/X sky130_fd_sc_hd__clkbuf_4
X_22381_ _22532_/A VGND VGND VPWR VPWR _22381_/X sky130_fd_sc_hd__buf_4
X_34367_ _35966_/CLK _34367_/D VGND VGND VPWR VPWR _34367_/Q sky130_fd_sc_hd__dfxtp_1
X_31579_ _31579_/A VGND VGND VPWR VPWR _35997_/D sky130_fd_sc_hd__clkbuf_1
X_36106_ _36172_/CLK _36106_/D VGND VGND VPWR VPWR _36106_/Q sky130_fd_sc_hd__dfxtp_1
X_24120_ _24120_/A VGND VGND VPWR VPWR _32594_/D sky130_fd_sc_hd__clkbuf_1
X_33318_ _33702_/CLK _33318_/D VGND VGND VPWR VPWR _33318_/Q sky130_fd_sc_hd__dfxtp_1
X_21332_ _21328_/X _21331_/X _21055_/X VGND VGND VPWR VPWR _21333_/D sky130_fd_sc_hd__o21ba_1
XFILLER_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34298_ _34298_/CLK _34298_/D VGND VGND VPWR VPWR _34298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36037_ _36037_/CLK _36037_/D VGND VGND VPWR VPWR _36037_/Q sky130_fd_sc_hd__dfxtp_1
X_24051_ _24051_/A VGND VGND VPWR VPWR _32562_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33249_ _36128_/CLK _33249_/D VGND VGND VPWR VPWR _33249_/Q sky130_fd_sc_hd__dfxtp_1
X_21263_ _33759_/Q _33695_/Q _33631_/Q _33567_/Q _21090_/X _21091_/X VGND VGND VPWR
+ VPWR _21263_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23002_ _23002_/A VGND VGND VPWR VPWR _32053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20214_ _32770_/Q _32706_/Q _32642_/Q _36098_/Q _19925_/X _20062_/X VGND VGND VPWR
+ VPWR _20214_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap283 _24401_/A VGND VGND VPWR VPWR _24441_/S sky130_fd_sc_hd__buf_8
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21194_ _34269_/Q _34205_/Q _34141_/Q _34077_/Q _20983_/X _20984_/X VGND VGND VPWR
+ VPWR _21194_/X sky130_fd_sc_hd__mux4_1
X_27810_ _27810_/A VGND VGND VPWR VPWR _34242_/D sky130_fd_sc_hd__clkbuf_1
X_20145_ _35840_/Q _32219_/Q _35712_/Q _35648_/Q _19966_/X _19967_/X VGND VGND VPWR
+ VPWR _20145_/X sky130_fd_sc_hd__mux4_1
X_28790_ _26838_/X _34707_/Q _28798_/S VGND VGND VPWR VPWR _28791_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24953_ _24953_/A VGND VGND VPWR VPWR _32956_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27741_ _27831_/S VGND VGND VPWR VPWR _27760_/S sky130_fd_sc_hd__buf_4
X_20076_ _35838_/Q _32217_/Q _35710_/Q _35646_/Q _19966_/X _19967_/X VGND VGND VPWR
+ VPWR _20076_/X sky130_fd_sc_hd__mux4_1
XTAP_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23904_ _22976_/X _32493_/Q _23920_/S VGND VGND VPWR VPWR _23905_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27672_ _34177_/Q _24404_/X _27688_/S VGND VGND VPWR VPWR _27673_/A sky130_fd_sc_hd__mux2_1
X_24884_ _24884_/A VGND VGND VPWR VPWR _32923_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29411_ _23124_/X _34970_/Q _29425_/S VGND VGND VPWR VPWR _29412_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23835_ _23835_/A VGND VGND VPWR VPWR _32461_/D sky130_fd_sc_hd__clkbuf_1
X_26623_ _25097_/X _33712_/Q _26633_/S VGND VGND VPWR VPWR _26624_/A sky130_fd_sc_hd__mux2_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_404 _36211_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_415 _36212_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_426 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26554_ _24995_/X _33679_/Q _26570_/S VGND VGND VPWR VPWR _26555_/A sky130_fd_sc_hd__mux2_1
X_29342_ _29342_/A VGND VGND VPWR VPWR _34937_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_437 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23766_ _22972_/X _32428_/Q _23784_/S VGND VGND VPWR VPWR _23767_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_448 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20978_ _20687_/X _20976_/X _20977_/X _20697_/X VGND VGND VPWR VPWR _20978_/X sky130_fd_sc_hd__a22o_1
XANTENNA_459 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22717_ _35336_/Q _35272_/Q _35208_/Q _32328_/Q _20688_/X _20690_/X VGND VGND VPWR
+ VPWR _22717_/X sky130_fd_sc_hd__mux4_1
X_25505_ _33185_/Q _24304_/X _25505_/S VGND VGND VPWR VPWR _25506_/A sky130_fd_sc_hd__mux2_1
X_29273_ _29273_/A VGND VGND VPWR VPWR _34904_/D sky130_fd_sc_hd__clkbuf_1
X_26485_ _25094_/X _33647_/Q _26497_/S VGND VGND VPWR VPWR _26486_/A sky130_fd_sc_hd__mux2_1
X_23697_ _23697_/A VGND VGND VPWR VPWR _32397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28224_ _26999_/X _34439_/Q _28228_/S VGND VGND VPWR VPWR _28225_/A sky130_fd_sc_hd__mux2_1
X_25436_ _25153_/X _33154_/Q _25450_/S VGND VGND VPWR VPWR _25437_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_1160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22648_ _22644_/X _22647_/X _22442_/X _22443_/X VGND VGND VPWR VPWR _22663_/B sky130_fd_sc_hd__o211a_2
XFILLER_201_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_194_CLK clkbuf_6_49__f_CLK/X VGND VGND VPWR VPWR _36169_/CLK sky130_fd_sc_hd__clkbuf_16
X_28155_ _26897_/X _34406_/Q _28165_/S VGND VGND VPWR VPWR _28156_/A sky130_fd_sc_hd__mux2_1
X_25367_ _25367_/A VGND VGND VPWR VPWR _33121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22579_ _32772_/Q _32708_/Q _32644_/Q _36100_/Q _22578_/X _22362_/X VGND VGND VPWR
+ VPWR _22579_/X sky130_fd_sc_hd__mux4_1
XFILLER_167_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27106_ _27154_/S VGND VGND VPWR VPWR _27125_/S sky130_fd_sc_hd__buf_4
XFILLER_127_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24318_ _32677_/Q _24317_/X _24336_/S VGND VGND VPWR VPWR _24319_/A sky130_fd_sc_hd__mux2_1
X_28086_ _28086_/A VGND VGND VPWR VPWR _34373_/D sky130_fd_sc_hd__clkbuf_1
X_25298_ _25150_/X _33089_/Q _25314_/S VGND VGND VPWR VPWR _25299_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27037_ _26844_/X _33877_/Q _27041_/S VGND VGND VPWR VPWR _27038_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_952 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24249_ input12/X VGND VGND VPWR VPWR _24249_/X sky130_fd_sc_hd__buf_4
XFILLER_135_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18810_ _35738_/Q _35098_/Q _34458_/Q _33818_/Q _18734_/X _18735_/X VGND VGND VPWR
+ VPWR _18810_/X sky130_fd_sc_hd__mux4_1
XTAP_6030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19790_ _20143_/A VGND VGND VPWR VPWR _19790_/X sky130_fd_sc_hd__clkbuf_4
X_28988_ _34801_/Q _24354_/X _28996_/S VGND VGND VPWR VPWR _28989_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput95 _31964_/Q VGND VGND VPWR VPWR D1[14] sky130_fd_sc_hd__buf_2
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18741_ _20153_/A VGND VGND VPWR VPWR _18741_/X sky130_fd_sc_hd__buf_2
XTAP_6085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27939_ _27966_/S VGND VGND VPWR VPWR _27958_/S sky130_fd_sc_hd__clkbuf_8
XTAP_5340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18672_ _18666_/X _18671_/X _18371_/X VGND VGND VPWR VPWR _18680_/C sky130_fd_sc_hd__o21ba_1
XFILLER_7_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30950_ _30950_/A VGND VGND VPWR VPWR _35699_/D sky130_fd_sc_hd__clkbuf_1
XTAP_5395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17623_ _17555_/X _17621_/X _17622_/X _17558_/X VGND VGND VPWR VPWR _17623_/X sky130_fd_sc_hd__a22o_1
X_29609_ _35064_/Q _29182_/X _29623_/S VGND VGND VPWR VPWR _29610_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30881_ _30881_/A VGND VGND VPWR VPWR _35666_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32620_ _36076_/CLK _32620_/D VGND VGND VPWR VPWR _32620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _17548_/X _17551_/X _17552_/X _17553_/X VGND VGND VPWR VPWR _17554_/X sky130_fd_sc_hd__a22o_1
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_960 _29922_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_971 _31678_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16505_ _32474_/Q _32346_/Q _32026_/Q _35994_/Q _16217_/X _16358_/X VGND VGND VPWR
+ VPWR _16505_/X sky130_fd_sc_hd__mux4_1
X_32551_ _35943_/CLK _32551_/D VGND VGND VPWR VPWR _32551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_982 _17906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17485_ _17408_/X _17483_/X _17484_/X _17414_/X VGND VGND VPWR VPWR _17485_/X sky130_fd_sc_hd__a22o_1
XANTENNA_993 _17860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31502_ _23280_/X _35961_/Q _31514_/S VGND VGND VPWR VPWR _31503_/A sky130_fd_sc_hd__mux2_1
X_19224_ _32486_/Q _32358_/Q _32038_/Q _36006_/Q _19223_/X _19011_/X VGND VGND VPWR
+ VPWR _19224_/X sky130_fd_sc_hd__mux4_1
X_35270_ _35334_/CLK _35270_/D VGND VGND VPWR VPWR _35270_/Q sky130_fd_sc_hd__dfxtp_1
X_16436_ _35736_/Q _35096_/Q _34456_/Q _33816_/Q _16434_/X _16435_/X VGND VGND VPWR
+ VPWR _16436_/X sky130_fd_sc_hd__mux4_1
X_32482_ _36004_/CLK _32482_/D VGND VGND VPWR VPWR _32482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34221_ _35575_/CLK _34221_/D VGND VGND VPWR VPWR _34221_/Q sky130_fd_sc_hd__dfxtp_1
X_31433_ _23117_/X _35928_/Q _31451_/S VGND VGND VPWR VPWR _31434_/A sky130_fd_sc_hd__mux2_1
X_19155_ _32740_/Q _32676_/Q _32612_/Q _36068_/Q _18866_/X _19003_/X VGND VGND VPWR
+ VPWR _19155_/X sky130_fd_sc_hd__mux4_1
X_16367_ _35542_/Q _35478_/Q _35414_/Q _35350_/Q _16191_/X _16192_/X VGND VGND VPWR
+ VPWR _16367_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_185_CLK clkbuf_leaf_66_CLK/A VGND VGND VPWR VPWR _35002_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_199_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18106_ _33032_/Q _32968_/Q _32904_/Q _32840_/Q _15980_/X _15983_/X VGND VGND VPWR
+ VPWR _18106_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34152_ _34279_/CLK _34152_/D VGND VGND VPWR VPWR _34152_/Q sky130_fd_sc_hd__dfxtp_1
X_16298_ _16292_/X _16297_/X _16071_/X VGND VGND VPWR VPWR _16308_/C sky130_fd_sc_hd__o21ba_1
X_19086_ _35810_/Q _32186_/Q _35682_/Q _35618_/Q _18907_/X _18908_/X VGND VGND VPWR
+ VPWR _19086_/X sky130_fd_sc_hd__mux4_1
X_31364_ _31364_/A VGND VGND VPWR VPWR _35895_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33103_ _36112_/CLK _33103_/D VGND VGND VPWR VPWR _33103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18037_ _17901_/X _18035_/X _18036_/X _17906_/X VGND VGND VPWR VPWR _18037_/X sky130_fd_sc_hd__a22o_1
XFILLER_219_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30315_ _35399_/Q _29228_/X _30319_/S VGND VGND VPWR VPWR _30316_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_33__f_CLK clkbuf_5_16_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_33__f_CLK/X sky130_fd_sc_hd__clkbuf_16
X_34083_ _34146_/CLK _34083_/D VGND VGND VPWR VPWR _34083_/Q sky130_fd_sc_hd__dfxtp_1
X_31295_ _35863_/Q input64/X _31295_/S VGND VGND VPWR VPWR _31296_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33034_ _35979_/CLK _33034_/D VGND VGND VPWR VPWR _33034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1001 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30246_ _35366_/Q _29126_/X _30256_/S VGND VGND VPWR VPWR _30247_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30177_ _30177_/A VGND VGND VPWR VPWR _35333_/D sky130_fd_sc_hd__clkbuf_1
X_19988_ _34044_/Q _33980_/Q _33916_/Q _32252_/Q _19673_/X _19674_/X VGND VGND VPWR
+ VPWR _19988_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18939_ _18657_/X _18935_/X _18938_/X _18661_/X VGND VGND VPWR VPWR _18939_/X sky130_fd_sc_hd__a22o_1
X_34985_ _34987_/CLK _34985_/D VGND VGND VPWR VPWR _34985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1370 _24407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1381 _28776_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33936_ _34004_/CLK _33936_/D VGND VGND VPWR VPWR _33936_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1392 _17154_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21950_ _22458_/A VGND VGND VPWR VPWR _21950_/X sky130_fd_sc_hd__buf_4
XFILLER_223_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20901_ _21607_/A VGND VGND VPWR VPWR _20901_/X sky130_fd_sc_hd__buf_4
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33867_ _35787_/CLK _33867_/D VGND VGND VPWR VPWR _33867_/Q sky130_fd_sc_hd__dfxtp_1
X_21881_ _35824_/Q _32201_/Q _35696_/Q _35632_/Q _21560_/X _21561_/X VGND VGND VPWR
+ VPWR _21881_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35606_ _35799_/CLK _35606_/D VGND VGND VPWR VPWR _35606_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23620_ _23620_/A VGND VGND VPWR VPWR _32360_/D sky130_fd_sc_hd__clkbuf_1
X_20832_ _35282_/Q _35218_/Q _35154_/Q _32274_/Q _20679_/X _20681_/X VGND VGND VPWR
+ VPWR _20832_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32818_ _35765_/CLK _32818_/D VGND VGND VPWR VPWR _32818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33798_ _34308_/CLK _33798_/D VGND VGND VPWR VPWR _33798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23551_ _23062_/X _32329_/Q _23551_/S VGND VGND VPWR VPWR _23552_/A sky130_fd_sc_hd__mux2_1
XFILLER_223_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35537_ _35921_/CLK _35537_/D VGND VGND VPWR VPWR _35537_/Q sky130_fd_sc_hd__dfxtp_1
X_20763_ _34768_/Q _34704_/Q _34640_/Q _34576_/Q _20675_/X _20676_/X VGND VGND VPWR
+ VPWR _20763_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32749_ _36077_/CLK _32749_/D VGND VGND VPWR VPWR _32749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22502_ _22502_/A VGND VGND VPWR VPWR _22502_/X sky130_fd_sc_hd__buf_8
XFILLER_168_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26270_ _26270_/A VGND VGND VPWR VPWR _33545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35468_ _35532_/CLK _35468_/D VGND VGND VPWR VPWR _35468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_958 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23482_ _22960_/X _32296_/Q _23488_/S VGND VGND VPWR VPWR _23483_/A sky130_fd_sc_hd__mux2_1
X_20694_ _21757_/A VGND VGND VPWR VPWR _20694_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25221_ _25221_/A VGND VGND VPWR VPWR _33052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_241_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22433_ _22155_/X _22431_/X _22432_/X _22158_/X VGND VGND VPWR VPWR _22433_/X sky130_fd_sc_hd__a22o_1
X_34419_ _34805_/CLK _34419_/D VGND VGND VPWR VPWR _34419_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_176_CLK clkbuf_6_27__f_CLK/X VGND VGND VPWR VPWR _34060_/CLK sky130_fd_sc_hd__clkbuf_16
X_35399_ _35590_/CLK _35399_/D VGND VGND VPWR VPWR _35399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25152_ _25152_/A VGND VGND VPWR VPWR _33025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22364_ _22582_/A VGND VGND VPWR VPWR _22364_/X sky130_fd_sc_hd__buf_4
XFILLER_248_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24103_ _24103_/A VGND VGND VPWR VPWR _32587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21315_ _21310_/X _21312_/X _21313_/X _21314_/X VGND VGND VPWR VPWR _21315_/X sky130_fd_sc_hd__a22o_1
XFILLER_184_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29960_ _29960_/A VGND VGND VPWR VPWR _35230_/D sky130_fd_sc_hd__clkbuf_1
X_25083_ _25083_/A VGND VGND VPWR VPWR _33003_/D sky130_fd_sc_hd__clkbuf_1
X_22295_ _22429_/A VGND VGND VPWR VPWR _22295_/X sky130_fd_sc_hd__buf_4
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28911_ _27017_/X _34765_/Q _28911_/S VGND VGND VPWR VPWR _28912_/A sky130_fd_sc_hd__mux2_1
X_24034_ _24034_/A VGND VGND VPWR VPWR _32554_/D sky130_fd_sc_hd__clkbuf_1
X_21246_ _22460_/A VGND VGND VPWR VPWR _21246_/X sky130_fd_sc_hd__clkbuf_4
X_29891_ _35198_/Q _29200_/X _29893_/S VGND VGND VPWR VPWR _29892_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28842_ _28911_/S VGND VGND VPWR VPWR _28861_/S sky130_fd_sc_hd__buf_4
X_21177_ _20888_/X _21175_/X _21176_/X _20891_/X VGND VGND VPWR VPWR _21177_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20128_ _19848_/X _20126_/X _20127_/X _19853_/X VGND VGND VPWR VPWR _20128_/X sky130_fd_sc_hd__a22o_1
X_28773_ _28773_/A VGND VGND VPWR VPWR _34699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_1142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25985_ _25153_/X _33410_/Q _25999_/S VGND VGND VPWR VPWR _25986_/A sky130_fd_sc_hd__mux2_1
XFILLER_219_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27724_ _27724_/A VGND VGND VPWR VPWR _34201_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_100_CLK clkbuf_leaf_99_CLK/A VGND VGND VPWR VPWR _36204_/CLK sky130_fd_sc_hd__clkbuf_16
X_20059_ _19855_/X _20057_/X _20058_/X _19858_/X VGND VGND VPWR VPWR _20059_/X sky130_fd_sc_hd__a22o_1
XFILLER_150_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24936_ _24936_/A VGND VGND VPWR VPWR _32948_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27655_ _34169_/Q _24379_/X _27667_/S VGND VGND VPWR VPWR _27656_/A sky130_fd_sc_hd__mux2_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24867_ _24867_/A VGND VGND VPWR VPWR _32915_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_212 _32135_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_223 _32136_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26606_ _25072_/X _33704_/Q _26612_/S VGND VGND VPWR VPWR _26607_/A sky130_fd_sc_hd__mux2_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23818_ _23050_/X _32453_/Q _23826_/S VGND VGND VPWR VPWR _23819_/A sky130_fd_sc_hd__mux2_1
XANTENNA_234 _32136_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_245 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27586_ _34136_/Q _24276_/X _27604_/S VGND VGND VPWR VPWR _27587_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24798_ _22994_/X _32883_/Q _24802_/S VGND VGND VPWR VPWR _24799_/A sky130_fd_sc_hd__mux2_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 _32137_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_267 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29325_ _29325_/A VGND VGND VPWR VPWR _34929_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26537_ _25171_/X _33672_/Q _26539_/S VGND VGND VPWR VPWR _26538_/A sky130_fd_sc_hd__mux2_1
XANTENNA_278 _32138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23749_ _22948_/X _32420_/Q _23763_/S VGND VGND VPWR VPWR _23750_/A sky130_fd_sc_hd__mux2_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_289 _32139_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29256_ _29256_/A VGND VGND VPWR VPWR _34896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_1247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17270_ _17202_/X _17268_/X _17269_/X _17205_/X VGND VGND VPWR VPWR _17270_/X sky130_fd_sc_hd__a22o_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26468_ _25069_/X _33639_/Q _26476_/S VGND VGND VPWR VPWR _26469_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28207_ _26974_/X _34431_/Q _28207_/S VGND VGND VPWR VPWR _28208_/A sky130_fd_sc_hd__mux2_1
X_16221_ _16216_/X _16220_/X _16040_/X _16042_/X VGND VGND VPWR VPWR _16238_/B sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_167_CLK clkbuf_6_28__f_CLK/X VGND VGND VPWR VPWR _36109_/CLK sky130_fd_sc_hd__clkbuf_16
X_25419_ _25128_/X _33146_/Q _25429_/S VGND VGND VPWR VPWR _25420_/A sky130_fd_sc_hd__mux2_1
X_26399_ _26399_/A VGND VGND VPWR VPWR _33606_/D sky130_fd_sc_hd__clkbuf_1
X_29187_ _29187_/A VGND VGND VPWR VPWR _34873_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16152_ _32464_/Q _32336_/Q _32016_/Q _35984_/Q _16028_/X _17863_/A VGND VGND VPWR
+ VPWR _16152_/X sky130_fd_sc_hd__mux4_1
XFILLER_220_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28138_ _26872_/X _34398_/Q _28144_/S VGND VGND VPWR VPWR _28139_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16083_ _17767_/A VGND VGND VPWR VPWR _17152_/A sky130_fd_sc_hd__buf_12
XFILLER_154_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28069_ _28069_/A VGND VGND VPWR VPWR _34365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19911_ _19802_/X _19909_/X _19910_/X _19805_/X VGND VGND VPWR VPWR _19911_/X sky130_fd_sc_hd__a22o_1
X_30100_ _35297_/Q _29110_/X _30100_/S VGND VGND VPWR VPWR _30101_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31080_ _35761_/Q _29160_/X _31088_/S VGND VGND VPWR VPWR _31081_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30031_ _35264_/Q _29206_/X _30049_/S VGND VGND VPWR VPWR _30032_/A sky130_fd_sc_hd__mux2_1
X_19842_ _34551_/Q _32439_/Q _34423_/Q _34359_/Q _19525_/X _19526_/X VGND VGND VPWR
+ VPWR _19842_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19773_ _33782_/Q _33718_/Q _33654_/Q _33590_/Q _19496_/X _19497_/X VGND VGND VPWR
+ VPWR _19773_/X sky130_fd_sc_hd__mux4_1
X_16985_ _32744_/Q _32680_/Q _32616_/Q _36072_/Q _16919_/X _16703_/X VGND VGND VPWR
+ VPWR _16985_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18724_ _32728_/Q _32664_/Q _32600_/Q _36056_/Q _18513_/X _18650_/X VGND VGND VPWR
+ VPWR _18724_/X sky130_fd_sc_hd__mux4_1
XTAP_5170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34770_ _35669_/CLK _34770_/D VGND VGND VPWR VPWR _34770_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31982_ _35293_/CLK _31982_/D VGND VGND VPWR VPWR _31982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33721_ _34297_/CLK _33721_/D VGND VGND VPWR VPWR _33721_/Q sky130_fd_sc_hd__dfxtp_1
X_18655_ _20206_/A VGND VGND VPWR VPWR _18655_/X sky130_fd_sc_hd__clkbuf_4
X_30933_ _30933_/A VGND VGND VPWR VPWR _35691_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17606_ _33209_/Q _32569_/Q _35961_/Q _35897_/Q _17427_/X _17428_/X VGND VGND VPWR
+ VPWR _17606_/X sky130_fd_sc_hd__mux4_1
X_33652_ _34289_/CLK _33652_/D VGND VGND VPWR VPWR _33652_/Q sky130_fd_sc_hd__dfxtp_1
X_30864_ _23339_/X _35659_/Q _30868_/S VGND VGND VPWR VPWR _30865_/A sky130_fd_sc_hd__mux2_1
X_18586_ _18326_/X _18582_/X _18585_/X _18337_/X VGND VGND VPWR VPWR _18586_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32603_ _36059_/CLK _32603_/D VGND VGND VPWR VPWR _32603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17537_ _17352_/X _17535_/X _17536_/X _17355_/X VGND VGND VPWR VPWR _17537_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33583_ _33775_/CLK _33583_/D VGND VGND VPWR VPWR _33583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30795_ _23231_/X _35626_/Q _30797_/S VGND VGND VPWR VPWR _30796_/A sky130_fd_sc_hd__mux2_1
XANTENNA_790 _22664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35322_ _35579_/CLK _35322_/D VGND VGND VPWR VPWR _35322_/Q sky130_fd_sc_hd__dfxtp_1
X_32534_ _36118_/CLK _32534_/D VGND VGND VPWR VPWR _32534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_958 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17468_ _35061_/Q _34997_/Q _34933_/Q _34869_/Q _17156_/X _17157_/X VGND VGND VPWR
+ VPWR _17468_/X sky130_fd_sc_hd__mux4_1
X_19207_ _35045_/Q _34981_/Q _34917_/Q _34853_/Q _19103_/X _19104_/X VGND VGND VPWR
+ VPWR _19207_/X sky130_fd_sc_hd__mux4_1
X_16419_ _33496_/Q _33432_/Q _33368_/Q _33304_/Q _16417_/X _16418_/X VGND VGND VPWR
+ VPWR _16419_/X sky130_fd_sc_hd__mux4_1
X_35253_ _35315_/CLK _35253_/D VGND VGND VPWR VPWR _35253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_158_CLK clkbuf_6_31__f_CLK/X VGND VGND VPWR VPWR _35851_/CLK sky130_fd_sc_hd__clkbuf_16
X_32465_ _35985_/CLK _32465_/D VGND VGND VPWR VPWR _32465_/Q sky130_fd_sc_hd__dfxtp_1
X_17399_ _17399_/A _17399_/B _17399_/C _17399_/D VGND VGND VPWR VPWR _17400_/A sky130_fd_sc_hd__or4_4
X_34204_ _34777_/CLK _34204_/D VGND VGND VPWR VPWR _34204_/Q sky130_fd_sc_hd__dfxtp_1
X_31416_ _23093_/X _35920_/Q _31430_/S VGND VGND VPWR VPWR _31417_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19138_ _19101_/X _19136_/X _19137_/X _19106_/X VGND VGND VPWR VPWR _19138_/X sky130_fd_sc_hd__a22o_1
XFILLER_160_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35184_ _35757_/CLK _35184_/D VGND VGND VPWR VPWR _35184_/Q sky130_fd_sc_hd__dfxtp_1
X_32396_ _36109_/CLK _32396_/D VGND VGND VPWR VPWR _32396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34135_ _35669_/CLK _34135_/D VGND VGND VPWR VPWR _34135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_218_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31347_ _31347_/A VGND VGND VPWR VPWR _35887_/D sky130_fd_sc_hd__clkbuf_1
X_19069_ _18789_/X _19067_/X _19068_/X _18794_/X VGND VGND VPWR VPWR _19069_/X sky130_fd_sc_hd__a22o_1
XFILLER_172_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21100_ _21096_/X _21097_/X _21098_/X _21099_/X VGND VGND VPWR VPWR _21100_/X sky130_fd_sc_hd__a22o_1
XFILLER_191_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34066_ _34256_/CLK _34066_/D VGND VGND VPWR VPWR _34066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22080_ _21802_/X _22078_/X _22079_/X _21805_/X VGND VGND VPWR VPWR _22080_/X sky130_fd_sc_hd__a22o_1
XFILLER_47_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31278_ _31278_/A VGND VGND VPWR VPWR _35854_/D sky130_fd_sc_hd__clkbuf_1
X_33017_ _36090_/CLK _33017_/D VGND VGND VPWR VPWR _33017_/Q sky130_fd_sc_hd__dfxtp_1
X_21031_ _22443_/A VGND VGND VPWR VPWR _21031_/X sky130_fd_sc_hd__buf_4
X_30229_ _35358_/Q _29101_/X _30235_/S VGND VGND VPWR VPWR _30230_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_330_CLK clkbuf_6_45__f_CLK/X VGND VGND VPWR VPWR _36022_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22982_ input27/X VGND VGND VPWR VPWR _22982_/X sky130_fd_sc_hd__clkbuf_4
X_34968_ _35292_/CLK _34968_/D VGND VGND VPWR VPWR _34968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25770_ _25035_/X _33308_/Q _25780_/S VGND VGND VPWR VPWR _25771_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24721_ _22875_/X _32846_/Q _24739_/S VGND VGND VPWR VPWR _24722_/A sky130_fd_sc_hd__mux2_1
X_21933_ _21795_/X _21931_/X _21932_/X _21800_/X VGND VGND VPWR VPWR _21933_/X sky130_fd_sc_hd__a22o_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33919_ _34046_/CLK _33919_/D VGND VGND VPWR VPWR _33919_/Q sky130_fd_sc_hd__dfxtp_1
X_34899_ _34967_/CLK _34899_/D VGND VGND VPWR VPWR _34899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27440_ _26841_/X _34068_/Q _27446_/S VGND VGND VPWR VPWR _27441_/A sky130_fd_sc_hd__mux2_1
X_24652_ _24652_/A VGND VGND VPWR VPWR _32814_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21864_ _21864_/A VGND VGND VPWR VPWR _36207_/D sky130_fd_sc_hd__buf_6
XFILLER_70_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23603_ _23603_/A VGND VGND VPWR VPWR _32352_/D sky130_fd_sc_hd__clkbuf_1
X_20815_ _33234_/Q _36114_/Q _33106_/Q _33042_/Q _20620_/X _20621_/X VGND VGND VPWR
+ VPWR _20815_/X sky130_fd_sc_hd__mux4_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24583_ _24715_/S VGND VGND VPWR VPWR _24602_/S sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_397_CLK clkbuf_6_34__f_CLK/X VGND VGND VPWR VPWR _35949_/CLK sky130_fd_sc_hd__clkbuf_16
X_27371_ _27371_/A VGND VGND VPWR VPWR _34035_/D sky130_fd_sc_hd__clkbuf_1
X_21795_ _22501_/A VGND VGND VPWR VPWR _21795_/X sky130_fd_sc_hd__buf_2
XFILLER_169_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29110_ input11/X VGND VGND VPWR VPWR _29110_/X sky130_fd_sc_hd__buf_2
XFILLER_93_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23534_ _23534_/A VGND VGND VPWR VPWR _32320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26322_ _26412_/S VGND VGND VPWR VPWR _26341_/S sky130_fd_sc_hd__buf_4
X_20746_ _22465_/A VGND VGND VPWR VPWR _20746_/X sky130_fd_sc_hd__buf_4
X_29041_ _29041_/A VGND VGND VPWR VPWR _34826_/D sky130_fd_sc_hd__clkbuf_1
X_26253_ _25150_/X _33537_/Q _26269_/S VGND VGND VPWR VPWR _26254_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_149_CLK clkbuf_6_29__f_CLK/X VGND VGND VPWR VPWR _35788_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_183_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23465_ _22935_/X _32288_/Q _23467_/S VGND VGND VPWR VPWR _23466_/A sky130_fd_sc_hd__mux2_1
X_20677_ _34766_/Q _34702_/Q _34638_/Q _34574_/Q _20675_/X _20676_/X VGND VGND VPWR
+ VPWR _20677_/X sky130_fd_sc_hd__mux4_1
X_25204_ _25204_/A VGND VGND VPWR VPWR _33044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22416_ _22412_/X _22415_/X _22100_/X VGND VGND VPWR VPWR _22424_/C sky130_fd_sc_hd__o21ba_1
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26184_ _26184_/A VGND VGND VPWR VPWR _33504_/D sky130_fd_sc_hd__clkbuf_1
X_23396_ _23396_/A VGND VGND VPWR VPWR _32256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25135_ _25134_/X _33020_/Q _25144_/S VGND VGND VPWR VPWR _25136_/A sky130_fd_sc_hd__mux2_1
X_22347_ _22102_/X _22345_/X _22346_/X _22105_/X VGND VGND VPWR VPWR _22347_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29943_ _29943_/A VGND VGND VPWR VPWR _35222_/D sky130_fd_sc_hd__clkbuf_1
X_25066_ input17/X VGND VGND VPWR VPWR _25066_/X sky130_fd_sc_hd__buf_2
XFILLER_163_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22278_ _34555_/Q _32443_/Q _34427_/Q _34363_/Q _22178_/X _22179_/X VGND VGND VPWR
+ VPWR _22278_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24017_ _22941_/X _32546_/Q _24035_/S VGND VGND VPWR VPWR _24018_/A sky130_fd_sc_hd__mux2_1
X_21229_ _34014_/Q _33950_/Q _33886_/Q _32158_/Q _20914_/X _20915_/X VGND VGND VPWR
+ VPWR _21229_/X sky130_fd_sc_hd__mux4_1
X_29874_ _29922_/S VGND VGND VPWR VPWR _29893_/S sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_321_CLK clkbuf_6_38__f_CLK/X VGND VGND VPWR VPWR _35252_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_104_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28825_ _28825_/A VGND VGND VPWR VPWR _34723_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28756_ _26987_/X _34691_/Q _28768_/S VGND VGND VPWR VPWR _28757_/A sky130_fd_sc_hd__mux2_1
X_16770_ _17829_/A VGND VGND VPWR VPWR _16770_/X sky130_fd_sc_hd__buf_4
XFILLER_219_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25968_ _25128_/X _33402_/Q _25978_/S VGND VGND VPWR VPWR _25969_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27707_ _27707_/A VGND VGND VPWR VPWR _34193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24919_ _22972_/X _32940_/Q _24937_/S VGND VGND VPWR VPWR _24920_/A sky130_fd_sc_hd__mux2_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28687_ _26884_/X _34658_/Q _28705_/S VGND VGND VPWR VPWR _28688_/A sky130_fd_sc_hd__mux2_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25899_ _25026_/X _33369_/Q _25915_/S VGND VGND VPWR VPWR _25900_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _34256_/Q _34192_/Q _34128_/Q _34064_/Q _18305_/X _18307_/X VGND VGND VPWR
+ VPWR _18440_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27638_ _34161_/Q _24354_/X _27646_/S VGND VGND VPWR VPWR _27639_/A sky130_fd_sc_hd__mux2_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _20153_/A VGND VGND VPWR VPWR _18371_/X sky130_fd_sc_hd__buf_2
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27569_ _34128_/Q _24252_/X _27583_/S VGND VGND VPWR VPWR _27570_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_388_CLK clkbuf_6_35__f_CLK/X VGND VGND VPWR VPWR _34866_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29308_ _29308_/A VGND VGND VPWR VPWR _34921_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _34801_/Q _34737_/Q _34673_/Q _34609_/Q _17288_/X _17289_/X VGND VGND VPWR
+ VPWR _17322_/X sky130_fd_sc_hd__mux4_1
X_30580_ _23316_/X _35524_/Q _30590_/S VGND VGND VPWR VPWR _30581_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29239_ _29239_/A VGND VGND VPWR VPWR _34890_/D sky130_fd_sc_hd__clkbuf_1
X_17253_ _33199_/Q _32559_/Q _35951_/Q _35887_/Q _17074_/X _17075_/X VGND VGND VPWR
+ VPWR _17253_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16204_ _16204_/A _16204_/B _16204_/C _16204_/D VGND VGND VPWR VPWR _16205_/A sky130_fd_sc_hd__or4_4
XFILLER_161_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32250_ _36154_/CLK _32250_/D VGND VGND VPWR VPWR _32250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17184_ _16999_/X _17182_/X _17183_/X _17002_/X VGND VGND VPWR VPWR _17184_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31201_ _31201_/A VGND VGND VPWR VPWR _35818_/D sky130_fd_sc_hd__clkbuf_1
X_16135_ _16135_/A VGND VGND VPWR VPWR _31951_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32181_ _35809_/CLK _32181_/D VGND VGND VPWR VPWR _32181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31132_ _35786_/Q _29237_/X _31138_/S VGND VGND VPWR VPWR _31133_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16066_ _33166_/Q _32526_/Q _35918_/Q _35854_/Q _16063_/X _16065_/X VGND VGND VPWR
+ VPWR _16066_/X sky130_fd_sc_hd__mux4_1
XFILLER_142_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31063_ _35753_/Q _29135_/X _31067_/S VGND VGND VPWR VPWR _31064_/A sky130_fd_sc_hd__mux2_1
X_35940_ _35940_/CLK _35940_/D VGND VGND VPWR VPWR _35940_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_312_CLK clkbuf_6_37__f_CLK/X VGND VGND VPWR VPWR _35318_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_151_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30014_ _35256_/Q _29182_/X _30028_/S VGND VGND VPWR VPWR _30015_/A sky130_fd_sc_hd__mux2_1
X_19825_ _32759_/Q _32695_/Q _32631_/Q _36087_/Q _19572_/X _19709_/X VGND VGND VPWR
+ VPWR _19825_/X sky130_fd_sc_hd__mux4_1
X_35871_ _35937_/CLK _35871_/D VGND VGND VPWR VPWR _35871_/Q sky130_fd_sc_hd__dfxtp_1
X_34822_ _34822_/CLK _34822_/D VGND VGND VPWR VPWR _34822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19756_ _19752_/X _19755_/X _19436_/X _19437_/X VGND VGND VPWR VPWR _19771_/B sky130_fd_sc_hd__o211a_1
XFILLER_238_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16968_ _16964_/X _16967_/X _16794_/X VGND VGND VPWR VPWR _16976_/C sky130_fd_sc_hd__o21ba_1
XFILLER_225_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18707_ _18374_/X _18705_/X _18706_/X _18384_/X VGND VGND VPWR VPWR _18707_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34753_ _34817_/CLK _34753_/D VGND VGND VPWR VPWR _34753_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_16_0_CLK clkbuf_2_2_0_CLK/X VGND VGND VPWR VPWR clkbuf_5_16_0_CLK/X sky130_fd_sc_hd__clkbuf_8
XFILLER_237_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31965_ _35166_/CLK _31965_/D VGND VGND VPWR VPWR _31965_/Q sky130_fd_sc_hd__dfxtp_1
X_19687_ _19647_/X _19685_/X _19686_/X _19650_/X VGND VGND VPWR VPWR _19687_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16899_ _35557_/Q _35493_/Q _35429_/Q _35365_/Q _16897_/X _16898_/X VGND VGND VPWR
+ VPWR _16899_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33704_ _34870_/CLK _33704_/D VGND VGND VPWR VPWR _33704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18638_ _18387_/X _18636_/X _18637_/X _18397_/X VGND VGND VPWR VPWR _18638_/X sky130_fd_sc_hd__a22o_1
X_30916_ _35683_/Q _29117_/X _30932_/S VGND VGND VPWR VPWR _30917_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34684_ _35707_/CLK _34684_/D VGND VGND VPWR VPWR _34684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31896_ _23264_/X _36148_/Q _31898_/S VGND VGND VPWR VPWR _31897_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33635_ _33635_/CLK _33635_/D VGND VGND VPWR VPWR _33635_/Q sky130_fd_sc_hd__dfxtp_1
X_30847_ _30847_/A VGND VGND VPWR VPWR _35650_/D sky130_fd_sc_hd__clkbuf_1
X_18569_ _18565_/X _18568_/X _18400_/X VGND VGND VPWR VPWR _18570_/D sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_379_CLK clkbuf_6_40__f_CLK/X VGND VGND VPWR VPWR _35951_/CLK sky130_fd_sc_hd__clkbuf_16
X_20600_ _33486_/Q _33422_/Q _33358_/Q _33294_/Q _20598_/X _20599_/X VGND VGND VPWR
+ VPWR _20600_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33566_ _34010_/CLK _33566_/D VGND VGND VPWR VPWR _33566_/Q sky130_fd_sc_hd__dfxtp_1
X_21580_ _21442_/X _21578_/X _21579_/X _21447_/X VGND VGND VPWR VPWR _21580_/X sky130_fd_sc_hd__a22o_1
XFILLER_244_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30778_ _30868_/S VGND VGND VPWR VPWR _30797_/S sky130_fd_sc_hd__buf_4
XFILLER_36_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35305_ _35307_/CLK _35305_/D VGND VGND VPWR VPWR _35305_/Q sky130_fd_sc_hd__dfxtp_1
X_20531_ _18277_/X _20529_/X _20530_/X _18287_/X VGND VGND VPWR VPWR _20531_/X sky130_fd_sc_hd__a22o_1
X_32517_ _36037_/CLK _32517_/D VGND VGND VPWR VPWR _32517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33497_ _34267_/CLK _33497_/D VGND VGND VPWR VPWR _33497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23250_ input28/X VGND VGND VPWR VPWR _23250_/X sky130_fd_sc_hd__clkbuf_4
X_35236_ _35300_/CLK _35236_/D VGND VGND VPWR VPWR _35236_/Q sky130_fd_sc_hd__dfxtp_1
X_32448_ _32967_/CLK _32448_/D VGND VGND VPWR VPWR _32448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20462_ _32778_/Q _32714_/Q _32650_/Q _36106_/Q _20278_/X _19173_/A VGND VGND VPWR
+ VPWR _20462_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22201_ _35769_/Q _35129_/Q _34489_/Q _33849_/Q _22093_/X _22094_/X VGND VGND VPWR
+ VPWR _22201_/X sky130_fd_sc_hd__mux4_1
X_23181_ _23181_/A VGND VGND VPWR VPWR _32173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35167_ _35294_/CLK _35167_/D VGND VGND VPWR VPWR _35167_/Q sky130_fd_sc_hd__dfxtp_1
X_20393_ _20393_/A _20393_/B _20393_/C _20393_/D VGND VGND VPWR VPWR _20394_/A sky130_fd_sc_hd__or4_1
X_32379_ _36028_/CLK _32379_/D VGND VGND VPWR VPWR _32379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34118_ _34312_/CLK _34118_/D VGND VGND VPWR VPWR _34118_/Q sky130_fd_sc_hd__dfxtp_1
X_22132_ _35831_/Q _32209_/Q _35703_/Q _35639_/Q _21913_/X _21914_/X VGND VGND VPWR
+ VPWR _22132_/X sky130_fd_sc_hd__mux4_1
XFILLER_134_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput230 _32098_/Q VGND VGND VPWR VPWR D3[20] sky130_fd_sc_hd__buf_2
X_35098_ _35098_/CLK _35098_/D VGND VGND VPWR VPWR _35098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput241 _32108_/Q VGND VGND VPWR VPWR D3[30] sky130_fd_sc_hd__buf_2
XFILLER_86_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput252 _32118_/Q VGND VGND VPWR VPWR D3[40] sky130_fd_sc_hd__buf_2
XTAP_6618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34049_ _34305_/CLK _34049_/D VGND VGND VPWR VPWR _34049_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput263 _32128_/Q VGND VGND VPWR VPWR D3[50] sky130_fd_sc_hd__buf_2
X_26940_ input32/X VGND VGND VPWR VPWR _26940_/X sky130_fd_sc_hd__clkbuf_4
X_22063_ _22059_/X _22062_/X _21747_/X VGND VGND VPWR VPWR _22071_/C sky130_fd_sc_hd__o21ba_1
XFILLER_82_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_303_CLK clkbuf_6_50__f_CLK/X VGND VGND VPWR VPWR _34811_/CLK sky130_fd_sc_hd__clkbuf_16
Xoutput274 _32138_/Q VGND VGND VPWR VPWR D3[60] sky130_fd_sc_hd__buf_2
XFILLER_58_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21014_ _33752_/Q _33688_/Q _33624_/Q _33560_/Q _20737_/X _20738_/X VGND VGND VPWR
+ VPWR _21014_/X sky130_fd_sc_hd__mux4_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26871_ _26871_/A VGND VGND VPWR VPWR _33821_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28610_ _26971_/X _34622_/Q _28612_/S VGND VGND VPWR VPWR _28611_/A sky130_fd_sc_hd__mux2_1
X_25822_ _25112_/X _33333_/Q _25822_/S VGND VGND VPWR VPWR _25823_/A sky130_fd_sc_hd__mux2_1
X_29590_ _35055_/Q _29154_/X _29602_/S VGND VGND VPWR VPWR _29591_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28541_ _26869_/X _34589_/Q _28549_/S VGND VGND VPWR VPWR _28542_/A sky130_fd_sc_hd__mux2_1
X_25753_ _25010_/X _33300_/Q _25759_/S VGND VGND VPWR VPWR _25754_/A sky130_fd_sc_hd__mux2_1
XFILLER_228_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22965_ _22965_/A VGND VGND VPWR VPWR _32041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24704_ _24704_/A VGND VGND VPWR VPWR _32839_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28472_ _28472_/A VGND VGND VPWR VPWR _34556_/D sky130_fd_sc_hd__clkbuf_1
X_21916_ _35761_/Q _35121_/Q _34481_/Q _33841_/Q _21740_/X _21741_/X VGND VGND VPWR
+ VPWR _21916_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22896_ _22895_/X _32019_/Q _22908_/S VGND VGND VPWR VPWR _22897_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25684_ _25684_/A VGND VGND VPWR VPWR _33268_/D sky130_fd_sc_hd__clkbuf_1
X_27423_ _27423_/A VGND VGND VPWR VPWR _34060_/D sky130_fd_sc_hd__clkbuf_1
X_21847_ _35823_/Q _32200_/Q _35695_/Q _35631_/Q _21560_/X _21561_/X VGND VGND VPWR
+ VPWR _21847_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_1350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24635_ _24635_/A VGND VGND VPWR VPWR _32806_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_231_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24566_ _24566_/A VGND VGND VPWR VPWR _32775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27354_ _27354_/A VGND VGND VPWR VPWR _34027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21778_ _21774_/X _21777_/X _21736_/X _21737_/X VGND VGND VPWR VPWR _21793_/B sky130_fd_sc_hd__o211a_1
XFILLER_19_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26305_ _26305_/A VGND VGND VPWR VPWR _33561_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20729_ _20674_/X _20727_/X _20728_/X _20684_/X VGND VGND VPWR VPWR _20729_/X sky130_fd_sc_hd__a22o_1
XFILLER_156_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23517_ _23517_/A VGND VGND VPWR VPWR _32312_/D sky130_fd_sc_hd__clkbuf_1
X_27285_ _27011_/X _33995_/Q _27289_/S VGND VGND VPWR VPWR _27286_/A sky130_fd_sc_hd__mux2_1
X_24497_ _24497_/A VGND VGND VPWR VPWR _32742_/D sky130_fd_sc_hd__clkbuf_1
X_29024_ _34818_/Q _24407_/X _29038_/S VGND VGND VPWR VPWR _29025_/A sky130_fd_sc_hd__mux2_1
X_26236_ _25125_/X _33529_/Q _26248_/S VGND VGND VPWR VPWR _26237_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23448_ _23559_/S VGND VGND VPWR VPWR _23467_/S sky130_fd_sc_hd__buf_4
XFILLER_184_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23379_ _23379_/A VGND VGND VPWR VPWR _32248_/D sky130_fd_sc_hd__clkbuf_1
X_26167_ _25022_/X _33496_/Q _26185_/S VGND VGND VPWR VPWR _26168_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25118_ _25118_/A VGND VGND VPWR VPWR _33014_/D sky130_fd_sc_hd__clkbuf_1
X_26098_ _26098_/A VGND VGND VPWR VPWR _33463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17940_ _34307_/Q _34243_/Q _34179_/Q _34115_/Q _17795_/X _17796_/X VGND VGND VPWR
+ VPWR _17940_/X sky130_fd_sc_hd__mux4_1
X_29926_ _35214_/Q _29048_/X _29944_/S VGND VGND VPWR VPWR _29927_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25049_ _25049_/A VGND VGND VPWR VPWR _32992_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_1302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1034 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17871_ _33793_/Q _33729_/Q _33665_/Q _33601_/Q _17549_/X _17550_/X VGND VGND VPWR
+ VPWR _17871_/X sky130_fd_sc_hd__mux4_1
X_29857_ _29857_/A VGND VGND VPWR VPWR _35181_/D sky130_fd_sc_hd__clkbuf_1
X_19610_ _33009_/Q _32945_/Q _32881_/Q _32817_/Q _19289_/X _19290_/X VGND VGND VPWR
+ VPWR _19610_/X sky130_fd_sc_hd__mux4_1
X_16822_ _32483_/Q _32355_/Q _32035_/Q _36003_/Q _16570_/X _16711_/X VGND VGND VPWR
+ VPWR _16822_/X sky130_fd_sc_hd__mux4_1
X_28808_ _28808_/A VGND VGND VPWR VPWR _34715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29788_ _29788_/A VGND VGND VPWR VPWR _35149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_948 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19541_ _33263_/Q _36143_/Q _33135_/Q _33071_/Q _19358_/X _19359_/X VGND VGND VPWR
+ VPWR _19541_/X sky130_fd_sc_hd__mux4_1
XFILLER_219_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28739_ _26962_/X _34683_/Q _28747_/S VGND VGND VPWR VPWR _28740_/A sky130_fd_sc_hd__mux2_1
X_16753_ _16641_/X _16751_/X _16752_/X _16644_/X VGND VGND VPWR VPWR _16753_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19472_ _32749_/Q _32685_/Q _32621_/Q _36077_/Q _19219_/X _19356_/X VGND VGND VPWR
+ VPWR _19472_/X sky130_fd_sc_hd__mux4_1
X_31750_ _31750_/A VGND VGND VPWR VPWR _36078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16684_ _16646_/X _16682_/X _16683_/X _16649_/X VGND VGND VPWR VPWR _16684_/X sky130_fd_sc_hd__a22o_1
XFILLER_94_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18423_ _35535_/Q _35471_/Q _35407_/Q _35343_/Q _18358_/X _18360_/X VGND VGND VPWR
+ VPWR _18423_/X sky130_fd_sc_hd__mux4_1
X_30701_ _30701_/A VGND VGND VPWR VPWR _35581_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31681_ _31813_/S VGND VGND VPWR VPWR _31700_/S sky130_fd_sc_hd__buf_4
XFILLER_37_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33420_ _34060_/CLK _33420_/D VGND VGND VPWR VPWR _33420_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18354_ _20158_/A VGND VGND VPWR VPWR _18354_/X sky130_fd_sc_hd__buf_4
X_30632_ _30632_/A VGND VGND VPWR VPWR _35548_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _17301_/X _17304_/X _17128_/X VGND VGND VPWR VPWR _17329_/A sky130_fd_sc_hd__o21ba_1
X_33351_ _33544_/CLK _33351_/D VGND VGND VPWR VPWR _33351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18285_ input79/X input80/X VGND VGND VPWR VPWR _20067_/A sky130_fd_sc_hd__nor2_4
X_30563_ _23289_/X _35516_/Q _30569_/S VGND VGND VPWR VPWR _30564_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32302_ _35054_/CLK _32302_/D VGND VGND VPWR VPWR _32302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17236_ _33519_/Q _33455_/Q _33391_/Q _33327_/Q _17123_/X _17124_/X VGND VGND VPWR
+ VPWR _17236_/X sky130_fd_sc_hd__mux4_1
X_36070_ _36070_/CLK _36070_/D VGND VGND VPWR VPWR _36070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33282_ _36165_/CLK _33282_/D VGND VGND VPWR VPWR _33282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30494_ _23127_/X _35483_/Q _30506_/S VGND VGND VPWR VPWR _30495_/A sky130_fd_sc_hd__mux2_1
X_35021_ _35021_/CLK _35021_/D VGND VGND VPWR VPWR _35021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32233_ _35853_/CLK _32233_/D VGND VGND VPWR VPWR _32233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17167_ _16842_/X _17165_/X _17166_/X _16847_/X VGND VGND VPWR VPWR _17167_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_982 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16118_ _16026_/X _16116_/X _16117_/X _16037_/X VGND VGND VPWR VPWR _16118_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32164_ _35727_/CLK _32164_/D VGND VGND VPWR VPWR _32164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17098_ _33259_/Q _36139_/Q _33131_/Q _33067_/Q _17058_/X _17059_/X VGND VGND VPWR
+ VPWR _17098_/X sky130_fd_sc_hd__mux4_1
XFILLER_100_1470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31115_ _31115_/A VGND VGND VPWR VPWR _35777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16049_ _17994_/A VGND VGND VPWR VPWR _16049_/X sky130_fd_sc_hd__buf_6
XFILLER_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32095_ _35807_/CLK _32095_/D VGND VGND VPWR VPWR _32095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35923_ _35925_/CLK _35923_/D VGND VGND VPWR VPWR _35923_/Q sky130_fd_sc_hd__dfxtp_1
X_31046_ _35745_/Q _29110_/X _31046_/S VGND VGND VPWR VPWR _31047_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19808_ _34550_/Q _32438_/Q _34422_/Q _34358_/Q _19525_/X _19526_/X VGND VGND VPWR
+ VPWR _19808_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35854_ _35919_/CLK _35854_/D VGND VGND VPWR VPWR _35854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34805_ _34805_/CLK _34805_/D VGND VGND VPWR VPWR _34805_/Q sky130_fd_sc_hd__dfxtp_1
X_19739_ _19739_/A _19739_/B _19739_/C _19739_/D VGND VGND VPWR VPWR _19740_/A sky130_fd_sc_hd__or4_2
X_35785_ _35845_/CLK _35785_/D VGND VGND VPWR VPWR _35785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32997_ _36007_/CLK _32997_/D VGND VGND VPWR VPWR _32997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_886 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22750_ _35081_/Q _35017_/Q _34953_/Q _34889_/Q _22462_/X _22463_/X VGND VGND VPWR
+ VPWR _22750_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31948_ _23345_/X _36173_/Q _31948_/S VGND VGND VPWR VPWR _31949_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_1342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34736_ _34797_/CLK _34736_/D VGND VGND VPWR VPWR _34736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21701_ _33003_/Q _32939_/Q _32875_/Q _32811_/Q _21589_/X _21590_/X VGND VGND VPWR
+ VPWR _21701_/X sky130_fd_sc_hd__mux4_1
X_22681_ _20577_/X _22679_/X _22680_/X _20587_/X VGND VGND VPWR VPWR _22681_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34667_ _34986_/CLK _34667_/D VGND VGND VPWR VPWR _34667_/Q sky130_fd_sc_hd__dfxtp_1
X_31879_ _31948_/S VGND VGND VPWR VPWR _31898_/S sky130_fd_sc_hd__buf_4
XFILLER_53_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24420_ _32710_/Q _24419_/X _24429_/S VGND VGND VPWR VPWR _24421_/A sky130_fd_sc_hd__mux2_1
X_33618_ _34194_/CLK _33618_/D VGND VGND VPWR VPWR _33618_/Q sky130_fd_sc_hd__dfxtp_1
X_21632_ _35817_/Q _32194_/Q _35689_/Q _35625_/Q _21560_/X _21561_/X VGND VGND VPWR
+ VPWR _21632_/X sky130_fd_sc_hd__mux4_1
X_34598_ _35302_/CLK _34598_/D VGND VGND VPWR VPWR _34598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24351_ input28/X VGND VGND VPWR VPWR _24351_/X sky130_fd_sc_hd__buf_6
X_33549_ _35984_/CLK _33549_/D VGND VGND VPWR VPWR _33549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21563_ _35751_/Q _35111_/Q _34471_/Q _33831_/Q _21387_/X _21388_/X VGND VGND VPWR
+ VPWR _21563_/X sky130_fd_sc_hd__mux4_1
X_23302_ _23302_/A VGND VGND VPWR VPWR _32218_/D sky130_fd_sc_hd__clkbuf_1
X_20514_ _20514_/A VGND VGND VPWR VPWR _32139_/D sky130_fd_sc_hd__buf_4
X_27070_ _27070_/A VGND VGND VPWR VPWR _33892_/D sky130_fd_sc_hd__clkbuf_1
X_24282_ _24282_/A VGND VGND VPWR VPWR _32665_/D sky130_fd_sc_hd__clkbuf_1
X_21494_ _35813_/Q _32189_/Q _35685_/Q _35621_/Q _21207_/X _21208_/X VGND VGND VPWR
+ VPWR _21494_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26021_ _25007_/X _33427_/Q _26029_/S VGND VGND VPWR VPWR _26022_/A sky130_fd_sc_hd__mux2_1
X_35219_ _36211_/CLK _35219_/D VGND VGND VPWR VPWR _35219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23233_ _23233_/A VGND VGND VPWR VPWR _32195_/D sky130_fd_sc_hd__clkbuf_1
X_20445_ _20441_/X _20444_/X _20153_/X VGND VGND VPWR VPWR _20453_/C sky130_fd_sc_hd__o21ba_1
XFILLER_101_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36199_ _36200_/CLK _36199_/D VGND VGND VPWR VPWR _36199_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_80_CLK clkbuf_leaf_80_CLK/A VGND VGND VPWR VPWR _35733_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23164_ _23164_/A VGND VGND VPWR VPWR _32165_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20376_ _33031_/Q _32967_/Q _32903_/Q _32839_/Q _18280_/X _18283_/X VGND VGND VPWR
+ VPWR _20376_/X sky130_fd_sc_hd__mux4_1
XFILLER_161_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22115_ _22106_/X _22113_/X _22114_/X VGND VGND VPWR VPWR _22116_/D sky130_fd_sc_hd__o21ba_1
XFILLER_106_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23095_ _23095_/A VGND VGND VPWR VPWR _32144_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27972_ _26826_/X _34319_/Q _27988_/S VGND VGND VPWR VPWR _27973_/A sky130_fd_sc_hd__mux2_1
XTAP_6426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29711_ _29711_/A VGND VGND VPWR VPWR _35112_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26923_ _26922_/X _33838_/Q _26944_/S VGND VGND VPWR VPWR _26924_/A sky130_fd_sc_hd__mux2_1
X_22046_ _33525_/Q _33461_/Q _33397_/Q _33333_/Q _21723_/X _21724_/X VGND VGND VPWR
+ VPWR _22046_/X sky130_fd_sc_hd__mux4_1
XTAP_6459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29642_ _35080_/Q _29231_/X _29644_/S VGND VGND VPWR VPWR _29643_/A sky130_fd_sc_hd__mux2_1
XTAP_5747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26854_ _27018_/S VGND VGND VPWR VPWR _26882_/S sky130_fd_sc_hd__buf_4
XFILLER_76_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25805_ _25805_/A VGND VGND VPWR VPWR _33324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29573_ _35047_/Q _29129_/X _29581_/S VGND VGND VPWR VPWR _29574_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26785_ _26785_/A VGND VGND VPWR VPWR _33788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23997_ _23997_/A VGND VGND VPWR VPWR _32536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28524_ _26844_/X _34581_/Q _28528_/S VGND VGND VPWR VPWR _28525_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25736_ _25736_/A VGND VGND VPWR VPWR _33293_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22948_ input15/X VGND VGND VPWR VPWR _22948_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_43_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28455_ _28455_/A VGND VGND VPWR VPWR _34548_/D sky130_fd_sc_hd__clkbuf_1
X_25667_ _33260_/Q _24338_/X _25685_/S VGND VGND VPWR VPWR _25668_/A sky130_fd_sc_hd__mux2_1
XFILLER_245_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22879_ _22879_/A VGND VGND VPWR VPWR _23075_/S sky130_fd_sc_hd__buf_12
XFILLER_232_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27406_ _34052_/Q _24413_/X _27416_/S VGND VGND VPWR VPWR _27407_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24618_ _24618_/A VGND VGND VPWR VPWR _32798_/D sky130_fd_sc_hd__clkbuf_1
X_28386_ _28386_/A VGND VGND VPWR VPWR _34515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25598_ _25598_/A VGND VGND VPWR VPWR _33229_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27337_ _34019_/Q _24311_/X _27353_/S VGND VGND VPWR VPWR _27338_/A sky130_fd_sc_hd__mux2_1
X_24549_ _24549_/A VGND VGND VPWR VPWR _32767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18070_ _17908_/X _18068_/X _18069_/X _17911_/X VGND VGND VPWR VPWR _18070_/X sky130_fd_sc_hd__a22o_1
X_27268_ _27268_/A VGND VGND VPWR VPWR _33986_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29007_ _34810_/Q _24382_/X _29017_/S VGND VGND VPWR VPWR _29008_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17021_ _17847_/A VGND VGND VPWR VPWR _17021_/X sky130_fd_sc_hd__buf_6
XFILLER_156_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26219_ _25100_/X _33521_/Q _26227_/S VGND VGND VPWR VPWR _26220_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27199_ _27289_/S VGND VGND VPWR VPWR _27218_/S sky130_fd_sc_hd__buf_4
XFILLER_166_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_CLK clkbuf_leaf_73_CLK/A VGND VGND VPWR VPWR _36117_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18972_ _32735_/Q _32671_/Q _32607_/Q _36063_/Q _18866_/X _18650_/X VGND VGND VPWR
+ VPWR _18972_/X sky130_fd_sc_hd__mux4_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ _17700_/X _17921_/X _17922_/X _17703_/X VGND VGND VPWR VPWR _17923_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29909_ _29909_/A VGND VGND VPWR VPWR _35206_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_234_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32920_ _35994_/CLK _32920_/D VGND VGND VPWR VPWR _32920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17854_ _17849_/X _17852_/X _17853_/X VGND VGND VPWR VPWR _17869_/C sky130_fd_sc_hd__o21ba_1
XTAP_6993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16805_ _35042_/Q _34978_/Q _34914_/Q _34850_/Q _16803_/X _16804_/X VGND VGND VPWR
+ VPWR _16805_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32851_ _32978_/CLK _32851_/D VGND VGND VPWR VPWR _32851_/Q sky130_fd_sc_hd__dfxtp_1
X_17785_ _34814_/Q _34750_/Q _34686_/Q _34622_/Q _17641_/X _17642_/X VGND VGND VPWR
+ VPWR _17785_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31802_ _31802_/A VGND VGND VPWR VPWR _36103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19524_ _19449_/X _19522_/X _19523_/X _19452_/X VGND VGND VPWR VPWR _19524_/X sky130_fd_sc_hd__a22o_1
X_35570_ _35955_/CLK _35570_/D VGND VGND VPWR VPWR _35570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16736_ _17956_/A VGND VGND VPWR VPWR _16736_/X sky130_fd_sc_hd__buf_4
X_32782_ _35982_/CLK _32782_/D VGND VGND VPWR VPWR _32782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34521_ _35293_/CLK _34521_/D VGND VGND VPWR VPWR _34521_/Q sky130_fd_sc_hd__dfxtp_1
X_19455_ _34540_/Q _32428_/Q _34412_/Q _34348_/Q _19172_/X _19173_/X VGND VGND VPWR
+ VPWR _19455_/X sky130_fd_sc_hd__mux4_1
X_31733_ _31733_/A VGND VGND VPWR VPWR _36070_/D sky130_fd_sc_hd__clkbuf_1
X_16667_ _17846_/A VGND VGND VPWR VPWR _16667_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_228_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18406_ _18277_/X _18404_/X _18405_/X _18287_/X VGND VGND VPWR VPWR _18406_/X sky130_fd_sc_hd__a22o_1
X_34452_ _35667_/CLK _34452_/D VGND VGND VPWR VPWR _34452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31664_ _36038_/Q input52/X _31670_/S VGND VGND VPWR VPWR _31665_/A sky130_fd_sc_hd__mux2_1
X_19386_ _19386_/A _19386_/B _19386_/C _19386_/D VGND VGND VPWR VPWR _19387_/A sky130_fd_sc_hd__or4_4
XFILLER_188_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16598_ _16496_/X _16596_/X _16597_/X _16499_/X VGND VGND VPWR VPWR _16598_/X sky130_fd_sc_hd__a22o_1
XFILLER_37_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33403_ _33787_/CLK _33403_/D VGND VGND VPWR VPWR _33403_/Q sky130_fd_sc_hd__dfxtp_1
X_30615_ _30615_/A VGND VGND VPWR VPWR _35540_/D sky130_fd_sc_hd__clkbuf_1
X_18337_ _20211_/A VGND VGND VPWR VPWR _18337_/X sky130_fd_sc_hd__clkbuf_4
X_34383_ _34638_/CLK _34383_/D VGND VGND VPWR VPWR _34383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31595_ _36005_/Q input16/X _31607_/S VGND VGND VPWR VPWR _31596_/A sky130_fd_sc_hd__mux2_1
XFILLER_241_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36122_ _36124_/CLK _36122_/D VGND VGND VPWR VPWR _36122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33334_ _34039_/CLK _33334_/D VGND VGND VPWR VPWR _33334_/Q sky130_fd_sc_hd__dfxtp_1
X_18268_ _16044_/X _18266_/X _18267_/X _16054_/X VGND VGND VPWR VPWR _18268_/X sky130_fd_sc_hd__a22o_1
X_30546_ _23264_/X _35508_/Q _30548_/S VGND VGND VPWR VPWR _30547_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36053_ _36116_/CLK _36053_/D VGND VGND VPWR VPWR _36053_/Q sky130_fd_sc_hd__dfxtp_1
X_17219_ _33198_/Q _32558_/Q _35950_/Q _35886_/Q _17074_/X _17075_/X VGND VGND VPWR
+ VPWR _17219_/X sky130_fd_sc_hd__mux4_1
X_33265_ _33520_/CLK _33265_/D VGND VGND VPWR VPWR _33265_/Q sky130_fd_sc_hd__dfxtp_1
X_18199_ _35851_/Q _32231_/Q _35723_/Q _35659_/Q _15989_/X _15991_/X VGND VGND VPWR
+ VPWR _18199_/X sky130_fd_sc_hd__mux4_1
X_30477_ _23102_/X _35475_/Q _30485_/S VGND VGND VPWR VPWR _30478_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_62_CLK clkbuf_leaf_66_CLK/A VGND VGND VPWR VPWR _33512_/CLK sky130_fd_sc_hd__clkbuf_16
X_35004_ _35515_/CLK _35004_/D VGND VGND VPWR VPWR _35004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20230_ _20155_/X _20228_/X _20229_/X _20158_/X VGND VGND VPWR VPWR _20230_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32216_ _35711_/CLK _32216_/D VGND VGND VPWR VPWR _32216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33196_ _35949_/CLK _33196_/D VGND VGND VPWR VPWR _33196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32147_ _36228_/CLK _32147_/D VGND VGND VPWR VPWR _32147_/Q sky130_fd_sc_hd__dfxtp_1
X_20161_ _34560_/Q _32448_/Q _34432_/Q _34368_/Q _19878_/X _19879_/X VGND VGND VPWR
+ VPWR _20161_/X sky130_fd_sc_hd__mux4_1
XFILLER_171_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20092_ _20092_/A _20092_/B _20092_/C _20092_/D VGND VGND VPWR VPWR _20093_/A sky130_fd_sc_hd__or4_1
X_32078_ _34973_/CLK _32078_/D VGND VGND VPWR VPWR _32078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35906_ _35906_/CLK _35906_/D VGND VGND VPWR VPWR _35906_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31029_ _31029_/A VGND VGND VPWR VPWR _35736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23920_ _23000_/X _32501_/Q _23920_/S VGND VGND VPWR VPWR _23921_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35837_ _35837_/CLK _35837_/D VGND VGND VPWR VPWR _35837_/Q sky130_fd_sc_hd__dfxtp_1
X_23851_ _22898_/X _32468_/Q _23857_/S VGND VGND VPWR VPWR _23852_/A sky130_fd_sc_hd__mux2_1
XTAP_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_918 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22802_ _35595_/Q _35531_/Q _35467_/Q _35403_/Q _22556_/X _22557_/X VGND VGND VPWR
+ VPWR _22802_/X sky130_fd_sc_hd__mux4_1
X_26570_ _25019_/X _33687_/Q _26570_/S VGND VGND VPWR VPWR _26571_/A sky130_fd_sc_hd__mux2_1
XANTENNA_608 _18435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_619 _18571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20994_ _32471_/Q _32343_/Q _32023_/Q _35991_/Q _20817_/X _20958_/X VGND VGND VPWR
+ VPWR _20994_/X sky130_fd_sc_hd__mux4_1
X_35768_ _35768_/CLK _35768_/D VGND VGND VPWR VPWR _35768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23782_ _22997_/X _32436_/Q _23784_/S VGND VGND VPWR VPWR _23783_/A sky130_fd_sc_hd__mux2_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25521_ _25521_/A VGND VGND VPWR VPWR _33192_/D sky130_fd_sc_hd__clkbuf_1
X_22733_ _33289_/Q _36169_/Q _33161_/Q _33097_/Q _20628_/X _21757_/A VGND VGND VPWR
+ VPWR _22733_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34719_ _35098_/CLK _34719_/D VGND VGND VPWR VPWR _34719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35699_ _35827_/CLK _35699_/D VGND VGND VPWR VPWR _35699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28240_ _34446_/Q _24244_/X _28258_/S VGND VGND VPWR VPWR _28241_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22664_ _22664_/A VGND VGND VPWR VPWR _36230_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25452_ _25177_/X _33162_/Q _25458_/S VGND VGND VPWR VPWR _25453_/A sky130_fd_sc_hd__mux2_1
XFILLER_240_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24403_ _24403_/A VGND VGND VPWR VPWR _32704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21615_ _21615_/A VGND VGND VPWR VPWR _36200_/D sky130_fd_sc_hd__clkbuf_1
X_28171_ _28171_/A VGND VGND VPWR VPWR _34413_/D sky130_fd_sc_hd__clkbuf_1
X_22595_ _22595_/A VGND VGND VPWR VPWR _22595_/X sky130_fd_sc_hd__buf_4
XFILLER_142_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25383_ _25075_/X _33129_/Q _25387_/S VGND VGND VPWR VPWR _25384_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27122_ _27122_/A VGND VGND VPWR VPWR _33917_/D sky130_fd_sc_hd__clkbuf_1
X_21546_ _33767_/Q _33703_/Q _33639_/Q _33575_/Q _21443_/X _21444_/X VGND VGND VPWR
+ VPWR _21546_/X sky130_fd_sc_hd__mux4_1
X_24334_ _24334_/A VGND VGND VPWR VPWR _32682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24265_ _32660_/Q _24264_/X _24274_/S VGND VGND VPWR VPWR _24266_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27053_ _27053_/A VGND VGND VPWR VPWR _33884_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21477_ _21471_/X _21476_/X _21408_/X VGND VGND VPWR VPWR _21478_/D sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_53_CLK clkbuf_leaf_57_CLK/A VGND VGND VPWR VPWR _35994_/CLK sky130_fd_sc_hd__clkbuf_16
X_26004_ _26004_/A VGND VGND VPWR VPWR _33419_/D sky130_fd_sc_hd__clkbuf_1
X_23216_ _23216_/A VGND VGND VPWR VPWR _32189_/D sky130_fd_sc_hd__clkbuf_1
X_20428_ _33545_/Q _33481_/Q _33417_/Q _33353_/Q _20129_/X _20130_/X VGND VGND VPWR
+ VPWR _20428_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24196_ _24196_/A VGND VGND VPWR VPWR _32630_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23147_ _23147_/A VGND VGND VPWR VPWR _32161_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20359_ _34566_/Q _32454_/Q _34438_/Q _34374_/Q _20231_/X _20232_/X VGND VGND VPWR
+ VPWR _20359_/X sky130_fd_sc_hd__mux4_1
XFILLER_175_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1007 _17862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1018 _17858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27955_ _27955_/A VGND VGND VPWR VPWR _34311_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23078_ input87/X VGND VGND VPWR VPWR _30329_/B sky130_fd_sc_hd__buf_4
XTAP_5500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1029 _17865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26906_ input20/X VGND VGND VPWR VPWR _26906_/X sky130_fd_sc_hd__clkbuf_4
X_22029_ _33204_/Q _32564_/Q _35956_/Q _35892_/Q _22027_/X _22028_/X VGND VGND VPWR
+ VPWR _22029_/X sky130_fd_sc_hd__mux4_1
XTAP_6289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27886_ _27886_/A VGND VGND VPWR VPWR _34278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29625_ _29652_/S VGND VGND VPWR VPWR _29644_/S sky130_fd_sc_hd__buf_4
XTAP_5577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26837_ _26837_/A VGND VGND VPWR VPWR _33810_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17570_ _17347_/X _17568_/X _17569_/X _17350_/X VGND VGND VPWR VPWR _17570_/X sky130_fd_sc_hd__a22o_1
X_29556_ _35039_/Q _29104_/X _29560_/S VGND VGND VPWR VPWR _29557_/A sky130_fd_sc_hd__mux2_1
XTAP_4898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26768_ _26768_/A VGND VGND VPWR VPWR _33780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_217_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28507_ _28507_/A VGND VGND VPWR VPWR _34573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16521_ _34522_/Q _32410_/Q _34394_/Q _34330_/Q _16519_/X _16520_/X VGND VGND VPWR
+ VPWR _16521_/X sky130_fd_sc_hd__mux4_1
X_25719_ _33285_/Q _24416_/X _25727_/S VGND VGND VPWR VPWR _25720_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29487_ _29487_/A VGND VGND VPWR VPWR _35006_/D sky130_fd_sc_hd__clkbuf_1
X_26699_ _26699_/A VGND VGND VPWR VPWR _33747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19240_ _34534_/Q _32422_/Q _34406_/Q _34342_/Q _19172_/X _19173_/X VGND VGND VPWR
+ VPWR _19240_/X sky130_fd_sc_hd__mux4_1
XFILLER_204_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28438_ _26915_/X _34540_/Q _28456_/S VGND VGND VPWR VPWR _28439_/A sky130_fd_sc_hd__mux2_1
X_16452_ _35032_/Q _34968_/Q _34904_/Q _34840_/Q _16450_/X _16451_/X VGND VGND VPWR
+ VPWR _16452_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19171_ _19096_/X _19169_/X _19170_/X _19099_/X VGND VGND VPWR VPWR _19171_/X sky130_fd_sc_hd__a22o_1
X_28369_ _34508_/Q _24437_/X _28371_/S VGND VGND VPWR VPWR _28370_/A sky130_fd_sc_hd__mux2_1
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16383_ _17956_/A VGND VGND VPWR VPWR _16383_/X sky130_fd_sc_hd__buf_6
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18122_ _18118_/X _18121_/X _17867_/X VGND VGND VPWR VPWR _18123_/D sky130_fd_sc_hd__o21ba_1
X_30400_ _30400_/A VGND VGND VPWR VPWR _35438_/D sky130_fd_sc_hd__clkbuf_1
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31380_ _31380_/A VGND VGND VPWR VPWR _35903_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18053_ _33222_/Q _32582_/Q _35974_/Q _35910_/Q _17780_/X _17781_/X VGND VGND VPWR
+ VPWR _18053_/X sky130_fd_sc_hd__mux4_1
X_30331_ _30463_/S VGND VGND VPWR VPWR _30350_/S sky130_fd_sc_hd__buf_4
XFILLER_172_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_44_CLK clkbuf_6_6__f_CLK/X VGND VGND VPWR VPWR _36125_/CLK sky130_fd_sc_hd__clkbuf_16
X_17004_ _16998_/X _17003_/X _16794_/X VGND VGND VPWR VPWR _17014_/C sky130_fd_sc_hd__o21ba_1
XANTENNA_4 _32114_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33050_ _36124_/CLK _33050_/D VGND VGND VPWR VPWR _33050_/Q sky130_fd_sc_hd__dfxtp_1
X_30262_ _30262_/A VGND VGND VPWR VPWR _35373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32001_ _34202_/CLK _32001_/D VGND VGND VPWR VPWR _32001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30193_ _30193_/A VGND VGND VPWR VPWR _35341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18955_ _35294_/Q _35230_/Q _35166_/Q _32286_/Q _18953_/X _18954_/X VGND VGND VPWR
+ VPWR _18955_/X sky130_fd_sc_hd__mux4_1
XFILLER_86_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17906_ _17906_/A VGND VGND VPWR VPWR _17906_/X sky130_fd_sc_hd__buf_4
X_18886_ _18743_/X _18884_/X _18885_/X _18746_/X VGND VGND VPWR VPWR _18886_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33952_ _36124_/CLK _33952_/D VGND VGND VPWR VPWR _33952_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32903_ _34752_/CLK _32903_/D VGND VGND VPWR VPWR _32903_/Q sky130_fd_sc_hd__dfxtp_1
X_17837_ _33280_/Q _36160_/Q _33152_/Q _33088_/Q _17764_/X _17765_/X VGND VGND VPWR
+ VPWR _17837_/X sky130_fd_sc_hd__mux4_1
X_33883_ _34202_/CLK _33883_/D VGND VGND VPWR VPWR _33883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32834_ _32962_/CLK _32834_/D VGND VGND VPWR VPWR _32834_/Q sky130_fd_sc_hd__dfxtp_1
X_35622_ _35814_/CLK _35622_/D VGND VGND VPWR VPWR _35622_/Q sky130_fd_sc_hd__dfxtp_1
X_17768_ _17761_/X _17763_/X _17766_/X _17767_/X VGND VGND VPWR VPWR _17768_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_1022 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16719_ _16641_/X _16717_/X _16718_/X _16644_/X VGND VGND VPWR VPWR _16719_/X sky130_fd_sc_hd__a22o_1
X_19507_ _19501_/X _19506_/X _19428_/X VGND VGND VPWR VPWR _19531_/A sky130_fd_sc_hd__o21ba_1
X_32765_ _36092_/CLK _32765_/D VGND VGND VPWR VPWR _32765_/Q sky130_fd_sc_hd__dfxtp_1
X_35553_ _35809_/CLK _35553_/D VGND VGND VPWR VPWR _35553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17699_ _17693_/X _17698_/X _17489_/X _17490_/X VGND VGND VPWR VPWR _17720_/B sky130_fd_sc_hd__o211a_1
Xclkbuf_6_56__f_CLK clkbuf_5_28_0_CLK/X VGND VGND VPWR VPWR clkbuf_6_56__f_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34504_ _35847_/CLK _34504_/D VGND VGND VPWR VPWR _34504_/Q sky130_fd_sc_hd__dfxtp_1
X_19438_ _19432_/X _19435_/X _19436_/X _19437_/X VGND VGND VPWR VPWR _19463_/B sky130_fd_sc_hd__o211a_1
X_31716_ _31716_/A VGND VGND VPWR VPWR _36062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35484_ _35932_/CLK _35484_/D VGND VGND VPWR VPWR _35484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32696_ _36088_/CLK _32696_/D VGND VGND VPWR VPWR _32696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34435_ _34947_/CLK _34435_/D VGND VGND VPWR VPWR _34435_/Q sky130_fd_sc_hd__dfxtp_1
X_31647_ _36030_/Q input43/X _31649_/S VGND VGND VPWR VPWR _31648_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19369_ _19362_/X _19368_/X _19083_/X _19084_/X VGND VGND VPWR VPWR _19386_/B sky130_fd_sc_hd__o211a_1
XFILLER_241_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21400_ _21396_/X _21397_/X _21398_/X _21399_/X VGND VGND VPWR VPWR _21400_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22380_ _22531_/A VGND VGND VPWR VPWR _22380_/X sky130_fd_sc_hd__buf_6
X_34366_ _35581_/CLK _34366_/D VGND VGND VPWR VPWR _34366_/Q sky130_fd_sc_hd__dfxtp_1
X_31578_ _35997_/Q input7/X _31586_/S VGND VGND VPWR VPWR _31579_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36105_ _36105_/CLK _36105_/D VGND VGND VPWR VPWR _36105_/Q sky130_fd_sc_hd__dfxtp_1
X_33317_ _33507_/CLK _33317_/D VGND VGND VPWR VPWR _33317_/Q sky130_fd_sc_hd__dfxtp_1
X_21331_ _21048_/X _21329_/X _21330_/X _21053_/X VGND VGND VPWR VPWR _21331_/X sky130_fd_sc_hd__a22o_1
X_30529_ _30598_/S VGND VGND VPWR VPWR _30548_/S sky130_fd_sc_hd__buf_6
X_34297_ _34297_/CLK _34297_/D VGND VGND VPWR VPWR _34297_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_35_CLK clkbuf_6_7__f_CLK/X VGND VGND VPWR VPWR _34145_/CLK sky130_fd_sc_hd__clkbuf_16
X_24050_ _22991_/X _32562_/Q _24056_/S VGND VGND VPWR VPWR _24051_/A sky130_fd_sc_hd__mux2_1
X_36036_ _36037_/CLK _36036_/D VGND VGND VPWR VPWR _36036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21262_ _21262_/A VGND VGND VPWR VPWR _36190_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33248_ _36128_/CLK _33248_/D VGND VGND VPWR VPWR _33248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23001_ _23000_/X _32053_/Q _23001_/S VGND VGND VPWR VPWR _23002_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20213_ _20207_/X _20212_/X _20134_/X VGND VGND VPWR VPWR _20237_/A sky130_fd_sc_hd__o21ba_1
XFILLER_144_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33179_ _35931_/CLK _33179_/D VGND VGND VPWR VPWR _33179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21193_ _33757_/Q _33693_/Q _33629_/Q _33565_/Q _21090_/X _21091_/X VGND VGND VPWR
+ VPWR _21193_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20144_ _20138_/X _20141_/X _20142_/X _20143_/X VGND VGND VPWR VPWR _20169_/B sky130_fd_sc_hd__o211a_1
XFILLER_213_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27740_ _27740_/A VGND VGND VPWR VPWR _34209_/D sky130_fd_sc_hd__clkbuf_1
X_20075_ _20068_/X _20074_/X _19789_/X _19790_/X VGND VGND VPWR VPWR _20092_/B sky130_fd_sc_hd__o211a_1
X_24952_ _23022_/X _32956_/Q _24958_/S VGND VGND VPWR VPWR _24953_/A sky130_fd_sc_hd__mux2_1
XTAP_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23903_ _23903_/A VGND VGND VPWR VPWR _32492_/D sky130_fd_sc_hd__clkbuf_1
X_27671_ _27671_/A VGND VGND VPWR VPWR _34176_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24883_ _22920_/X _32923_/Q _24895_/S VGND VGND VPWR VPWR _24884_/A sky130_fd_sc_hd__mux2_1
XTAP_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29410_ _29410_/A VGND VGND VPWR VPWR _34969_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26622_ _26622_/A VGND VGND VPWR VPWR _33711_/D sky130_fd_sc_hd__clkbuf_1
X_23834_ _23074_/X _32461_/Q _23834_/S VGND VGND VPWR VPWR _23835_/A sky130_fd_sc_hd__mux2_1
XTAP_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_405 _36211_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_416 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29341_ _23280_/X _34937_/Q _29353_/S VGND VGND VPWR VPWR _29342_/A sky130_fd_sc_hd__mux2_1
XANTENNA_427 _31989_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26553_ _26553_/A VGND VGND VPWR VPWR _33678_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_438 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20977_ _35030_/Q _34966_/Q _34902_/Q _34838_/Q _20692_/X _20694_/X VGND VGND VPWR
+ VPWR _20977_/X sky130_fd_sc_hd__mux4_1
X_23765_ _23834_/S VGND VGND VPWR VPWR _23784_/S sky130_fd_sc_hd__buf_6
XFILLER_82_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_449 _31990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25504_ _25504_/A VGND VGND VPWR VPWR _33184_/D sky130_fd_sc_hd__clkbuf_1
X_22716_ _34824_/Q _34760_/Q _34696_/Q _34632_/Q _22594_/X _22595_/X VGND VGND VPWR
+ VPWR _22716_/X sky130_fd_sc_hd__mux4_1
XFILLER_15_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29272_ _23117_/X _34904_/Q _29290_/S VGND VGND VPWR VPWR _29273_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26484_ _26484_/A VGND VGND VPWR VPWR _33646_/D sky130_fd_sc_hd__clkbuf_1
X_23696_ _32397_/Q _23345_/X _23696_/S VGND VGND VPWR VPWR _23697_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28223_ _28223_/A VGND VGND VPWR VPWR _34438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25435_ _25435_/A VGND VGND VPWR VPWR _33153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_213_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22647_ _22369_/X _22645_/X _22646_/X _22373_/X VGND VGND VPWR VPWR _22647_/X sky130_fd_sc_hd__a22o_1
XFILLER_201_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28154_ _28154_/A VGND VGND VPWR VPWR _34405_/D sky130_fd_sc_hd__clkbuf_1
X_22578_ _22578_/A VGND VGND VPWR VPWR _22578_/X sky130_fd_sc_hd__buf_6
XFILLER_16_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25366_ _25050_/X _33121_/Q _25366_/S VGND VGND VPWR VPWR _25367_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27105_ _27105_/A VGND VGND VPWR VPWR _33909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24317_ input16/X VGND VGND VPWR VPWR _24317_/X sky130_fd_sc_hd__buf_4
X_28085_ _26993_/X _34373_/Q _28093_/S VGND VGND VPWR VPWR _28086_/A sky130_fd_sc_hd__mux2_1
X_21529_ _35750_/Q _35110_/Q _34470_/Q _33830_/Q _21387_/X _21388_/X VGND VGND VPWR
+ VPWR _21529_/X sky130_fd_sc_hd__mux4_1
X_25297_ _25297_/A VGND VGND VPWR VPWR _33088_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_26_CLK clkbuf_6_5__f_CLK/X VGND VGND VPWR VPWR _34010_/CLK sky130_fd_sc_hd__clkbuf_16
X_27036_ _27036_/A VGND VGND VPWR VPWR _33876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24248_ _24248_/A VGND VGND VPWR VPWR _32654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24179_ _24179_/A VGND VGND VPWR VPWR _32622_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28987_ _28987_/A VGND VGND VPWR VPWR _34800_/D sky130_fd_sc_hd__clkbuf_1
XTAP_6042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput96 _31965_/Q VGND VGND VPWR VPWR D1[15] sky130_fd_sc_hd__buf_2
XTAP_6064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18740_ _18593_/X _18738_/X _18739_/X _18596_/X VGND VGND VPWR VPWR _18740_/X sky130_fd_sc_hd__a22o_1
XTAP_5330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27938_ _27938_/A VGND VGND VPWR VPWR _34303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18671_ _18593_/X _18667_/X _18670_/X _18596_/X VGND VGND VPWR VPWR _18671_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27869_ _27869_/A VGND VGND VPWR VPWR _34270_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17622_ _34042_/Q _33978_/Q _33914_/Q _32250_/Q _17373_/X _17374_/X VGND VGND VPWR
+ VPWR _17622_/X sky130_fd_sc_hd__mux4_1
XTAP_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29608_ _29608_/A VGND VGND VPWR VPWR _35063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30880_ _35666_/Q _29064_/X _30890_/S VGND VGND VPWR VPWR _30881_/A sky130_fd_sc_hd__mux2_1
XTAP_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17553_ _17906_/A VGND VGND VPWR VPWR _17553_/X sky130_fd_sc_hd__clkbuf_4
X_29539_ _35031_/Q _29079_/X _29539_/S VGND VGND VPWR VPWR _29540_/A sky130_fd_sc_hd__mux2_1
XTAP_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_950 _29652_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16504_ _16349_/X _16502_/X _16503_/X _16355_/X VGND VGND VPWR VPWR _16504_/X sky130_fd_sc_hd__a22o_1
X_32550_ _35942_/CLK _32550_/D VGND VGND VPWR VPWR _32550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_961 _30057_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_972 _31813_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17484_ _33270_/Q _36150_/Q _33142_/Q _33078_/Q _17411_/X _17412_/X VGND VGND VPWR
+ VPWR _17484_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_983 _17795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_994 _17860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31501_ _31501_/A VGND VGND VPWR VPWR _35960_/D sky130_fd_sc_hd__clkbuf_1
X_19223_ _20282_/A VGND VGND VPWR VPWR _19223_/X sky130_fd_sc_hd__buf_6
XFILLER_108_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16435_ _17995_/A VGND VGND VPWR VPWR _16435_/X sky130_fd_sc_hd__clkbuf_4
X_32481_ _36001_/CLK _32481_/D VGND VGND VPWR VPWR _32481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34220_ _35315_/CLK _34220_/D VGND VGND VPWR VPWR _34220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31432_ _31543_/S VGND VGND VPWR VPWR _31451_/S sky130_fd_sc_hd__buf_4
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19154_ _19148_/X _19153_/X _19075_/X VGND VGND VPWR VPWR _19178_/A sky130_fd_sc_hd__o21ba_1
X_16366_ _16288_/X _16364_/X _16365_/X _16291_/X VGND VGND VPWR VPWR _16366_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18105_ _32520_/Q _32392_/Q _32072_/Q _36040_/Q _17982_/X _17007_/A VGND VGND VPWR
+ VPWR _18105_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34151_ _34279_/CLK _34151_/D VGND VGND VPWR VPWR _34151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19085_ _19079_/X _19082_/X _19083_/X _19084_/X VGND VGND VPWR VPWR _19110_/B sky130_fd_sc_hd__o211a_1
X_31363_ _35895_/Q input36/X _31379_/S VGND VGND VPWR VPWR _31364_/A sky130_fd_sc_hd__mux2_1
X_16297_ _16293_/X _16294_/X _16295_/X _16296_/X VGND VGND VPWR VPWR _16297_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_17_CLK clkbuf_6_6__f_CLK/X VGND VGND VPWR VPWR _34271_/CLK sky130_fd_sc_hd__clkbuf_16
X_33102_ _36114_/CLK _33102_/D VGND VGND VPWR VPWR _33102_/Q sky130_fd_sc_hd__dfxtp_1
X_18036_ _34310_/Q _34246_/Q _34182_/Q _34118_/Q _17795_/X _17796_/X VGND VGND VPWR
+ VPWR _18036_/X sky130_fd_sc_hd__mux4_1
X_30314_ _30314_/A VGND VGND VPWR VPWR _35398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34082_ _34146_/CLK _34082_/D VGND VGND VPWR VPWR _34082_/Q sky130_fd_sc_hd__dfxtp_1
X_31294_ _31294_/A VGND VGND VPWR VPWR _35862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33033_ _36169_/CLK _33033_/D VGND VGND VPWR VPWR _33033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30245_ _30245_/A VGND VGND VPWR VPWR _35365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1013 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30176_ _35333_/Q _29222_/X _30184_/S VGND VGND VPWR VPWR _30177_/A sky130_fd_sc_hd__mux2_1
X_19987_ _33532_/Q _33468_/Q _33404_/Q _33340_/Q _19776_/X _19777_/X VGND VGND VPWR
+ VPWR _19987_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18938_ _32990_/Q _32926_/Q _32862_/Q _32798_/Q _18936_/X _18937_/X VGND VGND VPWR
+ VPWR _18938_/X sky130_fd_sc_hd__mux4_1
.ends

