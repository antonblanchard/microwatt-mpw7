VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM32_1RW1R
  CLASS BLOCK ;
  FOREIGN RAM32_1RW1R ;
  ORIGIN 0.000 0.000 ;
  SIZE 1173.460 BY 185.440 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 124.480 1173.460 125.080 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 137.400 1173.460 138.000 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 150.320 1173.460 150.920 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 163.240 1173.460 163.840 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 176.160 1173.460 176.760 ;
    END
  END A0[4]
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 2.000 40.080 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 2.000 66.600 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 2.000 93.120 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 2.000 119.640 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 2.000 146.160 ;
    END
  END A1[4]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 2.000 13.560 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 0.000 290.630 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 0.000 326.510 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 0.000 434.150 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 0.000 470.030 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 0.000 523.850 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 0.000 541.790 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 0.000 559.730 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 0.000 577.670 2.000 ;
    END
  END Di0[31]
  PIN Di0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 2.000 ;
    END
  END Di0[32]
  PIN Di0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 2.000 ;
    END
  END Di0[33]
  PIN Di0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 2.000 ;
    END
  END Di0[34]
  PIN Di0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.150 0.000 649.430 2.000 ;
    END
  END Di0[35]
  PIN Di0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 2.000 ;
    END
  END Di0[36]
  PIN Di0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 0.000 685.310 2.000 ;
    END
  END Di0[37]
  PIN Di0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.970 0.000 703.250 2.000 ;
    END
  END Di0[38]
  PIN Di0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 0.000 721.190 2.000 ;
    END
  END Di0[39]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 2.000 ;
    END
  END Di0[3]
  PIN Di0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 0.000 739.130 2.000 ;
    END
  END Di0[40]
  PIN Di0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 2.000 ;
    END
  END Di0[41]
  PIN Di0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 0.000 775.010 2.000 ;
    END
  END Di0[42]
  PIN Di0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.670 0.000 792.950 2.000 ;
    END
  END Di0[43]
  PIN Di0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.610 0.000 810.890 2.000 ;
    END
  END Di0[44]
  PIN Di0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 0.000 828.830 2.000 ;
    END
  END Di0[45]
  PIN Di0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 0.000 846.770 2.000 ;
    END
  END Di0[46]
  PIN Di0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.430 0.000 864.710 2.000 ;
    END
  END Di0[47]
  PIN Di0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 2.000 ;
    END
  END Di0[48]
  PIN Di0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.310 0.000 900.590 2.000 ;
    END
  END Di0[49]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 2.000 ;
    END
  END Di0[4]
  PIN Di0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 0.000 918.530 2.000 ;
    END
  END Di0[50]
  PIN Di0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.190 0.000 936.470 2.000 ;
    END
  END Di0[51]
  PIN Di0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.130 0.000 954.410 2.000 ;
    END
  END Di0[52]
  PIN Di0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.070 0.000 972.350 2.000 ;
    END
  END Di0[53]
  PIN Di0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.010 0.000 990.290 2.000 ;
    END
  END Di0[54]
  PIN Di0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 0.000 1008.230 2.000 ;
    END
  END Di0[55]
  PIN Di0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.890 0.000 1026.170 2.000 ;
    END
  END Di0[56]
  PIN Di0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.830 0.000 1044.110 2.000 ;
    END
  END Di0[57]
  PIN Di0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.770 0.000 1062.050 2.000 ;
    END
  END Di0[58]
  PIN Di0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.710 0.000 1079.990 2.000 ;
    END
  END Di0[59]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 2.000 ;
    END
  END Di0[5]
  PIN Di0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.650 0.000 1097.930 2.000 ;
    END
  END Di0[60]
  PIN Di0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.590 0.000 1115.870 2.000 ;
    END
  END Di0[61]
  PIN Di0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.530 0.000 1133.810 2.000 ;
    END
  END Di0[62]
  PIN Di0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.470 0.000 1151.750 2.000 ;
    END
  END Di0[63]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 183.440 31.650 185.440 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 183.440 119.050 185.440 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 183.440 136.530 185.440 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 183.440 154.010 185.440 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 183.440 171.490 185.440 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 183.440 188.970 185.440 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 183.440 206.450 185.440 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 183.440 223.930 185.440 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 183.440 241.410 185.440 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 183.440 258.890 185.440 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 183.440 276.370 185.440 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 183.440 40.390 185.440 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 183.440 293.850 185.440 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 183.440 302.590 185.440 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 183.440 311.330 185.440 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 183.440 320.070 185.440 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 183.440 328.810 185.440 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 183.440 337.550 185.440 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 183.440 346.290 185.440 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 183.440 355.030 185.440 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 183.440 363.770 185.440 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 183.440 372.510 185.440 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 183.440 49.130 185.440 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 183.440 381.250 185.440 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 183.440 389.990 185.440 ;
    END
  END Do0[31]
  PIN Do0[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 183.440 398.730 185.440 ;
    END
  END Do0[32]
  PIN Do0[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 183.440 407.470 185.440 ;
    END
  END Do0[33]
  PIN Do0[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 183.440 416.210 185.440 ;
    END
  END Do0[34]
  PIN Do0[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 183.440 424.950 185.440 ;
    END
  END Do0[35]
  PIN Do0[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 183.440 433.690 185.440 ;
    END
  END Do0[36]
  PIN Do0[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 183.440 442.430 185.440 ;
    END
  END Do0[37]
  PIN Do0[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 183.440 451.170 185.440 ;
    END
  END Do0[38]
  PIN Do0[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 183.440 459.910 185.440 ;
    END
  END Do0[39]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 183.440 57.870 185.440 ;
    END
  END Do0[3]
  PIN Do0[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 183.440 468.650 185.440 ;
    END
  END Do0[40]
  PIN Do0[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 183.440 477.390 185.440 ;
    END
  END Do0[41]
  PIN Do0[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 183.440 486.130 185.440 ;
    END
  END Do0[42]
  PIN Do0[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 183.440 494.870 185.440 ;
    END
  END Do0[43]
  PIN Do0[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 183.440 503.610 185.440 ;
    END
  END Do0[44]
  PIN Do0[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 183.440 512.350 185.440 ;
    END
  END Do0[45]
  PIN Do0[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 183.440 521.090 185.440 ;
    END
  END Do0[46]
  PIN Do0[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 183.440 529.830 185.440 ;
    END
  END Do0[47]
  PIN Do0[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 183.440 538.570 185.440 ;
    END
  END Do0[48]
  PIN Do0[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 183.440 547.310 185.440 ;
    END
  END Do0[49]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 183.440 66.610 185.440 ;
    END
  END Do0[4]
  PIN Do0[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 183.440 556.050 185.440 ;
    END
  END Do0[50]
  PIN Do0[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 183.440 564.790 185.440 ;
    END
  END Do0[51]
  PIN Do0[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 183.440 573.530 185.440 ;
    END
  END Do0[52]
  PIN Do0[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 183.440 582.270 185.440 ;
    END
  END Do0[53]
  PIN Do0[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 183.440 591.010 185.440 ;
    END
  END Do0[54]
  PIN Do0[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 183.440 599.750 185.440 ;
    END
  END Do0[55]
  PIN Do0[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 183.440 608.490 185.440 ;
    END
  END Do0[56]
  PIN Do0[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 183.440 617.230 185.440 ;
    END
  END Do0[57]
  PIN Do0[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 183.440 625.970 185.440 ;
    END
  END Do0[58]
  PIN Do0[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 183.440 634.710 185.440 ;
    END
  END Do0[59]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 183.440 75.350 185.440 ;
    END
  END Do0[5]
  PIN Do0[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 183.440 643.450 185.440 ;
    END
  END Do0[60]
  PIN Do0[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 183.440 652.190 185.440 ;
    END
  END Do0[61]
  PIN Do0[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 183.440 660.930 185.440 ;
    END
  END Do0[62]
  PIN Do0[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 183.440 669.670 185.440 ;
    END
  END Do0[63]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 183.440 84.090 185.440 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 183.440 92.830 185.440 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 183.440 101.570 185.440 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 183.440 110.310 185.440 ;
    END
  END Do0[9]
  PIN Do1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 183.440 127.790 185.440 ;
    END
  END Do1[0]
  PIN Do1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 183.440 678.410 185.440 ;
    END
  END Do1[10]
  PIN Do1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 183.440 687.150 185.440 ;
    END
  END Do1[11]
  PIN Do1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 183.440 695.890 185.440 ;
    END
  END Do1[12]
  PIN Do1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 183.440 704.630 185.440 ;
    END
  END Do1[13]
  PIN Do1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 183.440 713.370 185.440 ;
    END
  END Do1[14]
  PIN Do1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 183.440 722.110 185.440 ;
    END
  END Do1[15]
  PIN Do1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 183.440 730.850 185.440 ;
    END
  END Do1[16]
  PIN Do1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 183.440 739.590 185.440 ;
    END
  END Do1[17]
  PIN Do1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 183.440 748.330 185.440 ;
    END
  END Do1[18]
  PIN Do1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 183.440 757.070 185.440 ;
    END
  END Do1[19]
  PIN Do1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 183.440 145.270 185.440 ;
    END
  END Do1[1]
  PIN Do1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 183.440 765.810 185.440 ;
    END
  END Do1[20]
  PIN Do1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 183.440 774.550 185.440 ;
    END
  END Do1[21]
  PIN Do1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 183.440 783.290 185.440 ;
    END
  END Do1[22]
  PIN Do1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.750 183.440 792.030 185.440 ;
    END
  END Do1[23]
  PIN Do1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 183.440 800.770 185.440 ;
    END
  END Do1[24]
  PIN Do1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.230 183.440 809.510 185.440 ;
    END
  END Do1[25]
  PIN Do1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 183.440 818.250 185.440 ;
    END
  END Do1[26]
  PIN Do1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 183.440 826.990 185.440 ;
    END
  END Do1[27]
  PIN Do1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.450 183.440 835.730 185.440 ;
    END
  END Do1[28]
  PIN Do1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.190 183.440 844.470 185.440 ;
    END
  END Do1[29]
  PIN Do1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 183.440 162.750 185.440 ;
    END
  END Do1[2]
  PIN Do1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.930 183.440 853.210 185.440 ;
    END
  END Do1[30]
  PIN Do1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.670 183.440 861.950 185.440 ;
    END
  END Do1[31]
  PIN Do1[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 183.440 870.690 185.440 ;
    END
  END Do1[32]
  PIN Do1[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 183.440 879.430 185.440 ;
    END
  END Do1[33]
  PIN Do1[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 183.440 888.170 185.440 ;
    END
  END Do1[34]
  PIN Do1[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.630 183.440 896.910 185.440 ;
    END
  END Do1[35]
  PIN Do1[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.370 183.440 905.650 185.440 ;
    END
  END Do1[36]
  PIN Do1[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.110 183.440 914.390 185.440 ;
    END
  END Do1[37]
  PIN Do1[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.850 183.440 923.130 185.440 ;
    END
  END Do1[38]
  PIN Do1[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.590 183.440 931.870 185.440 ;
    END
  END Do1[39]
  PIN Do1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 183.440 180.230 185.440 ;
    END
  END Do1[3]
  PIN Do1[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 183.440 940.610 185.440 ;
    END
  END Do1[40]
  PIN Do1[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 183.440 949.350 185.440 ;
    END
  END Do1[41]
  PIN Do1[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.810 183.440 958.090 185.440 ;
    END
  END Do1[42]
  PIN Do1[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 183.440 966.830 185.440 ;
    END
  END Do1[43]
  PIN Do1[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.290 183.440 975.570 185.440 ;
    END
  END Do1[44]
  PIN Do1[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.030 183.440 984.310 185.440 ;
    END
  END Do1[45]
  PIN Do1[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.770 183.440 993.050 185.440 ;
    END
  END Do1[46]
  PIN Do1[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 183.440 1001.790 185.440 ;
    END
  END Do1[47]
  PIN Do1[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.250 183.440 1010.530 185.440 ;
    END
  END Do1[48]
  PIN Do1[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.990 183.440 1019.270 185.440 ;
    END
  END Do1[49]
  PIN Do1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 183.440 197.710 185.440 ;
    END
  END Do1[4]
  PIN Do1[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.730 183.440 1028.010 185.440 ;
    END
  END Do1[50]
  PIN Do1[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.470 183.440 1036.750 185.440 ;
    END
  END Do1[51]
  PIN Do1[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.210 183.440 1045.490 185.440 ;
    END
  END Do1[52]
  PIN Do1[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.950 183.440 1054.230 185.440 ;
    END
  END Do1[53]
  PIN Do1[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 183.440 1062.970 185.440 ;
    END
  END Do1[54]
  PIN Do1[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.430 183.440 1071.710 185.440 ;
    END
  END Do1[55]
  PIN Do1[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.170 183.440 1080.450 185.440 ;
    END
  END Do1[56]
  PIN Do1[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.910 183.440 1089.190 185.440 ;
    END
  END Do1[57]
  PIN Do1[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.650 183.440 1097.930 185.440 ;
    END
  END Do1[58]
  PIN Do1[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.390 183.440 1106.670 185.440 ;
    END
  END Do1[59]
  PIN Do1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 183.440 215.190 185.440 ;
    END
  END Do1[5]
  PIN Do1[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.130 183.440 1115.410 185.440 ;
    END
  END Do1[60]
  PIN Do1[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 183.440 1124.150 185.440 ;
    END
  END Do1[61]
  PIN Do1[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.610 183.440 1132.890 185.440 ;
    END
  END Do1[62]
  PIN Do1[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.350 183.440 1141.630 185.440 ;
    END
  END Do1[63]
  PIN Do1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 183.440 232.670 185.440 ;
    END
  END Do1[6]
  PIN Do1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 183.440 250.150 185.440 ;
    END
  END Do1[7]
  PIN Do1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 183.440 267.630 185.440 ;
    END
  END Do1[8]
  PIN Do1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 183.440 285.110 185.440 ;
    END
  END Do1[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 8.200 1173.460 8.800 ;
    END
  END EN0
  PIN EN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 2.000 172.680 ;
    END
  END EN1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.210 2.480 99.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 276.210 2.480 279.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 456.210 2.480 459.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.210 2.480 639.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 816.210 2.480 819.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.210 2.480 999.310 182.480 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 6.210 2.480 9.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 186.210 2.480 189.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 366.210 2.480 369.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.210 2.480 549.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 726.210 2.480 729.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 906.210 2.480 909.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1086.210 2.480 1089.310 182.480 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 21.120 1173.460 21.720 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 34.040 1173.460 34.640 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 46.960 1173.460 47.560 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 59.880 1173.460 60.480 ;
    END
  END WE0[3]
  PIN WE0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 72.800 1173.460 73.400 ;
    END
  END WE0[4]
  PIN WE0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 85.720 1173.460 86.320 ;
    END
  END WE0[5]
  PIN WE0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 98.640 1173.460 99.240 ;
    END
  END WE0[6]
  PIN WE0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 111.560 1173.460 112.160 ;
    END
  END WE0[7]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 1170.700 98.005 ;
      LAYER met1 ;
        RECT 1.450 0.040 1170.700 182.480 ;
      LAYER met2 ;
        RECT 1.470 183.160 31.090 184.805 ;
        RECT 31.930 183.160 39.830 184.805 ;
        RECT 40.670 183.160 48.570 184.805 ;
        RECT 49.410 183.160 57.310 184.805 ;
        RECT 58.150 183.160 66.050 184.805 ;
        RECT 66.890 183.160 74.790 184.805 ;
        RECT 75.630 183.160 83.530 184.805 ;
        RECT 84.370 183.160 92.270 184.805 ;
        RECT 93.110 183.160 101.010 184.805 ;
        RECT 101.850 183.160 109.750 184.805 ;
        RECT 110.590 183.160 118.490 184.805 ;
        RECT 119.330 183.160 127.230 184.805 ;
        RECT 128.070 183.160 135.970 184.805 ;
        RECT 136.810 183.160 144.710 184.805 ;
        RECT 145.550 183.160 153.450 184.805 ;
        RECT 154.290 183.160 162.190 184.805 ;
        RECT 163.030 183.160 170.930 184.805 ;
        RECT 171.770 183.160 179.670 184.805 ;
        RECT 180.510 183.160 188.410 184.805 ;
        RECT 189.250 183.160 197.150 184.805 ;
        RECT 197.990 183.160 205.890 184.805 ;
        RECT 206.730 183.160 214.630 184.805 ;
        RECT 215.470 183.160 223.370 184.805 ;
        RECT 224.210 183.160 232.110 184.805 ;
        RECT 232.950 183.160 240.850 184.805 ;
        RECT 241.690 183.160 249.590 184.805 ;
        RECT 250.430 183.160 258.330 184.805 ;
        RECT 259.170 183.160 267.070 184.805 ;
        RECT 267.910 183.160 275.810 184.805 ;
        RECT 276.650 183.160 284.550 184.805 ;
        RECT 285.390 183.160 293.290 184.805 ;
        RECT 294.130 183.160 302.030 184.805 ;
        RECT 302.870 183.160 310.770 184.805 ;
        RECT 311.610 183.160 319.510 184.805 ;
        RECT 320.350 183.160 328.250 184.805 ;
        RECT 329.090 183.160 336.990 184.805 ;
        RECT 337.830 183.160 345.730 184.805 ;
        RECT 346.570 183.160 354.470 184.805 ;
        RECT 355.310 183.160 363.210 184.805 ;
        RECT 364.050 183.160 371.950 184.805 ;
        RECT 372.790 183.160 380.690 184.805 ;
        RECT 381.530 183.160 389.430 184.805 ;
        RECT 390.270 183.160 398.170 184.805 ;
        RECT 399.010 183.160 406.910 184.805 ;
        RECT 407.750 183.160 415.650 184.805 ;
        RECT 416.490 183.160 424.390 184.805 ;
        RECT 425.230 183.160 433.130 184.805 ;
        RECT 433.970 183.160 441.870 184.805 ;
        RECT 442.710 183.160 450.610 184.805 ;
        RECT 451.450 183.160 459.350 184.805 ;
        RECT 460.190 183.160 468.090 184.805 ;
        RECT 468.930 183.160 476.830 184.805 ;
        RECT 477.670 183.160 485.570 184.805 ;
        RECT 486.410 183.160 494.310 184.805 ;
        RECT 495.150 183.160 503.050 184.805 ;
        RECT 503.890 183.160 511.790 184.805 ;
        RECT 512.630 183.160 520.530 184.805 ;
        RECT 521.370 183.160 529.270 184.805 ;
        RECT 530.110 183.160 538.010 184.805 ;
        RECT 538.850 183.160 546.750 184.805 ;
        RECT 547.590 183.160 555.490 184.805 ;
        RECT 556.330 183.160 564.230 184.805 ;
        RECT 565.070 183.160 572.970 184.805 ;
        RECT 573.810 183.160 581.710 184.805 ;
        RECT 582.550 183.160 590.450 184.805 ;
        RECT 591.290 183.160 599.190 184.805 ;
        RECT 600.030 183.160 607.930 184.805 ;
        RECT 608.770 183.160 616.670 184.805 ;
        RECT 617.510 183.160 625.410 184.805 ;
        RECT 626.250 183.160 634.150 184.805 ;
        RECT 634.990 183.160 642.890 184.805 ;
        RECT 643.730 183.160 651.630 184.805 ;
        RECT 652.470 183.160 660.370 184.805 ;
        RECT 661.210 183.160 669.110 184.805 ;
        RECT 669.950 183.160 677.850 184.805 ;
        RECT 678.690 183.160 686.590 184.805 ;
        RECT 687.430 183.160 695.330 184.805 ;
        RECT 696.170 183.160 704.070 184.805 ;
        RECT 704.910 183.160 712.810 184.805 ;
        RECT 713.650 183.160 721.550 184.805 ;
        RECT 722.390 183.160 730.290 184.805 ;
        RECT 731.130 183.160 739.030 184.805 ;
        RECT 739.870 183.160 747.770 184.805 ;
        RECT 748.610 183.160 756.510 184.805 ;
        RECT 757.350 183.160 765.250 184.805 ;
        RECT 766.090 183.160 773.990 184.805 ;
        RECT 774.830 183.160 782.730 184.805 ;
        RECT 783.570 183.160 791.470 184.805 ;
        RECT 792.310 183.160 800.210 184.805 ;
        RECT 801.050 183.160 808.950 184.805 ;
        RECT 809.790 183.160 817.690 184.805 ;
        RECT 818.530 183.160 826.430 184.805 ;
        RECT 827.270 183.160 835.170 184.805 ;
        RECT 836.010 183.160 843.910 184.805 ;
        RECT 844.750 183.160 852.650 184.805 ;
        RECT 853.490 183.160 861.390 184.805 ;
        RECT 862.230 183.160 870.130 184.805 ;
        RECT 870.970 183.160 878.870 184.805 ;
        RECT 879.710 183.160 887.610 184.805 ;
        RECT 888.450 183.160 896.350 184.805 ;
        RECT 897.190 183.160 905.090 184.805 ;
        RECT 905.930 183.160 913.830 184.805 ;
        RECT 914.670 183.160 922.570 184.805 ;
        RECT 923.410 183.160 931.310 184.805 ;
        RECT 932.150 183.160 940.050 184.805 ;
        RECT 940.890 183.160 948.790 184.805 ;
        RECT 949.630 183.160 957.530 184.805 ;
        RECT 958.370 183.160 966.270 184.805 ;
        RECT 967.110 183.160 975.010 184.805 ;
        RECT 975.850 183.160 983.750 184.805 ;
        RECT 984.590 183.160 992.490 184.805 ;
        RECT 993.330 183.160 1001.230 184.805 ;
        RECT 1002.070 183.160 1009.970 184.805 ;
        RECT 1010.810 183.160 1018.710 184.805 ;
        RECT 1019.550 183.160 1027.450 184.805 ;
        RECT 1028.290 183.160 1036.190 184.805 ;
        RECT 1037.030 183.160 1044.930 184.805 ;
        RECT 1045.770 183.160 1053.670 184.805 ;
        RECT 1054.510 183.160 1062.410 184.805 ;
        RECT 1063.250 183.160 1071.150 184.805 ;
        RECT 1071.990 183.160 1079.890 184.805 ;
        RECT 1080.730 183.160 1088.630 184.805 ;
        RECT 1089.470 183.160 1097.370 184.805 ;
        RECT 1098.210 183.160 1106.110 184.805 ;
        RECT 1106.950 183.160 1114.850 184.805 ;
        RECT 1115.690 183.160 1123.590 184.805 ;
        RECT 1124.430 183.160 1132.330 184.805 ;
        RECT 1133.170 183.160 1141.070 184.805 ;
        RECT 1141.910 183.160 1169.680 184.805 ;
        RECT 1.470 2.280 1169.680 183.160 ;
        RECT 1.470 0.010 20.970 2.280 ;
        RECT 21.810 0.010 38.910 2.280 ;
        RECT 39.750 0.010 56.850 2.280 ;
        RECT 57.690 0.010 74.790 2.280 ;
        RECT 75.630 0.010 92.730 2.280 ;
        RECT 93.570 0.010 110.670 2.280 ;
        RECT 111.510 0.010 128.610 2.280 ;
        RECT 129.450 0.010 146.550 2.280 ;
        RECT 147.390 0.010 164.490 2.280 ;
        RECT 165.330 0.010 182.430 2.280 ;
        RECT 183.270 0.010 200.370 2.280 ;
        RECT 201.210 0.010 218.310 2.280 ;
        RECT 219.150 0.010 236.250 2.280 ;
        RECT 237.090 0.010 254.190 2.280 ;
        RECT 255.030 0.010 272.130 2.280 ;
        RECT 272.970 0.010 290.070 2.280 ;
        RECT 290.910 0.010 308.010 2.280 ;
        RECT 308.850 0.010 325.950 2.280 ;
        RECT 326.790 0.010 343.890 2.280 ;
        RECT 344.730 0.010 361.830 2.280 ;
        RECT 362.670 0.010 379.770 2.280 ;
        RECT 380.610 0.010 397.710 2.280 ;
        RECT 398.550 0.010 415.650 2.280 ;
        RECT 416.490 0.010 433.590 2.280 ;
        RECT 434.430 0.010 451.530 2.280 ;
        RECT 452.370 0.010 469.470 2.280 ;
        RECT 470.310 0.010 487.410 2.280 ;
        RECT 488.250 0.010 505.350 2.280 ;
        RECT 506.190 0.010 523.290 2.280 ;
        RECT 524.130 0.010 541.230 2.280 ;
        RECT 542.070 0.010 559.170 2.280 ;
        RECT 560.010 0.010 577.110 2.280 ;
        RECT 577.950 0.010 595.050 2.280 ;
        RECT 595.890 0.010 612.990 2.280 ;
        RECT 613.830 0.010 630.930 2.280 ;
        RECT 631.770 0.010 648.870 2.280 ;
        RECT 649.710 0.010 666.810 2.280 ;
        RECT 667.650 0.010 684.750 2.280 ;
        RECT 685.590 0.010 702.690 2.280 ;
        RECT 703.530 0.010 720.630 2.280 ;
        RECT 721.470 0.010 738.570 2.280 ;
        RECT 739.410 0.010 756.510 2.280 ;
        RECT 757.350 0.010 774.450 2.280 ;
        RECT 775.290 0.010 792.390 2.280 ;
        RECT 793.230 0.010 810.330 2.280 ;
        RECT 811.170 0.010 828.270 2.280 ;
        RECT 829.110 0.010 846.210 2.280 ;
        RECT 847.050 0.010 864.150 2.280 ;
        RECT 864.990 0.010 882.090 2.280 ;
        RECT 882.930 0.010 900.030 2.280 ;
        RECT 900.870 0.010 917.970 2.280 ;
        RECT 918.810 0.010 935.910 2.280 ;
        RECT 936.750 0.010 953.850 2.280 ;
        RECT 954.690 0.010 971.790 2.280 ;
        RECT 972.630 0.010 989.730 2.280 ;
        RECT 990.570 0.010 1007.670 2.280 ;
        RECT 1008.510 0.010 1025.610 2.280 ;
        RECT 1026.450 0.010 1043.550 2.280 ;
        RECT 1044.390 0.010 1061.490 2.280 ;
        RECT 1062.330 0.010 1079.430 2.280 ;
        RECT 1080.270 0.010 1097.370 2.280 ;
        RECT 1098.210 0.010 1115.310 2.280 ;
        RECT 1116.150 0.010 1133.250 2.280 ;
        RECT 1134.090 0.010 1151.190 2.280 ;
        RECT 1152.030 0.010 1169.680 2.280 ;
      LAYER met3 ;
        RECT 1.445 177.160 1171.460 184.785 ;
        RECT 1.445 175.760 1171.060 177.160 ;
        RECT 1.445 173.080 1171.460 175.760 ;
        RECT 2.400 171.680 1171.460 173.080 ;
        RECT 1.445 164.240 1171.460 171.680 ;
        RECT 1.445 162.840 1171.060 164.240 ;
        RECT 1.445 151.320 1171.460 162.840 ;
        RECT 1.445 149.920 1171.060 151.320 ;
        RECT 1.445 146.560 1171.460 149.920 ;
        RECT 2.400 145.160 1171.460 146.560 ;
        RECT 1.445 138.400 1171.460 145.160 ;
        RECT 1.445 137.000 1171.060 138.400 ;
        RECT 1.445 125.480 1171.460 137.000 ;
        RECT 1.445 124.080 1171.060 125.480 ;
        RECT 1.445 120.040 1171.460 124.080 ;
        RECT 2.400 118.640 1171.460 120.040 ;
        RECT 1.445 112.560 1171.460 118.640 ;
        RECT 1.445 111.160 1171.060 112.560 ;
        RECT 1.445 99.640 1171.460 111.160 ;
        RECT 1.445 98.240 1171.060 99.640 ;
        RECT 1.445 93.520 1171.460 98.240 ;
        RECT 2.400 92.120 1171.460 93.520 ;
        RECT 1.445 86.720 1171.460 92.120 ;
        RECT 1.445 85.320 1171.060 86.720 ;
        RECT 1.445 73.800 1171.460 85.320 ;
        RECT 1.445 72.400 1171.060 73.800 ;
        RECT 1.445 67.000 1171.460 72.400 ;
        RECT 2.400 65.600 1171.460 67.000 ;
        RECT 1.445 60.880 1171.460 65.600 ;
        RECT 1.445 59.480 1171.060 60.880 ;
        RECT 1.445 47.960 1171.460 59.480 ;
        RECT 1.445 46.560 1171.060 47.960 ;
        RECT 1.445 40.480 1171.460 46.560 ;
        RECT 2.400 39.080 1171.460 40.480 ;
        RECT 1.445 35.040 1171.460 39.080 ;
        RECT 1.445 33.640 1171.060 35.040 ;
        RECT 1.445 22.120 1171.460 33.640 ;
        RECT 1.445 20.720 1171.060 22.120 ;
        RECT 1.445 13.960 1171.460 20.720 ;
        RECT 2.400 12.560 1171.460 13.960 ;
        RECT 1.445 9.200 1171.460 12.560 ;
        RECT 1.445 7.800 1171.060 9.200 ;
        RECT 1.445 0.175 1171.460 7.800 ;
      LAYER met4 ;
        RECT 4.895 182.880 1060.465 184.785 ;
        RECT 4.895 2.215 5.810 182.880 ;
        RECT 9.710 2.215 95.810 182.880 ;
        RECT 99.710 2.215 185.810 182.880 ;
        RECT 189.710 2.215 275.810 182.880 ;
        RECT 279.710 2.215 365.810 182.880 ;
        RECT 369.710 2.215 455.810 182.880 ;
        RECT 459.710 2.215 545.810 182.880 ;
        RECT 549.710 2.215 635.810 182.880 ;
        RECT 639.710 2.215 725.810 182.880 ;
        RECT 729.710 2.215 815.810 182.880 ;
        RECT 819.710 2.215 905.810 182.880 ;
        RECT 909.710 2.215 995.810 182.880 ;
        RECT 999.710 2.215 1060.465 182.880 ;
  END
END RAM32_1RW1R
END LIBRARY

