VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM512
  CLASS BLOCK ;
  FOREIGN RAM512 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1587.460 BY 987.360 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 520.240 1587.460 520.840 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 574.640 1587.460 575.240 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 629.040 1587.460 629.640 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 683.440 1587.460 684.040 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 737.840 1587.460 738.440 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 792.240 1587.460 792.840 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 846.640 1587.460 847.240 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 901.040 1587.460 901.640 ;
    END
  END A0[7]
  PIN A0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 955.440 1587.460 956.040 ;
    END
  END A0[8]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 2.000 493.640 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 0.000 464.510 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 0.000 513.270 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 0.000 635.170 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.270 0.000 659.550 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.650 0.000 683.930 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 0.000 708.310 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 0.000 732.690 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 2.000 ;
    END
  END Di0[31]
  PIN Di0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 0.000 805.830 2.000 ;
    END
  END Di0[32]
  PIN Di0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.930 0.000 830.210 2.000 ;
    END
  END Di0[33]
  PIN Di0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.310 0.000 854.590 2.000 ;
    END
  END Di0[34]
  PIN Di0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 0.000 878.970 2.000 ;
    END
  END Di0[35]
  PIN Di0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.070 0.000 903.350 2.000 ;
    END
  END Di0[36]
  PIN Di0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 2.000 ;
    END
  END Di0[37]
  PIN Di0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.830 0.000 952.110 2.000 ;
    END
  END Di0[38]
  PIN Di0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.210 0.000 976.490 2.000 ;
    END
  END Di0[39]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 2.000 ;
    END
  END Di0[3]
  PIN Di0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.590 0.000 1000.870 2.000 ;
    END
  END Di0[40]
  PIN Di0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.970 0.000 1025.250 2.000 ;
    END
  END Di0[41]
  PIN Di0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.350 0.000 1049.630 2.000 ;
    END
  END Di0[42]
  PIN Di0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.730 0.000 1074.010 2.000 ;
    END
  END Di0[43]
  PIN Di0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 2.000 ;
    END
  END Di0[44]
  PIN Di0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.490 0.000 1122.770 2.000 ;
    END
  END Di0[45]
  PIN Di0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.870 0.000 1147.150 2.000 ;
    END
  END Di0[46]
  PIN Di0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.250 0.000 1171.530 2.000 ;
    END
  END Di0[47]
  PIN Di0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.630 0.000 1195.910 2.000 ;
    END
  END Di0[48]
  PIN Di0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.010 0.000 1220.290 2.000 ;
    END
  END Di0[49]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 2.000 ;
    END
  END Di0[4]
  PIN Di0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.390 0.000 1244.670 2.000 ;
    END
  END Di0[50]
  PIN Di0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 0.000 1269.050 2.000 ;
    END
  END Di0[51]
  PIN Di0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.150 0.000 1293.430 2.000 ;
    END
  END Di0[52]
  PIN Di0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.530 0.000 1317.810 2.000 ;
    END
  END Di0[53]
  PIN Di0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.910 0.000 1342.190 2.000 ;
    END
  END Di0[54]
  PIN Di0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.290 0.000 1366.570 2.000 ;
    END
  END Di0[55]
  PIN Di0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.670 0.000 1390.950 2.000 ;
    END
  END Di0[56]
  PIN Di0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.050 0.000 1415.330 2.000 ;
    END
  END Di0[57]
  PIN Di0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 0.000 1439.710 2.000 ;
    END
  END Di0[58]
  PIN Di0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1463.810 0.000 1464.090 2.000 ;
    END
  END Di0[59]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 2.000 ;
    END
  END Di0[5]
  PIN Di0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1488.190 0.000 1488.470 2.000 ;
    END
  END Di0[60]
  PIN Di0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.570 0.000 1512.850 2.000 ;
    END
  END Di0[61]
  PIN Di0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.950 0.000 1537.230 2.000 ;
    END
  END Di0[62]
  PIN Di0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.330 0.000 1561.610 2.000 ;
    END
  END Di0[63]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 985.360 25.670 987.360 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 985.360 269.470 987.360 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 985.360 293.850 987.360 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 985.360 318.230 987.360 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 985.360 342.610 987.360 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 985.360 366.990 987.360 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 985.360 391.370 987.360 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 985.360 415.750 987.360 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 985.360 440.130 987.360 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 985.360 464.510 987.360 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 985.360 488.890 987.360 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 985.360 50.050 987.360 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 985.360 513.270 987.360 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 985.360 537.650 987.360 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 985.360 562.030 987.360 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 985.360 586.410 987.360 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 985.360 610.790 987.360 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 985.360 635.170 987.360 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.270 985.360 659.550 987.360 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.650 985.360 683.930 987.360 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 985.360 708.310 987.360 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 985.360 732.690 987.360 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 985.360 74.430 987.360 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 985.360 757.070 987.360 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 985.360 781.450 987.360 ;
    END
  END Do0[31]
  PIN Do0[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 985.360 805.830 987.360 ;
    END
  END Do0[32]
  PIN Do0[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.930 985.360 830.210 987.360 ;
    END
  END Do0[33]
  PIN Do0[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.310 985.360 854.590 987.360 ;
    END
  END Do0[34]
  PIN Do0[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 985.360 878.970 987.360 ;
    END
  END Do0[35]
  PIN Do0[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.070 985.360 903.350 987.360 ;
    END
  END Do0[36]
  PIN Do0[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 985.360 927.730 987.360 ;
    END
  END Do0[37]
  PIN Do0[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.830 985.360 952.110 987.360 ;
    END
  END Do0[38]
  PIN Do0[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.210 985.360 976.490 987.360 ;
    END
  END Do0[39]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 985.360 98.810 987.360 ;
    END
  END Do0[3]
  PIN Do0[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.590 985.360 1000.870 987.360 ;
    END
  END Do0[40]
  PIN Do0[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.970 985.360 1025.250 987.360 ;
    END
  END Do0[41]
  PIN Do0[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.350 985.360 1049.630 987.360 ;
    END
  END Do0[42]
  PIN Do0[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.730 985.360 1074.010 987.360 ;
    END
  END Do0[43]
  PIN Do0[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 985.360 1098.390 987.360 ;
    END
  END Do0[44]
  PIN Do0[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.490 985.360 1122.770 987.360 ;
    END
  END Do0[45]
  PIN Do0[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.870 985.360 1147.150 987.360 ;
    END
  END Do0[46]
  PIN Do0[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.250 985.360 1171.530 987.360 ;
    END
  END Do0[47]
  PIN Do0[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.630 985.360 1195.910 987.360 ;
    END
  END Do0[48]
  PIN Do0[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.010 985.360 1220.290 987.360 ;
    END
  END Do0[49]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 985.360 123.190 987.360 ;
    END
  END Do0[4]
  PIN Do0[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.390 985.360 1244.670 987.360 ;
    END
  END Do0[50]
  PIN Do0[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 985.360 1269.050 987.360 ;
    END
  END Do0[51]
  PIN Do0[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.150 985.360 1293.430 987.360 ;
    END
  END Do0[52]
  PIN Do0[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.530 985.360 1317.810 987.360 ;
    END
  END Do0[53]
  PIN Do0[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.910 985.360 1342.190 987.360 ;
    END
  END Do0[54]
  PIN Do0[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.290 985.360 1366.570 987.360 ;
    END
  END Do0[55]
  PIN Do0[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.670 985.360 1390.950 987.360 ;
    END
  END Do0[56]
  PIN Do0[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.050 985.360 1415.330 987.360 ;
    END
  END Do0[57]
  PIN Do0[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 985.360 1439.710 987.360 ;
    END
  END Do0[58]
  PIN Do0[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1463.810 985.360 1464.090 987.360 ;
    END
  END Do0[59]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 985.360 147.570 987.360 ;
    END
  END Do0[5]
  PIN Do0[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1488.190 985.360 1488.470 987.360 ;
    END
  END Do0[60]
  PIN Do0[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.570 985.360 1512.850 987.360 ;
    END
  END Do0[61]
  PIN Do0[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.950 985.360 1537.230 987.360 ;
    END
  END Do0[62]
  PIN Do0[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.330 985.360 1561.610 987.360 ;
    END
  END Do0[63]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 985.360 171.950 987.360 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 985.360 196.330 987.360 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 985.360 220.710 987.360 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 985.360 245.090 987.360 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 30.640 1587.460 31.240 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 113.690 100.400 116.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 293.690 100.400 296.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 473.690 100.400 476.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 653.690 100.400 656.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 833.690 100.400 836.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.690 100.400 1016.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1193.690 100.400 1196.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.690 100.400 1376.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1553.690 100.400 1556.790 886.960 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.690 100.400 26.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.690 100.400 206.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.690 100.400 386.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.690 100.400 566.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.690 100.400 746.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.690 100.400 926.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.690 100.400 1106.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1283.690 100.400 1286.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.690 100.400 1466.790 886.960 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 85.040 1587.460 85.640 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 139.440 1587.460 140.040 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 193.840 1587.460 194.440 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 248.240 1587.460 248.840 ;
    END
  END WE0[3]
  PIN WE0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 302.640 1587.460 303.240 ;
    END
  END WE0[4]
  PIN WE0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 357.040 1587.460 357.640 ;
    END
  END WE0[5]
  PIN WE0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 411.440 1587.460 412.040 ;
    END
  END WE0[6]
  PIN WE0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1585.460 465.840 1587.460 466.440 ;
    END
  END WE0[7]
  OBS
      LAYER li1 ;
        RECT 20.240 100.555 1567.220 886.805 ;
      LAYER met1 ;
        RECT 3.290 0.380 1574.510 987.320 ;
      LAYER met2 ;
        RECT 3.320 985.080 25.110 987.350 ;
        RECT 25.950 985.080 49.490 987.350 ;
        RECT 50.330 985.080 73.870 987.350 ;
        RECT 74.710 985.080 98.250 987.350 ;
        RECT 99.090 985.080 122.630 987.350 ;
        RECT 123.470 985.080 147.010 987.350 ;
        RECT 147.850 985.080 171.390 987.350 ;
        RECT 172.230 985.080 195.770 987.350 ;
        RECT 196.610 985.080 220.150 987.350 ;
        RECT 220.990 985.080 244.530 987.350 ;
        RECT 245.370 985.080 268.910 987.350 ;
        RECT 269.750 985.080 293.290 987.350 ;
        RECT 294.130 985.080 317.670 987.350 ;
        RECT 318.510 985.080 342.050 987.350 ;
        RECT 342.890 985.080 366.430 987.350 ;
        RECT 367.270 985.080 390.810 987.350 ;
        RECT 391.650 985.080 415.190 987.350 ;
        RECT 416.030 985.080 439.570 987.350 ;
        RECT 440.410 985.080 463.950 987.350 ;
        RECT 464.790 985.080 488.330 987.350 ;
        RECT 489.170 985.080 512.710 987.350 ;
        RECT 513.550 985.080 537.090 987.350 ;
        RECT 537.930 985.080 561.470 987.350 ;
        RECT 562.310 985.080 585.850 987.350 ;
        RECT 586.690 985.080 610.230 987.350 ;
        RECT 611.070 985.080 634.610 987.350 ;
        RECT 635.450 985.080 658.990 987.350 ;
        RECT 659.830 985.080 683.370 987.350 ;
        RECT 684.210 985.080 707.750 987.350 ;
        RECT 708.590 985.080 732.130 987.350 ;
        RECT 732.970 985.080 756.510 987.350 ;
        RECT 757.350 985.080 780.890 987.350 ;
        RECT 781.730 985.080 805.270 987.350 ;
        RECT 806.110 985.080 829.650 987.350 ;
        RECT 830.490 985.080 854.030 987.350 ;
        RECT 854.870 985.080 878.410 987.350 ;
        RECT 879.250 985.080 902.790 987.350 ;
        RECT 903.630 985.080 927.170 987.350 ;
        RECT 928.010 985.080 951.550 987.350 ;
        RECT 952.390 985.080 975.930 987.350 ;
        RECT 976.770 985.080 1000.310 987.350 ;
        RECT 1001.150 985.080 1024.690 987.350 ;
        RECT 1025.530 985.080 1049.070 987.350 ;
        RECT 1049.910 985.080 1073.450 987.350 ;
        RECT 1074.290 985.080 1097.830 987.350 ;
        RECT 1098.670 985.080 1122.210 987.350 ;
        RECT 1123.050 985.080 1146.590 987.350 ;
        RECT 1147.430 985.080 1170.970 987.350 ;
        RECT 1171.810 985.080 1195.350 987.350 ;
        RECT 1196.190 985.080 1219.730 987.350 ;
        RECT 1220.570 985.080 1244.110 987.350 ;
        RECT 1244.950 985.080 1268.490 987.350 ;
        RECT 1269.330 985.080 1292.870 987.350 ;
        RECT 1293.710 985.080 1317.250 987.350 ;
        RECT 1318.090 985.080 1341.630 987.350 ;
        RECT 1342.470 985.080 1366.010 987.350 ;
        RECT 1366.850 985.080 1390.390 987.350 ;
        RECT 1391.230 985.080 1414.770 987.350 ;
        RECT 1415.610 985.080 1439.150 987.350 ;
        RECT 1439.990 985.080 1463.530 987.350 ;
        RECT 1464.370 985.080 1487.910 987.350 ;
        RECT 1488.750 985.080 1512.290 987.350 ;
        RECT 1513.130 985.080 1536.670 987.350 ;
        RECT 1537.510 985.080 1561.050 987.350 ;
        RECT 1561.890 985.080 1574.480 987.350 ;
        RECT 3.320 2.280 1574.480 985.080 ;
        RECT 3.320 0.350 25.110 2.280 ;
        RECT 25.950 0.350 49.490 2.280 ;
        RECT 50.330 0.350 73.870 2.280 ;
        RECT 74.710 0.350 98.250 2.280 ;
        RECT 99.090 0.350 122.630 2.280 ;
        RECT 123.470 0.350 147.010 2.280 ;
        RECT 147.850 0.350 171.390 2.280 ;
        RECT 172.230 0.350 195.770 2.280 ;
        RECT 196.610 0.350 220.150 2.280 ;
        RECT 220.990 0.350 244.530 2.280 ;
        RECT 245.370 0.350 268.910 2.280 ;
        RECT 269.750 0.350 293.290 2.280 ;
        RECT 294.130 0.350 317.670 2.280 ;
        RECT 318.510 0.350 342.050 2.280 ;
        RECT 342.890 0.350 366.430 2.280 ;
        RECT 367.270 0.350 390.810 2.280 ;
        RECT 391.650 0.350 415.190 2.280 ;
        RECT 416.030 0.350 439.570 2.280 ;
        RECT 440.410 0.350 463.950 2.280 ;
        RECT 464.790 0.350 488.330 2.280 ;
        RECT 489.170 0.350 512.710 2.280 ;
        RECT 513.550 0.350 537.090 2.280 ;
        RECT 537.930 0.350 561.470 2.280 ;
        RECT 562.310 0.350 585.850 2.280 ;
        RECT 586.690 0.350 610.230 2.280 ;
        RECT 611.070 0.350 634.610 2.280 ;
        RECT 635.450 0.350 658.990 2.280 ;
        RECT 659.830 0.350 683.370 2.280 ;
        RECT 684.210 0.350 707.750 2.280 ;
        RECT 708.590 0.350 732.130 2.280 ;
        RECT 732.970 0.350 756.510 2.280 ;
        RECT 757.350 0.350 780.890 2.280 ;
        RECT 781.730 0.350 805.270 2.280 ;
        RECT 806.110 0.350 829.650 2.280 ;
        RECT 830.490 0.350 854.030 2.280 ;
        RECT 854.870 0.350 878.410 2.280 ;
        RECT 879.250 0.350 902.790 2.280 ;
        RECT 903.630 0.350 927.170 2.280 ;
        RECT 928.010 0.350 951.550 2.280 ;
        RECT 952.390 0.350 975.930 2.280 ;
        RECT 976.770 0.350 1000.310 2.280 ;
        RECT 1001.150 0.350 1024.690 2.280 ;
        RECT 1025.530 0.350 1049.070 2.280 ;
        RECT 1049.910 0.350 1073.450 2.280 ;
        RECT 1074.290 0.350 1097.830 2.280 ;
        RECT 1098.670 0.350 1122.210 2.280 ;
        RECT 1123.050 0.350 1146.590 2.280 ;
        RECT 1147.430 0.350 1170.970 2.280 ;
        RECT 1171.810 0.350 1195.350 2.280 ;
        RECT 1196.190 0.350 1219.730 2.280 ;
        RECT 1220.570 0.350 1244.110 2.280 ;
        RECT 1244.950 0.350 1268.490 2.280 ;
        RECT 1269.330 0.350 1292.870 2.280 ;
        RECT 1293.710 0.350 1317.250 2.280 ;
        RECT 1318.090 0.350 1341.630 2.280 ;
        RECT 1342.470 0.350 1366.010 2.280 ;
        RECT 1366.850 0.350 1390.390 2.280 ;
        RECT 1391.230 0.350 1414.770 2.280 ;
        RECT 1415.610 0.350 1439.150 2.280 ;
        RECT 1439.990 0.350 1463.530 2.280 ;
        RECT 1464.370 0.350 1487.910 2.280 ;
        RECT 1488.750 0.350 1512.290 2.280 ;
        RECT 1513.130 0.350 1536.670 2.280 ;
        RECT 1537.510 0.350 1561.050 2.280 ;
        RECT 1561.890 0.350 1574.480 2.280 ;
      LAYER met3 ;
        RECT 2.000 956.440 1585.460 987.185 ;
        RECT 2.000 955.040 1585.060 956.440 ;
        RECT 2.000 902.040 1585.460 955.040 ;
        RECT 2.000 900.640 1585.060 902.040 ;
        RECT 2.000 847.640 1585.460 900.640 ;
        RECT 2.000 846.240 1585.060 847.640 ;
        RECT 2.000 793.240 1585.460 846.240 ;
        RECT 2.000 791.840 1585.060 793.240 ;
        RECT 2.000 738.840 1585.460 791.840 ;
        RECT 2.000 737.440 1585.060 738.840 ;
        RECT 2.000 684.440 1585.460 737.440 ;
        RECT 2.000 683.040 1585.060 684.440 ;
        RECT 2.000 630.040 1585.460 683.040 ;
        RECT 2.000 628.640 1585.060 630.040 ;
        RECT 2.000 575.640 1585.460 628.640 ;
        RECT 2.000 574.240 1585.060 575.640 ;
        RECT 2.000 521.240 1585.460 574.240 ;
        RECT 2.000 519.840 1585.060 521.240 ;
        RECT 2.000 494.040 1585.460 519.840 ;
        RECT 2.400 492.640 1585.460 494.040 ;
        RECT 2.000 466.840 1585.460 492.640 ;
        RECT 2.000 465.440 1585.060 466.840 ;
        RECT 2.000 412.440 1585.460 465.440 ;
        RECT 2.000 411.040 1585.060 412.440 ;
        RECT 2.000 358.040 1585.460 411.040 ;
        RECT 2.000 356.640 1585.060 358.040 ;
        RECT 2.000 303.640 1585.460 356.640 ;
        RECT 2.000 302.240 1585.060 303.640 ;
        RECT 2.000 249.240 1585.460 302.240 ;
        RECT 2.000 247.840 1585.060 249.240 ;
        RECT 2.000 194.840 1585.460 247.840 ;
        RECT 2.000 193.440 1585.060 194.840 ;
        RECT 2.000 140.440 1585.460 193.440 ;
        RECT 2.000 139.040 1585.060 140.440 ;
        RECT 2.000 86.040 1585.460 139.040 ;
        RECT 2.000 84.640 1585.060 86.040 ;
        RECT 2.000 31.640 1585.460 84.640 ;
        RECT 2.000 30.240 1585.060 31.640 ;
        RECT 2.000 0.855 1585.460 30.240 ;
      LAYER met4 ;
        RECT 42.615 887.360 1570.145 987.185 ;
        RECT 42.615 100.000 113.290 887.360 ;
        RECT 117.190 100.000 203.290 887.360 ;
        RECT 207.190 100.000 293.290 887.360 ;
        RECT 297.190 100.000 383.290 887.360 ;
        RECT 387.190 100.000 473.290 887.360 ;
        RECT 477.190 100.000 563.290 887.360 ;
        RECT 567.190 100.000 653.290 887.360 ;
        RECT 657.190 100.000 743.290 887.360 ;
        RECT 747.190 100.000 833.290 887.360 ;
        RECT 837.190 100.000 923.290 887.360 ;
        RECT 927.190 100.000 1013.290 887.360 ;
        RECT 1017.190 100.000 1103.290 887.360 ;
        RECT 1107.190 100.000 1193.290 887.360 ;
        RECT 1197.190 100.000 1283.290 887.360 ;
        RECT 1287.190 100.000 1373.290 887.360 ;
        RECT 1377.190 100.000 1463.290 887.360 ;
        RECT 1467.190 100.000 1553.290 887.360 ;
        RECT 1557.190 100.000 1570.145 887.360 ;
        RECT 42.615 0.855 1570.145 100.000 ;
  END
END RAM512
END LIBRARY

