magic
tech sky130A
magscale 1 2
timestamp 1662543620
<< obsli1 >>
rect 4048 20111 312708 177361
<< obsm1 >>
rect 658 76 315086 197464
<< metal2 >>
rect 4710 197072 4766 197472
rect 9586 197072 9642 197472
rect 14462 197072 14518 197472
rect 19338 197072 19394 197472
rect 24214 197072 24270 197472
rect 29090 197072 29146 197472
rect 33966 197072 34022 197472
rect 38842 197072 38898 197472
rect 43718 197072 43774 197472
rect 48594 197072 48650 197472
rect 53470 197072 53526 197472
rect 58346 197072 58402 197472
rect 63222 197072 63278 197472
rect 68098 197072 68154 197472
rect 72974 197072 73030 197472
rect 77850 197072 77906 197472
rect 82726 197072 82782 197472
rect 87602 197072 87658 197472
rect 92478 197072 92534 197472
rect 97354 197072 97410 197472
rect 102230 197072 102286 197472
rect 107106 197072 107162 197472
rect 111982 197072 112038 197472
rect 116858 197072 116914 197472
rect 121734 197072 121790 197472
rect 126610 197072 126666 197472
rect 131486 197072 131542 197472
rect 136362 197072 136418 197472
rect 141238 197072 141294 197472
rect 146114 197072 146170 197472
rect 150990 197072 151046 197472
rect 155866 197072 155922 197472
rect 160742 197072 160798 197472
rect 165618 197072 165674 197472
rect 170494 197072 170550 197472
rect 175370 197072 175426 197472
rect 180246 197072 180302 197472
rect 185122 197072 185178 197472
rect 189998 197072 190054 197472
rect 194874 197072 194930 197472
rect 199750 197072 199806 197472
rect 204626 197072 204682 197472
rect 209502 197072 209558 197472
rect 214378 197072 214434 197472
rect 219254 197072 219310 197472
rect 224130 197072 224186 197472
rect 229006 197072 229062 197472
rect 233882 197072 233938 197472
rect 238758 197072 238814 197472
rect 243634 197072 243690 197472
rect 248510 197072 248566 197472
rect 253386 197072 253442 197472
rect 258262 197072 258318 197472
rect 263138 197072 263194 197472
rect 268014 197072 268070 197472
rect 272890 197072 272946 197472
rect 277766 197072 277822 197472
rect 282642 197072 282698 197472
rect 287518 197072 287574 197472
rect 292394 197072 292450 197472
rect 297270 197072 297326 197472
rect 302146 197072 302202 197472
rect 307022 197072 307078 197472
rect 311898 197072 311954 197472
rect 4710 0 4766 400
rect 9586 0 9642 400
rect 14462 0 14518 400
rect 19338 0 19394 400
rect 24214 0 24270 400
rect 29090 0 29146 400
rect 33966 0 34022 400
rect 38842 0 38898 400
rect 43718 0 43774 400
rect 48594 0 48650 400
rect 53470 0 53526 400
rect 58346 0 58402 400
rect 63222 0 63278 400
rect 68098 0 68154 400
rect 72974 0 73030 400
rect 77850 0 77906 400
rect 82726 0 82782 400
rect 87602 0 87658 400
rect 92478 0 92534 400
rect 97354 0 97410 400
rect 102230 0 102286 400
rect 107106 0 107162 400
rect 111982 0 112038 400
rect 116858 0 116914 400
rect 121734 0 121790 400
rect 126610 0 126666 400
rect 131486 0 131542 400
rect 136362 0 136418 400
rect 141238 0 141294 400
rect 146114 0 146170 400
rect 150990 0 151046 400
rect 155866 0 155922 400
rect 160742 0 160798 400
rect 165618 0 165674 400
rect 170494 0 170550 400
rect 175370 0 175426 400
rect 180246 0 180302 400
rect 185122 0 185178 400
rect 189998 0 190054 400
rect 194874 0 194930 400
rect 199750 0 199806 400
rect 204626 0 204682 400
rect 209502 0 209558 400
rect 214378 0 214434 400
rect 219254 0 219310 400
rect 224130 0 224186 400
rect 229006 0 229062 400
rect 233882 0 233938 400
rect 238758 0 238814 400
rect 243634 0 243690 400
rect 248510 0 248566 400
rect 253386 0 253442 400
rect 258262 0 258318 400
rect 263138 0 263194 400
rect 268014 0 268070 400
rect 272890 0 272946 400
rect 277766 0 277822 400
rect 282642 0 282698 400
rect 287518 0 287574 400
rect 292394 0 292450 400
rect 297270 0 297326 400
rect 302146 0 302202 400
rect 307022 0 307078 400
rect 311898 0 311954 400
<< obsm2 >>
rect 664 197016 4654 197470
rect 4822 197016 9530 197470
rect 9698 197016 14406 197470
rect 14574 197016 19282 197470
rect 19450 197016 24158 197470
rect 24326 197016 29034 197470
rect 29202 197016 33910 197470
rect 34078 197016 38786 197470
rect 38954 197016 43662 197470
rect 43830 197016 48538 197470
rect 48706 197016 53414 197470
rect 53582 197016 58290 197470
rect 58458 197016 63166 197470
rect 63334 197016 68042 197470
rect 68210 197016 72918 197470
rect 73086 197016 77794 197470
rect 77962 197016 82670 197470
rect 82838 197016 87546 197470
rect 87714 197016 92422 197470
rect 92590 197016 97298 197470
rect 97466 197016 102174 197470
rect 102342 197016 107050 197470
rect 107218 197016 111926 197470
rect 112094 197016 116802 197470
rect 116970 197016 121678 197470
rect 121846 197016 126554 197470
rect 126722 197016 131430 197470
rect 131598 197016 136306 197470
rect 136474 197016 141182 197470
rect 141350 197016 146058 197470
rect 146226 197016 150934 197470
rect 151102 197016 155810 197470
rect 155978 197016 160686 197470
rect 160854 197016 165562 197470
rect 165730 197016 170438 197470
rect 170606 197016 175314 197470
rect 175482 197016 180190 197470
rect 180358 197016 185066 197470
rect 185234 197016 189942 197470
rect 190110 197016 194818 197470
rect 194986 197016 199694 197470
rect 199862 197016 204570 197470
rect 204738 197016 209446 197470
rect 209614 197016 214322 197470
rect 214490 197016 219198 197470
rect 219366 197016 224074 197470
rect 224242 197016 228950 197470
rect 229118 197016 233826 197470
rect 233994 197016 238702 197470
rect 238870 197016 243578 197470
rect 243746 197016 248454 197470
rect 248622 197016 253330 197470
rect 253498 197016 258206 197470
rect 258374 197016 263082 197470
rect 263250 197016 267958 197470
rect 268126 197016 272834 197470
rect 273002 197016 277710 197470
rect 277878 197016 282586 197470
rect 282754 197016 287462 197470
rect 287630 197016 292338 197470
rect 292506 197016 297214 197470
rect 297382 197016 302090 197470
rect 302258 197016 306966 197470
rect 307134 197016 311842 197470
rect 312010 197016 315082 197470
rect 664 456 315082 197016
rect 664 70 4654 456
rect 4822 70 9530 456
rect 9698 70 14406 456
rect 14574 70 19282 456
rect 19450 70 24158 456
rect 24326 70 29034 456
rect 29202 70 33910 456
rect 34078 70 38786 456
rect 38954 70 43662 456
rect 43830 70 48538 456
rect 48706 70 53414 456
rect 53582 70 58290 456
rect 58458 70 63166 456
rect 63334 70 68042 456
rect 68210 70 72918 456
rect 73086 70 77794 456
rect 77962 70 82670 456
rect 82838 70 87546 456
rect 87714 70 92422 456
rect 92590 70 97298 456
rect 97466 70 102174 456
rect 102342 70 107050 456
rect 107218 70 111926 456
rect 112094 70 116802 456
rect 116970 70 121678 456
rect 121846 70 126554 456
rect 126722 70 131430 456
rect 131598 70 136306 456
rect 136474 70 141182 456
rect 141350 70 146058 456
rect 146226 70 150934 456
rect 151102 70 155810 456
rect 155978 70 160686 456
rect 160854 70 165562 456
rect 165730 70 170438 456
rect 170606 70 175314 456
rect 175482 70 180190 456
rect 180358 70 185066 456
rect 185234 70 189942 456
rect 190110 70 194818 456
rect 194986 70 199694 456
rect 199862 70 204570 456
rect 204738 70 209446 456
rect 209614 70 214322 456
rect 214490 70 219198 456
rect 219366 70 224074 456
rect 224242 70 228950 456
rect 229118 70 233826 456
rect 233994 70 238702 456
rect 238870 70 243578 456
rect 243746 70 248454 456
rect 248622 70 253330 456
rect 253498 70 258206 456
rect 258374 70 263082 456
rect 263250 70 267958 456
rect 268126 70 272834 456
rect 273002 70 277710 456
rect 277878 70 282586 456
rect 282754 70 287462 456
rect 287630 70 292338 456
rect 292506 70 297214 456
rect 297382 70 302090 456
rect 302258 70 306966 456
rect 307134 70 311842 456
rect 312010 70 315082 456
<< metal3 >>
rect 316356 191088 316756 191208
rect 316356 180208 316756 180328
rect 316356 169328 316756 169448
rect 316356 158448 316756 158568
rect 316356 147568 316756 147688
rect 316356 136688 316756 136808
rect 316356 125808 316756 125928
rect 316356 114928 316756 115048
rect 316356 104048 316756 104168
rect 0 98608 400 98728
rect 316356 93168 316756 93288
rect 316356 82288 316756 82408
rect 316356 71408 316756 71528
rect 316356 60528 316756 60648
rect 316356 49648 316756 49768
rect 316356 38768 316756 38888
rect 316356 27888 316756 28008
rect 316356 17008 316756 17128
rect 316356 6128 316756 6248
<< obsm3 >>
rect 400 191288 316356 197437
rect 400 191008 316276 191288
rect 400 180408 316356 191008
rect 400 180128 316276 180408
rect 400 169528 316356 180128
rect 400 169248 316276 169528
rect 400 158648 316356 169248
rect 400 158368 316276 158648
rect 400 147768 316356 158368
rect 400 147488 316276 147768
rect 400 136888 316356 147488
rect 400 136608 316276 136888
rect 400 126008 316356 136608
rect 400 125728 316276 126008
rect 400 115128 316356 125728
rect 400 114848 316276 115128
rect 400 104248 316356 114848
rect 400 103968 316276 104248
rect 400 98808 316356 103968
rect 480 98528 316356 98808
rect 400 93368 316356 98528
rect 400 93088 316276 93368
rect 400 82488 316356 93088
rect 400 82208 316276 82488
rect 400 71608 316356 82208
rect 400 71328 316276 71608
rect 400 60728 316356 71328
rect 400 60448 316276 60728
rect 400 49848 316356 60448
rect 400 49568 316276 49848
rect 400 38968 316356 49568
rect 400 38688 316276 38968
rect 400 28088 316356 38688
rect 400 27808 316276 28088
rect 400 17208 316356 27808
rect 400 16928 316276 17208
rect 400 6328 316356 16928
rect 400 6048 316276 6328
rect 400 171 316356 6048
<< metal4 >>
rect 4738 20080 5358 177392
rect 22738 20080 23358 177392
rect 40738 20080 41358 177392
rect 58738 20080 59358 177392
rect 76738 20080 77358 177392
rect 94738 20080 95358 177392
rect 112738 20080 113358 177392
rect 130738 20080 131358 177392
rect 148738 20080 149358 177392
rect 166738 20080 167358 177392
rect 184738 20080 185358 177392
rect 202738 20080 203358 177392
rect 220738 20080 221358 177392
rect 238738 20080 239358 177392
rect 256738 20080 257358 177392
rect 274738 20080 275358 177392
rect 292738 20080 293358 177392
rect 310738 20080 311358 177392
<< obsm4 >>
rect 8339 177472 313293 197437
rect 8339 20000 22658 177472
rect 23438 20000 40658 177472
rect 41438 20000 58658 177472
rect 59438 20000 76658 177472
rect 77438 20000 94658 177472
rect 95438 20000 112658 177472
rect 113438 20000 130658 177472
rect 131438 20000 148658 177472
rect 149438 20000 166658 177472
rect 167438 20000 184658 177472
rect 185438 20000 202658 177472
rect 203438 20000 220658 177472
rect 221438 20000 238658 177472
rect 239438 20000 256658 177472
rect 257438 20000 274658 177472
rect 275438 20000 292658 177472
rect 293438 20000 310658 177472
rect 311438 20000 313293 177472
rect 8339 851 313293 20000
<< labels >>
rlabel metal3 s 316356 104048 316756 104168 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 316356 114928 316756 115048 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 316356 125808 316756 125928 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 316356 136688 316756 136808 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 316356 147568 316756 147688 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 316356 158448 316756 158568 6 A0[5]
port 6 nsew signal input
rlabel metal3 s 316356 169328 316756 169448 6 A0[6]
port 7 nsew signal input
rlabel metal3 s 316356 180208 316756 180328 6 A0[7]
port 8 nsew signal input
rlabel metal3 s 316356 191088 316756 191208 6 A0[8]
port 9 nsew signal input
rlabel metal3 s 0 98608 400 98728 6 CLK
port 10 nsew signal input
rlabel metal2 s 4710 0 4766 400 6 Di0[0]
port 11 nsew signal input
rlabel metal2 s 53470 0 53526 400 6 Di0[10]
port 12 nsew signal input
rlabel metal2 s 58346 0 58402 400 6 Di0[11]
port 13 nsew signal input
rlabel metal2 s 63222 0 63278 400 6 Di0[12]
port 14 nsew signal input
rlabel metal2 s 68098 0 68154 400 6 Di0[13]
port 15 nsew signal input
rlabel metal2 s 72974 0 73030 400 6 Di0[14]
port 16 nsew signal input
rlabel metal2 s 77850 0 77906 400 6 Di0[15]
port 17 nsew signal input
rlabel metal2 s 82726 0 82782 400 6 Di0[16]
port 18 nsew signal input
rlabel metal2 s 87602 0 87658 400 6 Di0[17]
port 19 nsew signal input
rlabel metal2 s 92478 0 92534 400 6 Di0[18]
port 20 nsew signal input
rlabel metal2 s 97354 0 97410 400 6 Di0[19]
port 21 nsew signal input
rlabel metal2 s 9586 0 9642 400 6 Di0[1]
port 22 nsew signal input
rlabel metal2 s 102230 0 102286 400 6 Di0[20]
port 23 nsew signal input
rlabel metal2 s 107106 0 107162 400 6 Di0[21]
port 24 nsew signal input
rlabel metal2 s 111982 0 112038 400 6 Di0[22]
port 25 nsew signal input
rlabel metal2 s 116858 0 116914 400 6 Di0[23]
port 26 nsew signal input
rlabel metal2 s 121734 0 121790 400 6 Di0[24]
port 27 nsew signal input
rlabel metal2 s 126610 0 126666 400 6 Di0[25]
port 28 nsew signal input
rlabel metal2 s 131486 0 131542 400 6 Di0[26]
port 29 nsew signal input
rlabel metal2 s 136362 0 136418 400 6 Di0[27]
port 30 nsew signal input
rlabel metal2 s 141238 0 141294 400 6 Di0[28]
port 31 nsew signal input
rlabel metal2 s 146114 0 146170 400 6 Di0[29]
port 32 nsew signal input
rlabel metal2 s 14462 0 14518 400 6 Di0[2]
port 33 nsew signal input
rlabel metal2 s 150990 0 151046 400 6 Di0[30]
port 34 nsew signal input
rlabel metal2 s 155866 0 155922 400 6 Di0[31]
port 35 nsew signal input
rlabel metal2 s 160742 0 160798 400 6 Di0[32]
port 36 nsew signal input
rlabel metal2 s 165618 0 165674 400 6 Di0[33]
port 37 nsew signal input
rlabel metal2 s 170494 0 170550 400 6 Di0[34]
port 38 nsew signal input
rlabel metal2 s 175370 0 175426 400 6 Di0[35]
port 39 nsew signal input
rlabel metal2 s 180246 0 180302 400 6 Di0[36]
port 40 nsew signal input
rlabel metal2 s 185122 0 185178 400 6 Di0[37]
port 41 nsew signal input
rlabel metal2 s 189998 0 190054 400 6 Di0[38]
port 42 nsew signal input
rlabel metal2 s 194874 0 194930 400 6 Di0[39]
port 43 nsew signal input
rlabel metal2 s 19338 0 19394 400 6 Di0[3]
port 44 nsew signal input
rlabel metal2 s 199750 0 199806 400 6 Di0[40]
port 45 nsew signal input
rlabel metal2 s 204626 0 204682 400 6 Di0[41]
port 46 nsew signal input
rlabel metal2 s 209502 0 209558 400 6 Di0[42]
port 47 nsew signal input
rlabel metal2 s 214378 0 214434 400 6 Di0[43]
port 48 nsew signal input
rlabel metal2 s 219254 0 219310 400 6 Di0[44]
port 49 nsew signal input
rlabel metal2 s 224130 0 224186 400 6 Di0[45]
port 50 nsew signal input
rlabel metal2 s 229006 0 229062 400 6 Di0[46]
port 51 nsew signal input
rlabel metal2 s 233882 0 233938 400 6 Di0[47]
port 52 nsew signal input
rlabel metal2 s 238758 0 238814 400 6 Di0[48]
port 53 nsew signal input
rlabel metal2 s 243634 0 243690 400 6 Di0[49]
port 54 nsew signal input
rlabel metal2 s 24214 0 24270 400 6 Di0[4]
port 55 nsew signal input
rlabel metal2 s 248510 0 248566 400 6 Di0[50]
port 56 nsew signal input
rlabel metal2 s 253386 0 253442 400 6 Di0[51]
port 57 nsew signal input
rlabel metal2 s 258262 0 258318 400 6 Di0[52]
port 58 nsew signal input
rlabel metal2 s 263138 0 263194 400 6 Di0[53]
port 59 nsew signal input
rlabel metal2 s 268014 0 268070 400 6 Di0[54]
port 60 nsew signal input
rlabel metal2 s 272890 0 272946 400 6 Di0[55]
port 61 nsew signal input
rlabel metal2 s 277766 0 277822 400 6 Di0[56]
port 62 nsew signal input
rlabel metal2 s 282642 0 282698 400 6 Di0[57]
port 63 nsew signal input
rlabel metal2 s 287518 0 287574 400 6 Di0[58]
port 64 nsew signal input
rlabel metal2 s 292394 0 292450 400 6 Di0[59]
port 65 nsew signal input
rlabel metal2 s 29090 0 29146 400 6 Di0[5]
port 66 nsew signal input
rlabel metal2 s 297270 0 297326 400 6 Di0[60]
port 67 nsew signal input
rlabel metal2 s 302146 0 302202 400 6 Di0[61]
port 68 nsew signal input
rlabel metal2 s 307022 0 307078 400 6 Di0[62]
port 69 nsew signal input
rlabel metal2 s 311898 0 311954 400 6 Di0[63]
port 70 nsew signal input
rlabel metal2 s 33966 0 34022 400 6 Di0[6]
port 71 nsew signal input
rlabel metal2 s 38842 0 38898 400 6 Di0[7]
port 72 nsew signal input
rlabel metal2 s 43718 0 43774 400 6 Di0[8]
port 73 nsew signal input
rlabel metal2 s 48594 0 48650 400 6 Di0[9]
port 74 nsew signal input
rlabel metal2 s 4710 197072 4766 197472 6 Do0[0]
port 75 nsew signal output
rlabel metal2 s 53470 197072 53526 197472 6 Do0[10]
port 76 nsew signal output
rlabel metal2 s 58346 197072 58402 197472 6 Do0[11]
port 77 nsew signal output
rlabel metal2 s 63222 197072 63278 197472 6 Do0[12]
port 78 nsew signal output
rlabel metal2 s 68098 197072 68154 197472 6 Do0[13]
port 79 nsew signal output
rlabel metal2 s 72974 197072 73030 197472 6 Do0[14]
port 80 nsew signal output
rlabel metal2 s 77850 197072 77906 197472 6 Do0[15]
port 81 nsew signal output
rlabel metal2 s 82726 197072 82782 197472 6 Do0[16]
port 82 nsew signal output
rlabel metal2 s 87602 197072 87658 197472 6 Do0[17]
port 83 nsew signal output
rlabel metal2 s 92478 197072 92534 197472 6 Do0[18]
port 84 nsew signal output
rlabel metal2 s 97354 197072 97410 197472 6 Do0[19]
port 85 nsew signal output
rlabel metal2 s 9586 197072 9642 197472 6 Do0[1]
port 86 nsew signal output
rlabel metal2 s 102230 197072 102286 197472 6 Do0[20]
port 87 nsew signal output
rlabel metal2 s 107106 197072 107162 197472 6 Do0[21]
port 88 nsew signal output
rlabel metal2 s 111982 197072 112038 197472 6 Do0[22]
port 89 nsew signal output
rlabel metal2 s 116858 197072 116914 197472 6 Do0[23]
port 90 nsew signal output
rlabel metal2 s 121734 197072 121790 197472 6 Do0[24]
port 91 nsew signal output
rlabel metal2 s 126610 197072 126666 197472 6 Do0[25]
port 92 nsew signal output
rlabel metal2 s 131486 197072 131542 197472 6 Do0[26]
port 93 nsew signal output
rlabel metal2 s 136362 197072 136418 197472 6 Do0[27]
port 94 nsew signal output
rlabel metal2 s 141238 197072 141294 197472 6 Do0[28]
port 95 nsew signal output
rlabel metal2 s 146114 197072 146170 197472 6 Do0[29]
port 96 nsew signal output
rlabel metal2 s 14462 197072 14518 197472 6 Do0[2]
port 97 nsew signal output
rlabel metal2 s 150990 197072 151046 197472 6 Do0[30]
port 98 nsew signal output
rlabel metal2 s 155866 197072 155922 197472 6 Do0[31]
port 99 nsew signal output
rlabel metal2 s 160742 197072 160798 197472 6 Do0[32]
port 100 nsew signal output
rlabel metal2 s 165618 197072 165674 197472 6 Do0[33]
port 101 nsew signal output
rlabel metal2 s 170494 197072 170550 197472 6 Do0[34]
port 102 nsew signal output
rlabel metal2 s 175370 197072 175426 197472 6 Do0[35]
port 103 nsew signal output
rlabel metal2 s 180246 197072 180302 197472 6 Do0[36]
port 104 nsew signal output
rlabel metal2 s 185122 197072 185178 197472 6 Do0[37]
port 105 nsew signal output
rlabel metal2 s 189998 197072 190054 197472 6 Do0[38]
port 106 nsew signal output
rlabel metal2 s 194874 197072 194930 197472 6 Do0[39]
port 107 nsew signal output
rlabel metal2 s 19338 197072 19394 197472 6 Do0[3]
port 108 nsew signal output
rlabel metal2 s 199750 197072 199806 197472 6 Do0[40]
port 109 nsew signal output
rlabel metal2 s 204626 197072 204682 197472 6 Do0[41]
port 110 nsew signal output
rlabel metal2 s 209502 197072 209558 197472 6 Do0[42]
port 111 nsew signal output
rlabel metal2 s 214378 197072 214434 197472 6 Do0[43]
port 112 nsew signal output
rlabel metal2 s 219254 197072 219310 197472 6 Do0[44]
port 113 nsew signal output
rlabel metal2 s 224130 197072 224186 197472 6 Do0[45]
port 114 nsew signal output
rlabel metal2 s 229006 197072 229062 197472 6 Do0[46]
port 115 nsew signal output
rlabel metal2 s 233882 197072 233938 197472 6 Do0[47]
port 116 nsew signal output
rlabel metal2 s 238758 197072 238814 197472 6 Do0[48]
port 117 nsew signal output
rlabel metal2 s 243634 197072 243690 197472 6 Do0[49]
port 118 nsew signal output
rlabel metal2 s 24214 197072 24270 197472 6 Do0[4]
port 119 nsew signal output
rlabel metal2 s 248510 197072 248566 197472 6 Do0[50]
port 120 nsew signal output
rlabel metal2 s 253386 197072 253442 197472 6 Do0[51]
port 121 nsew signal output
rlabel metal2 s 258262 197072 258318 197472 6 Do0[52]
port 122 nsew signal output
rlabel metal2 s 263138 197072 263194 197472 6 Do0[53]
port 123 nsew signal output
rlabel metal2 s 268014 197072 268070 197472 6 Do0[54]
port 124 nsew signal output
rlabel metal2 s 272890 197072 272946 197472 6 Do0[55]
port 125 nsew signal output
rlabel metal2 s 277766 197072 277822 197472 6 Do0[56]
port 126 nsew signal output
rlabel metal2 s 282642 197072 282698 197472 6 Do0[57]
port 127 nsew signal output
rlabel metal2 s 287518 197072 287574 197472 6 Do0[58]
port 128 nsew signal output
rlabel metal2 s 292394 197072 292450 197472 6 Do0[59]
port 129 nsew signal output
rlabel metal2 s 29090 197072 29146 197472 6 Do0[5]
port 130 nsew signal output
rlabel metal2 s 297270 197072 297326 197472 6 Do0[60]
port 131 nsew signal output
rlabel metal2 s 302146 197072 302202 197472 6 Do0[61]
port 132 nsew signal output
rlabel metal2 s 307022 197072 307078 197472 6 Do0[62]
port 133 nsew signal output
rlabel metal2 s 311898 197072 311954 197472 6 Do0[63]
port 134 nsew signal output
rlabel metal2 s 33966 197072 34022 197472 6 Do0[6]
port 135 nsew signal output
rlabel metal2 s 38842 197072 38898 197472 6 Do0[7]
port 136 nsew signal output
rlabel metal2 s 43718 197072 43774 197472 6 Do0[8]
port 137 nsew signal output
rlabel metal2 s 48594 197072 48650 197472 6 Do0[9]
port 138 nsew signal output
rlabel metal3 s 316356 6128 316756 6248 6 EN0
port 139 nsew signal input
rlabel metal4 s 22738 20080 23358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 58738 20080 59358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 94738 20080 95358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 130738 20080 131358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 166738 20080 167358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 202738 20080 203358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 238738 20080 239358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 274738 20080 275358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 310738 20080 311358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 4738 20080 5358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 40738 20080 41358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 76738 20080 77358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 112738 20080 113358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 148738 20080 149358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 184738 20080 185358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 220738 20080 221358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 256738 20080 257358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 292738 20080 293358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal3 s 316356 17008 316756 17128 6 WE0[0]
port 142 nsew signal input
rlabel metal3 s 316356 27888 316756 28008 6 WE0[1]
port 143 nsew signal input
rlabel metal3 s 316356 38768 316756 38888 6 WE0[2]
port 144 nsew signal input
rlabel metal3 s 316356 49648 316756 49768 6 WE0[3]
port 145 nsew signal input
rlabel metal3 s 316356 60528 316756 60648 6 WE0[4]
port 146 nsew signal input
rlabel metal3 s 316356 71408 316756 71528 6 WE0[5]
port 147 nsew signal input
rlabel metal3 s 316356 82288 316756 82408 6 WE0[6]
port 148 nsew signal input
rlabel metal3 s 316356 93168 316756 93288 6 WE0[7]
port 149 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 316756 197472
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 189974424
string GDS_FILE /mnt/dffram/build/512x64_DEFAULT/openlane/runs/RUN_2022.09.07_08.02.44/results/signoff/RAM512.magic.gds
string GDS_START 165654
<< end >>

