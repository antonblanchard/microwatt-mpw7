VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiply_add_64x64
  CLASS BLOCK ;
  FOREIGN multiply_add_64x64 ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 98.970 10.640 102.070 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 10.640 282.070 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 10.640 462.070 487.120 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 8.970 10.640 12.070 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 10.640 192.070 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 10.640 372.070 487.120 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 33.360 500.000 33.960 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 67.360 500.000 67.960 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 70.760 500.000 71.360 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 74.160 500.000 74.760 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 77.560 500.000 78.160 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 80.960 500.000 81.560 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 84.360 500.000 84.960 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 87.760 500.000 88.360 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 91.160 500.000 91.760 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 94.560 500.000 95.160 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 97.960 500.000 98.560 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 36.760 500.000 37.360 ;
    END
  END a[1]
  PIN a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 101.360 500.000 101.960 ;
    END
  END a[20]
  PIN a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 104.760 500.000 105.360 ;
    END
  END a[21]
  PIN a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 108.160 500.000 108.760 ;
    END
  END a[22]
  PIN a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 111.560 500.000 112.160 ;
    END
  END a[23]
  PIN a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 114.960 500.000 115.560 ;
    END
  END a[24]
  PIN a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 118.360 500.000 118.960 ;
    END
  END a[25]
  PIN a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 121.760 500.000 122.360 ;
    END
  END a[26]
  PIN a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 125.160 500.000 125.760 ;
    END
  END a[27]
  PIN a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 128.560 500.000 129.160 ;
    END
  END a[28]
  PIN a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 131.960 500.000 132.560 ;
    END
  END a[29]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 40.160 500.000 40.760 ;
    END
  END a[2]
  PIN a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 135.360 500.000 135.960 ;
    END
  END a[30]
  PIN a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 138.760 500.000 139.360 ;
    END
  END a[31]
  PIN a[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 142.160 500.000 142.760 ;
    END
  END a[32]
  PIN a[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 145.560 500.000 146.160 ;
    END
  END a[33]
  PIN a[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 148.960 500.000 149.560 ;
    END
  END a[34]
  PIN a[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 152.360 500.000 152.960 ;
    END
  END a[35]
  PIN a[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 155.760 500.000 156.360 ;
    END
  END a[36]
  PIN a[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 159.160 500.000 159.760 ;
    END
  END a[37]
  PIN a[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 162.560 500.000 163.160 ;
    END
  END a[38]
  PIN a[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 165.960 500.000 166.560 ;
    END
  END a[39]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 43.560 500.000 44.160 ;
    END
  END a[3]
  PIN a[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 169.360 500.000 169.960 ;
    END
  END a[40]
  PIN a[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 172.760 500.000 173.360 ;
    END
  END a[41]
  PIN a[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 176.160 500.000 176.760 ;
    END
  END a[42]
  PIN a[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 179.560 500.000 180.160 ;
    END
  END a[43]
  PIN a[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 182.960 500.000 183.560 ;
    END
  END a[44]
  PIN a[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 186.360 500.000 186.960 ;
    END
  END a[45]
  PIN a[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 189.760 500.000 190.360 ;
    END
  END a[46]
  PIN a[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 193.160 500.000 193.760 ;
    END
  END a[47]
  PIN a[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 196.560 500.000 197.160 ;
    END
  END a[48]
  PIN a[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 199.960 500.000 200.560 ;
    END
  END a[49]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 46.960 500.000 47.560 ;
    END
  END a[4]
  PIN a[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 203.360 500.000 203.960 ;
    END
  END a[50]
  PIN a[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 206.760 500.000 207.360 ;
    END
  END a[51]
  PIN a[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 210.160 500.000 210.760 ;
    END
  END a[52]
  PIN a[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 213.560 500.000 214.160 ;
    END
  END a[53]
  PIN a[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 216.960 500.000 217.560 ;
    END
  END a[54]
  PIN a[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 220.360 500.000 220.960 ;
    END
  END a[55]
  PIN a[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 223.760 500.000 224.360 ;
    END
  END a[56]
  PIN a[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 227.160 500.000 227.760 ;
    END
  END a[57]
  PIN a[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 230.560 500.000 231.160 ;
    END
  END a[58]
  PIN a[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 233.960 500.000 234.560 ;
    END
  END a[59]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 50.360 500.000 50.960 ;
    END
  END a[5]
  PIN a[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 237.360 500.000 237.960 ;
    END
  END a[60]
  PIN a[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 240.760 500.000 241.360 ;
    END
  END a[61]
  PIN a[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 244.160 500.000 244.760 ;
    END
  END a[62]
  PIN a[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 247.560 500.000 248.160 ;
    END
  END a[63]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 53.760 500.000 54.360 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 57.160 500.000 57.760 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 60.560 500.000 61.160 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 63.960 500.000 64.560 ;
    END
  END a[9]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 250.960 500.000 251.560 ;
    END
  END b[0]
  PIN b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 284.960 500.000 285.560 ;
    END
  END b[10]
  PIN b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 288.360 500.000 288.960 ;
    END
  END b[11]
  PIN b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 291.760 500.000 292.360 ;
    END
  END b[12]
  PIN b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 295.160 500.000 295.760 ;
    END
  END b[13]
  PIN b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 298.560 500.000 299.160 ;
    END
  END b[14]
  PIN b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 301.960 500.000 302.560 ;
    END
  END b[15]
  PIN b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 305.360 500.000 305.960 ;
    END
  END b[16]
  PIN b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 308.760 500.000 309.360 ;
    END
  END b[17]
  PIN b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 312.160 500.000 312.760 ;
    END
  END b[18]
  PIN b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 315.560 500.000 316.160 ;
    END
  END b[19]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 254.360 500.000 254.960 ;
    END
  END b[1]
  PIN b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 318.960 500.000 319.560 ;
    END
  END b[20]
  PIN b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 322.360 500.000 322.960 ;
    END
  END b[21]
  PIN b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 325.760 500.000 326.360 ;
    END
  END b[22]
  PIN b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 329.160 500.000 329.760 ;
    END
  END b[23]
  PIN b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 332.560 500.000 333.160 ;
    END
  END b[24]
  PIN b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 335.960 500.000 336.560 ;
    END
  END b[25]
  PIN b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 339.360 500.000 339.960 ;
    END
  END b[26]
  PIN b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 342.760 500.000 343.360 ;
    END
  END b[27]
  PIN b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 346.160 500.000 346.760 ;
    END
  END b[28]
  PIN b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 349.560 500.000 350.160 ;
    END
  END b[29]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 257.760 500.000 258.360 ;
    END
  END b[2]
  PIN b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 352.960 500.000 353.560 ;
    END
  END b[30]
  PIN b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 356.360 500.000 356.960 ;
    END
  END b[31]
  PIN b[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 359.760 500.000 360.360 ;
    END
  END b[32]
  PIN b[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 363.160 500.000 363.760 ;
    END
  END b[33]
  PIN b[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 366.560 500.000 367.160 ;
    END
  END b[34]
  PIN b[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 369.960 500.000 370.560 ;
    END
  END b[35]
  PIN b[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 373.360 500.000 373.960 ;
    END
  END b[36]
  PIN b[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 376.760 500.000 377.360 ;
    END
  END b[37]
  PIN b[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 380.160 500.000 380.760 ;
    END
  END b[38]
  PIN b[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 383.560 500.000 384.160 ;
    END
  END b[39]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 261.160 500.000 261.760 ;
    END
  END b[3]
  PIN b[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 386.960 500.000 387.560 ;
    END
  END b[40]
  PIN b[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 390.360 500.000 390.960 ;
    END
  END b[41]
  PIN b[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 393.760 500.000 394.360 ;
    END
  END b[42]
  PIN b[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 397.160 500.000 397.760 ;
    END
  END b[43]
  PIN b[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 400.560 500.000 401.160 ;
    END
  END b[44]
  PIN b[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 403.960 500.000 404.560 ;
    END
  END b[45]
  PIN b[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 407.360 500.000 407.960 ;
    END
  END b[46]
  PIN b[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 410.760 500.000 411.360 ;
    END
  END b[47]
  PIN b[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 414.160 500.000 414.760 ;
    END
  END b[48]
  PIN b[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 417.560 500.000 418.160 ;
    END
  END b[49]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 264.560 500.000 265.160 ;
    END
  END b[4]
  PIN b[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 420.960 500.000 421.560 ;
    END
  END b[50]
  PIN b[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 424.360 500.000 424.960 ;
    END
  END b[51]
  PIN b[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 427.760 500.000 428.360 ;
    END
  END b[52]
  PIN b[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 431.160 500.000 431.760 ;
    END
  END b[53]
  PIN b[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 434.560 500.000 435.160 ;
    END
  END b[54]
  PIN b[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 437.960 500.000 438.560 ;
    END
  END b[55]
  PIN b[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 441.360 500.000 441.960 ;
    END
  END b[56]
  PIN b[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 444.760 500.000 445.360 ;
    END
  END b[57]
  PIN b[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 448.160 500.000 448.760 ;
    END
  END b[58]
  PIN b[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 451.560 500.000 452.160 ;
    END
  END b[59]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 267.960 500.000 268.560 ;
    END
  END b[5]
  PIN b[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 454.960 500.000 455.560 ;
    END
  END b[60]
  PIN b[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 458.360 500.000 458.960 ;
    END
  END b[61]
  PIN b[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 461.760 500.000 462.360 ;
    END
  END b[62]
  PIN b[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 465.160 500.000 465.760 ;
    END
  END b[63]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 271.360 500.000 271.960 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 274.760 500.000 275.360 ;
    END
  END b[7]
  PIN b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 278.160 500.000 278.760 ;
    END
  END b[8]
  PIN b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 281.560 500.000 282.160 ;
    END
  END b[9]
  PIN c[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END c[0]
  PIN c[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END c[100]
  PIN c[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END c[101]
  PIN c[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END c[102]
  PIN c[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 0.000 395.510 4.000 ;
    END
  END c[103]
  PIN c[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END c[104]
  PIN c[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END c[105]
  PIN c[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END c[106]
  PIN c[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END c[107]
  PIN c[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END c[108]
  PIN c[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END c[109]
  PIN c[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END c[10]
  PIN c[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END c[110]
  PIN c[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END c[111]
  PIN c[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END c[112]
  PIN c[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END c[113]
  PIN c[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 0.000 435.990 4.000 ;
    END
  END c[114]
  PIN c[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END c[115]
  PIN c[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END c[116]
  PIN c[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END c[117]
  PIN c[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END c[118]
  PIN c[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END c[119]
  PIN c[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END c[11]
  PIN c[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END c[120]
  PIN c[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END c[121]
  PIN c[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 0.000 465.430 4.000 ;
    END
  END c[122]
  PIN c[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END c[123]
  PIN c[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 0.000 472.790 4.000 ;
    END
  END c[124]
  PIN c[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END c[125]
  PIN c[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END c[126]
  PIN c[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 0.000 483.830 4.000 ;
    END
  END c[127]
  PIN c[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END c[12]
  PIN c[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END c[13]
  PIN c[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END c[14]
  PIN c[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END c[15]
  PIN c[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END c[16]
  PIN c[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END c[17]
  PIN c[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END c[18]
  PIN c[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END c[19]
  PIN c[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END c[1]
  PIN c[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END c[20]
  PIN c[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END c[21]
  PIN c[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END c[22]
  PIN c[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END c[23]
  PIN c[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END c[24]
  PIN c[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END c[25]
  PIN c[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END c[26]
  PIN c[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END c[27]
  PIN c[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END c[28]
  PIN c[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END c[29]
  PIN c[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END c[2]
  PIN c[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END c[30]
  PIN c[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END c[31]
  PIN c[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END c[32]
  PIN c[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END c[33]
  PIN c[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END c[34]
  PIN c[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END c[35]
  PIN c[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END c[36]
  PIN c[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END c[37]
  PIN c[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END c[38]
  PIN c[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END c[39]
  PIN c[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END c[3]
  PIN c[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END c[40]
  PIN c[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END c[41]
  PIN c[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END c[42]
  PIN c[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END c[43]
  PIN c[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END c[44]
  PIN c[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END c[45]
  PIN c[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END c[46]
  PIN c[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END c[47]
  PIN c[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END c[48]
  PIN c[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END c[49]
  PIN c[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END c[4]
  PIN c[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END c[50]
  PIN c[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END c[51]
  PIN c[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END c[52]
  PIN c[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END c[53]
  PIN c[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END c[54]
  PIN c[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END c[55]
  PIN c[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END c[56]
  PIN c[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END c[57]
  PIN c[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END c[58]
  PIN c[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END c[59]
  PIN c[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END c[5]
  PIN c[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END c[60]
  PIN c[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END c[61]
  PIN c[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END c[62]
  PIN c[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END c[63]
  PIN c[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END c[64]
  PIN c[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END c[65]
  PIN c[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 4.000 ;
    END
  END c[66]
  PIN c[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END c[67]
  PIN c[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END c[68]
  PIN c[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END c[69]
  PIN c[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END c[6]
  PIN c[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END c[70]
  PIN c[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 4.000 ;
    END
  END c[71]
  PIN c[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END c[72]
  PIN c[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END c[73]
  PIN c[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END c[74]
  PIN c[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END c[75]
  PIN c[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END c[76]
  PIN c[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END c[77]
  PIN c[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END c[78]
  PIN c[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END c[79]
  PIN c[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END c[7]
  PIN c[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END c[80]
  PIN c[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END c[81]
  PIN c[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END c[82]
  PIN c[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END c[83]
  PIN c[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END c[84]
  PIN c[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END c[85]
  PIN c[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END c[86]
  PIN c[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END c[87]
  PIN c[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END c[88]
  PIN c[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END c[89]
  PIN c[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END c[8]
  PIN c[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END c[90]
  PIN c[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END c[91]
  PIN c[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END c[92]
  PIN c[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END c[93]
  PIN c[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END c[94]
  PIN c[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END c[95]
  PIN c[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END c[96]
  PIN c[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END c[97]
  PIN c[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END c[98]
  PIN c[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END c[99]
  PIN c[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END c[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 496.000 487.510 500.000 ;
    END
  END clk
  PIN o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 496.000 12.790 500.000 ;
    END
  END o[0]
  PIN o[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 496.000 380.790 500.000 ;
    END
  END o[100]
  PIN o[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 496.000 384.470 500.000 ;
    END
  END o[101]
  PIN o[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 496.000 388.150 500.000 ;
    END
  END o[102]
  PIN o[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 496.000 391.830 500.000 ;
    END
  END o[103]
  PIN o[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 496.000 395.510 500.000 ;
    END
  END o[104]
  PIN o[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 496.000 399.190 500.000 ;
    END
  END o[105]
  PIN o[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 496.000 402.870 500.000 ;
    END
  END o[106]
  PIN o[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 496.000 406.550 500.000 ;
    END
  END o[107]
  PIN o[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 496.000 410.230 500.000 ;
    END
  END o[108]
  PIN o[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 496.000 413.910 500.000 ;
    END
  END o[109]
  PIN o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 496.000 49.590 500.000 ;
    END
  END o[10]
  PIN o[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 496.000 417.590 500.000 ;
    END
  END o[110]
  PIN o[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 496.000 421.270 500.000 ;
    END
  END o[111]
  PIN o[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 496.000 424.950 500.000 ;
    END
  END o[112]
  PIN o[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 496.000 428.630 500.000 ;
    END
  END o[113]
  PIN o[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 496.000 432.310 500.000 ;
    END
  END o[114]
  PIN o[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 496.000 435.990 500.000 ;
    END
  END o[115]
  PIN o[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 496.000 439.670 500.000 ;
    END
  END o[116]
  PIN o[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 496.000 443.350 500.000 ;
    END
  END o[117]
  PIN o[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 496.000 447.030 500.000 ;
    END
  END o[118]
  PIN o[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 496.000 450.710 500.000 ;
    END
  END o[119]
  PIN o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 496.000 53.270 500.000 ;
    END
  END o[11]
  PIN o[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 496.000 454.390 500.000 ;
    END
  END o[120]
  PIN o[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 496.000 458.070 500.000 ;
    END
  END o[121]
  PIN o[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 496.000 461.750 500.000 ;
    END
  END o[122]
  PIN o[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 496.000 465.430 500.000 ;
    END
  END o[123]
  PIN o[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 496.000 469.110 500.000 ;
    END
  END o[124]
  PIN o[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 496.000 472.790 500.000 ;
    END
  END o[125]
  PIN o[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 496.000 476.470 500.000 ;
    END
  END o[126]
  PIN o[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 496.000 480.150 500.000 ;
    END
  END o[127]
  PIN o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 496.000 56.950 500.000 ;
    END
  END o[12]
  PIN o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 496.000 60.630 500.000 ;
    END
  END o[13]
  PIN o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 496.000 64.310 500.000 ;
    END
  END o[14]
  PIN o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 496.000 67.990 500.000 ;
    END
  END o[15]
  PIN o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 496.000 71.670 500.000 ;
    END
  END o[16]
  PIN o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 496.000 75.350 500.000 ;
    END
  END o[17]
  PIN o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 496.000 79.030 500.000 ;
    END
  END o[18]
  PIN o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 496.000 82.710 500.000 ;
    END
  END o[19]
  PIN o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 496.000 16.470 500.000 ;
    END
  END o[1]
  PIN o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 496.000 86.390 500.000 ;
    END
  END o[20]
  PIN o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 496.000 90.070 500.000 ;
    END
  END o[21]
  PIN o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 496.000 93.750 500.000 ;
    END
  END o[22]
  PIN o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 496.000 97.430 500.000 ;
    END
  END o[23]
  PIN o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 496.000 101.110 500.000 ;
    END
  END o[24]
  PIN o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 496.000 104.790 500.000 ;
    END
  END o[25]
  PIN o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 496.000 108.470 500.000 ;
    END
  END o[26]
  PIN o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 496.000 112.150 500.000 ;
    END
  END o[27]
  PIN o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 496.000 115.830 500.000 ;
    END
  END o[28]
  PIN o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 496.000 119.510 500.000 ;
    END
  END o[29]
  PIN o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 496.000 20.150 500.000 ;
    END
  END o[2]
  PIN o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 496.000 123.190 500.000 ;
    END
  END o[30]
  PIN o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 496.000 126.870 500.000 ;
    END
  END o[31]
  PIN o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 496.000 130.550 500.000 ;
    END
  END o[32]
  PIN o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 496.000 134.230 500.000 ;
    END
  END o[33]
  PIN o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 496.000 137.910 500.000 ;
    END
  END o[34]
  PIN o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 496.000 141.590 500.000 ;
    END
  END o[35]
  PIN o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 496.000 145.270 500.000 ;
    END
  END o[36]
  PIN o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 496.000 148.950 500.000 ;
    END
  END o[37]
  PIN o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 496.000 152.630 500.000 ;
    END
  END o[38]
  PIN o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 496.000 156.310 500.000 ;
    END
  END o[39]
  PIN o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 496.000 23.830 500.000 ;
    END
  END o[3]
  PIN o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 496.000 159.990 500.000 ;
    END
  END o[40]
  PIN o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 496.000 163.670 500.000 ;
    END
  END o[41]
  PIN o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 496.000 167.350 500.000 ;
    END
  END o[42]
  PIN o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 496.000 171.030 500.000 ;
    END
  END o[43]
  PIN o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 496.000 174.710 500.000 ;
    END
  END o[44]
  PIN o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 496.000 178.390 500.000 ;
    END
  END o[45]
  PIN o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 496.000 182.070 500.000 ;
    END
  END o[46]
  PIN o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 496.000 185.750 500.000 ;
    END
  END o[47]
  PIN o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 496.000 189.430 500.000 ;
    END
  END o[48]
  PIN o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 496.000 193.110 500.000 ;
    END
  END o[49]
  PIN o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 496.000 27.510 500.000 ;
    END
  END o[4]
  PIN o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 496.000 196.790 500.000 ;
    END
  END o[50]
  PIN o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 496.000 200.470 500.000 ;
    END
  END o[51]
  PIN o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 496.000 204.150 500.000 ;
    END
  END o[52]
  PIN o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 496.000 207.830 500.000 ;
    END
  END o[53]
  PIN o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 496.000 211.510 500.000 ;
    END
  END o[54]
  PIN o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 496.000 215.190 500.000 ;
    END
  END o[55]
  PIN o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 496.000 218.870 500.000 ;
    END
  END o[56]
  PIN o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 496.000 222.550 500.000 ;
    END
  END o[57]
  PIN o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 496.000 226.230 500.000 ;
    END
  END o[58]
  PIN o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 496.000 229.910 500.000 ;
    END
  END o[59]
  PIN o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 496.000 31.190 500.000 ;
    END
  END o[5]
  PIN o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 496.000 233.590 500.000 ;
    END
  END o[60]
  PIN o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 496.000 237.270 500.000 ;
    END
  END o[61]
  PIN o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 496.000 240.950 500.000 ;
    END
  END o[62]
  PIN o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 496.000 244.630 500.000 ;
    END
  END o[63]
  PIN o[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 496.000 248.310 500.000 ;
    END
  END o[64]
  PIN o[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 496.000 251.990 500.000 ;
    END
  END o[65]
  PIN o[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 496.000 255.670 500.000 ;
    END
  END o[66]
  PIN o[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 496.000 259.350 500.000 ;
    END
  END o[67]
  PIN o[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 496.000 263.030 500.000 ;
    END
  END o[68]
  PIN o[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 496.000 266.710 500.000 ;
    END
  END o[69]
  PIN o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 496.000 34.870 500.000 ;
    END
  END o[6]
  PIN o[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 496.000 270.390 500.000 ;
    END
  END o[70]
  PIN o[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 496.000 274.070 500.000 ;
    END
  END o[71]
  PIN o[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 496.000 277.750 500.000 ;
    END
  END o[72]
  PIN o[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 496.000 281.430 500.000 ;
    END
  END o[73]
  PIN o[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 496.000 285.110 500.000 ;
    END
  END o[74]
  PIN o[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 496.000 288.790 500.000 ;
    END
  END o[75]
  PIN o[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 496.000 292.470 500.000 ;
    END
  END o[76]
  PIN o[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 496.000 296.150 500.000 ;
    END
  END o[77]
  PIN o[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 496.000 299.830 500.000 ;
    END
  END o[78]
  PIN o[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 496.000 303.510 500.000 ;
    END
  END o[79]
  PIN o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 496.000 38.550 500.000 ;
    END
  END o[7]
  PIN o[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 496.000 307.190 500.000 ;
    END
  END o[80]
  PIN o[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 496.000 310.870 500.000 ;
    END
  END o[81]
  PIN o[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 496.000 314.550 500.000 ;
    END
  END o[82]
  PIN o[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 496.000 318.230 500.000 ;
    END
  END o[83]
  PIN o[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 496.000 321.910 500.000 ;
    END
  END o[84]
  PIN o[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 496.000 325.590 500.000 ;
    END
  END o[85]
  PIN o[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 496.000 329.270 500.000 ;
    END
  END o[86]
  PIN o[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 496.000 332.950 500.000 ;
    END
  END o[87]
  PIN o[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 496.000 336.630 500.000 ;
    END
  END o[88]
  PIN o[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 496.000 340.310 500.000 ;
    END
  END o[89]
  PIN o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 496.000 42.230 500.000 ;
    END
  END o[8]
  PIN o[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 496.000 343.990 500.000 ;
    END
  END o[90]
  PIN o[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 496.000 347.670 500.000 ;
    END
  END o[91]
  PIN o[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 496.000 351.350 500.000 ;
    END
  END o[92]
  PIN o[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 496.000 355.030 500.000 ;
    END
  END o[93]
  PIN o[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 496.000 358.710 500.000 ;
    END
  END o[94]
  PIN o[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 496.000 362.390 500.000 ;
    END
  END o[95]
  PIN o[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 496.000 366.070 500.000 ;
    END
  END o[96]
  PIN o[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 496.000 369.750 500.000 ;
    END
  END o[97]
  PIN o[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 496.000 373.430 500.000 ;
    END
  END o[98]
  PIN o[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 496.000 377.110 500.000 ;
    END
  END o[99]
  PIN o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 496.000 45.910 500.000 ;
    END
  END o[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 496.000 483.830 500.000 ;
    END
  END rst
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 1.450 8.540 499.950 492.620 ;
      LAYER met2 ;
        RECT 1.010 495.720 12.230 496.810 ;
        RECT 13.070 495.720 15.910 496.810 ;
        RECT 16.750 495.720 19.590 496.810 ;
        RECT 20.430 495.720 23.270 496.810 ;
        RECT 24.110 495.720 26.950 496.810 ;
        RECT 27.790 495.720 30.630 496.810 ;
        RECT 31.470 495.720 34.310 496.810 ;
        RECT 35.150 495.720 37.990 496.810 ;
        RECT 38.830 495.720 41.670 496.810 ;
        RECT 42.510 495.720 45.350 496.810 ;
        RECT 46.190 495.720 49.030 496.810 ;
        RECT 49.870 495.720 52.710 496.810 ;
        RECT 53.550 495.720 56.390 496.810 ;
        RECT 57.230 495.720 60.070 496.810 ;
        RECT 60.910 495.720 63.750 496.810 ;
        RECT 64.590 495.720 67.430 496.810 ;
        RECT 68.270 495.720 71.110 496.810 ;
        RECT 71.950 495.720 74.790 496.810 ;
        RECT 75.630 495.720 78.470 496.810 ;
        RECT 79.310 495.720 82.150 496.810 ;
        RECT 82.990 495.720 85.830 496.810 ;
        RECT 86.670 495.720 89.510 496.810 ;
        RECT 90.350 495.720 93.190 496.810 ;
        RECT 94.030 495.720 96.870 496.810 ;
        RECT 97.710 495.720 100.550 496.810 ;
        RECT 101.390 495.720 104.230 496.810 ;
        RECT 105.070 495.720 107.910 496.810 ;
        RECT 108.750 495.720 111.590 496.810 ;
        RECT 112.430 495.720 115.270 496.810 ;
        RECT 116.110 495.720 118.950 496.810 ;
        RECT 119.790 495.720 122.630 496.810 ;
        RECT 123.470 495.720 126.310 496.810 ;
        RECT 127.150 495.720 129.990 496.810 ;
        RECT 130.830 495.720 133.670 496.810 ;
        RECT 134.510 495.720 137.350 496.810 ;
        RECT 138.190 495.720 141.030 496.810 ;
        RECT 141.870 495.720 144.710 496.810 ;
        RECT 145.550 495.720 148.390 496.810 ;
        RECT 149.230 495.720 152.070 496.810 ;
        RECT 152.910 495.720 155.750 496.810 ;
        RECT 156.590 495.720 159.430 496.810 ;
        RECT 160.270 495.720 163.110 496.810 ;
        RECT 163.950 495.720 166.790 496.810 ;
        RECT 167.630 495.720 170.470 496.810 ;
        RECT 171.310 495.720 174.150 496.810 ;
        RECT 174.990 495.720 177.830 496.810 ;
        RECT 178.670 495.720 181.510 496.810 ;
        RECT 182.350 495.720 185.190 496.810 ;
        RECT 186.030 495.720 188.870 496.810 ;
        RECT 189.710 495.720 192.550 496.810 ;
        RECT 193.390 495.720 196.230 496.810 ;
        RECT 197.070 495.720 199.910 496.810 ;
        RECT 200.750 495.720 203.590 496.810 ;
        RECT 204.430 495.720 207.270 496.810 ;
        RECT 208.110 495.720 210.950 496.810 ;
        RECT 211.790 495.720 214.630 496.810 ;
        RECT 215.470 495.720 218.310 496.810 ;
        RECT 219.150 495.720 221.990 496.810 ;
        RECT 222.830 495.720 225.670 496.810 ;
        RECT 226.510 495.720 229.350 496.810 ;
        RECT 230.190 495.720 233.030 496.810 ;
        RECT 233.870 495.720 236.710 496.810 ;
        RECT 237.550 495.720 240.390 496.810 ;
        RECT 241.230 495.720 244.070 496.810 ;
        RECT 244.910 495.720 247.750 496.810 ;
        RECT 248.590 495.720 251.430 496.810 ;
        RECT 252.270 495.720 255.110 496.810 ;
        RECT 255.950 495.720 258.790 496.810 ;
        RECT 259.630 495.720 262.470 496.810 ;
        RECT 263.310 495.720 266.150 496.810 ;
        RECT 266.990 495.720 269.830 496.810 ;
        RECT 270.670 495.720 273.510 496.810 ;
        RECT 274.350 495.720 277.190 496.810 ;
        RECT 278.030 495.720 280.870 496.810 ;
        RECT 281.710 495.720 284.550 496.810 ;
        RECT 285.390 495.720 288.230 496.810 ;
        RECT 289.070 495.720 291.910 496.810 ;
        RECT 292.750 495.720 295.590 496.810 ;
        RECT 296.430 495.720 299.270 496.810 ;
        RECT 300.110 495.720 302.950 496.810 ;
        RECT 303.790 495.720 306.630 496.810 ;
        RECT 307.470 495.720 310.310 496.810 ;
        RECT 311.150 495.720 313.990 496.810 ;
        RECT 314.830 495.720 317.670 496.810 ;
        RECT 318.510 495.720 321.350 496.810 ;
        RECT 322.190 495.720 325.030 496.810 ;
        RECT 325.870 495.720 328.710 496.810 ;
        RECT 329.550 495.720 332.390 496.810 ;
        RECT 333.230 495.720 336.070 496.810 ;
        RECT 336.910 495.720 339.750 496.810 ;
        RECT 340.590 495.720 343.430 496.810 ;
        RECT 344.270 495.720 347.110 496.810 ;
        RECT 347.950 495.720 350.790 496.810 ;
        RECT 351.630 495.720 354.470 496.810 ;
        RECT 355.310 495.720 358.150 496.810 ;
        RECT 358.990 495.720 361.830 496.810 ;
        RECT 362.670 495.720 365.510 496.810 ;
        RECT 366.350 495.720 369.190 496.810 ;
        RECT 370.030 495.720 372.870 496.810 ;
        RECT 373.710 495.720 376.550 496.810 ;
        RECT 377.390 495.720 380.230 496.810 ;
        RECT 381.070 495.720 383.910 496.810 ;
        RECT 384.750 495.720 387.590 496.810 ;
        RECT 388.430 495.720 391.270 496.810 ;
        RECT 392.110 495.720 394.950 496.810 ;
        RECT 395.790 495.720 398.630 496.810 ;
        RECT 399.470 495.720 402.310 496.810 ;
        RECT 403.150 495.720 405.990 496.810 ;
        RECT 406.830 495.720 409.670 496.810 ;
        RECT 410.510 495.720 413.350 496.810 ;
        RECT 414.190 495.720 417.030 496.810 ;
        RECT 417.870 495.720 420.710 496.810 ;
        RECT 421.550 495.720 424.390 496.810 ;
        RECT 425.230 495.720 428.070 496.810 ;
        RECT 428.910 495.720 431.750 496.810 ;
        RECT 432.590 495.720 435.430 496.810 ;
        RECT 436.270 495.720 439.110 496.810 ;
        RECT 439.950 495.720 442.790 496.810 ;
        RECT 443.630 495.720 446.470 496.810 ;
        RECT 447.310 495.720 450.150 496.810 ;
        RECT 450.990 495.720 453.830 496.810 ;
        RECT 454.670 495.720 457.510 496.810 ;
        RECT 458.350 495.720 461.190 496.810 ;
        RECT 462.030 495.720 464.870 496.810 ;
        RECT 465.710 495.720 468.550 496.810 ;
        RECT 469.390 495.720 472.230 496.810 ;
        RECT 473.070 495.720 475.910 496.810 ;
        RECT 476.750 495.720 479.590 496.810 ;
        RECT 480.430 495.720 483.270 496.810 ;
        RECT 484.110 495.720 486.950 496.810 ;
        RECT 487.790 495.720 499.930 496.810 ;
        RECT 1.010 4.280 499.930 495.720 ;
        RECT 1.010 3.670 15.910 4.280 ;
        RECT 16.750 3.670 19.590 4.280 ;
        RECT 20.430 3.670 23.270 4.280 ;
        RECT 24.110 3.670 26.950 4.280 ;
        RECT 27.790 3.670 30.630 4.280 ;
        RECT 31.470 3.670 34.310 4.280 ;
        RECT 35.150 3.670 37.990 4.280 ;
        RECT 38.830 3.670 41.670 4.280 ;
        RECT 42.510 3.670 45.350 4.280 ;
        RECT 46.190 3.670 49.030 4.280 ;
        RECT 49.870 3.670 52.710 4.280 ;
        RECT 53.550 3.670 56.390 4.280 ;
        RECT 57.230 3.670 60.070 4.280 ;
        RECT 60.910 3.670 63.750 4.280 ;
        RECT 64.590 3.670 67.430 4.280 ;
        RECT 68.270 3.670 71.110 4.280 ;
        RECT 71.950 3.670 74.790 4.280 ;
        RECT 75.630 3.670 78.470 4.280 ;
        RECT 79.310 3.670 82.150 4.280 ;
        RECT 82.990 3.670 85.830 4.280 ;
        RECT 86.670 3.670 89.510 4.280 ;
        RECT 90.350 3.670 93.190 4.280 ;
        RECT 94.030 3.670 96.870 4.280 ;
        RECT 97.710 3.670 100.550 4.280 ;
        RECT 101.390 3.670 104.230 4.280 ;
        RECT 105.070 3.670 107.910 4.280 ;
        RECT 108.750 3.670 111.590 4.280 ;
        RECT 112.430 3.670 115.270 4.280 ;
        RECT 116.110 3.670 118.950 4.280 ;
        RECT 119.790 3.670 122.630 4.280 ;
        RECT 123.470 3.670 126.310 4.280 ;
        RECT 127.150 3.670 129.990 4.280 ;
        RECT 130.830 3.670 133.670 4.280 ;
        RECT 134.510 3.670 137.350 4.280 ;
        RECT 138.190 3.670 141.030 4.280 ;
        RECT 141.870 3.670 144.710 4.280 ;
        RECT 145.550 3.670 148.390 4.280 ;
        RECT 149.230 3.670 152.070 4.280 ;
        RECT 152.910 3.670 155.750 4.280 ;
        RECT 156.590 3.670 159.430 4.280 ;
        RECT 160.270 3.670 163.110 4.280 ;
        RECT 163.950 3.670 166.790 4.280 ;
        RECT 167.630 3.670 170.470 4.280 ;
        RECT 171.310 3.670 174.150 4.280 ;
        RECT 174.990 3.670 177.830 4.280 ;
        RECT 178.670 3.670 181.510 4.280 ;
        RECT 182.350 3.670 185.190 4.280 ;
        RECT 186.030 3.670 188.870 4.280 ;
        RECT 189.710 3.670 192.550 4.280 ;
        RECT 193.390 3.670 196.230 4.280 ;
        RECT 197.070 3.670 199.910 4.280 ;
        RECT 200.750 3.670 203.590 4.280 ;
        RECT 204.430 3.670 207.270 4.280 ;
        RECT 208.110 3.670 210.950 4.280 ;
        RECT 211.790 3.670 214.630 4.280 ;
        RECT 215.470 3.670 218.310 4.280 ;
        RECT 219.150 3.670 221.990 4.280 ;
        RECT 222.830 3.670 225.670 4.280 ;
        RECT 226.510 3.670 229.350 4.280 ;
        RECT 230.190 3.670 233.030 4.280 ;
        RECT 233.870 3.670 236.710 4.280 ;
        RECT 237.550 3.670 240.390 4.280 ;
        RECT 241.230 3.670 244.070 4.280 ;
        RECT 244.910 3.670 247.750 4.280 ;
        RECT 248.590 3.670 251.430 4.280 ;
        RECT 252.270 3.670 255.110 4.280 ;
        RECT 255.950 3.670 258.790 4.280 ;
        RECT 259.630 3.670 262.470 4.280 ;
        RECT 263.310 3.670 266.150 4.280 ;
        RECT 266.990 3.670 269.830 4.280 ;
        RECT 270.670 3.670 273.510 4.280 ;
        RECT 274.350 3.670 277.190 4.280 ;
        RECT 278.030 3.670 280.870 4.280 ;
        RECT 281.710 3.670 284.550 4.280 ;
        RECT 285.390 3.670 288.230 4.280 ;
        RECT 289.070 3.670 291.910 4.280 ;
        RECT 292.750 3.670 295.590 4.280 ;
        RECT 296.430 3.670 299.270 4.280 ;
        RECT 300.110 3.670 302.950 4.280 ;
        RECT 303.790 3.670 306.630 4.280 ;
        RECT 307.470 3.670 310.310 4.280 ;
        RECT 311.150 3.670 313.990 4.280 ;
        RECT 314.830 3.670 317.670 4.280 ;
        RECT 318.510 3.670 321.350 4.280 ;
        RECT 322.190 3.670 325.030 4.280 ;
        RECT 325.870 3.670 328.710 4.280 ;
        RECT 329.550 3.670 332.390 4.280 ;
        RECT 333.230 3.670 336.070 4.280 ;
        RECT 336.910 3.670 339.750 4.280 ;
        RECT 340.590 3.670 343.430 4.280 ;
        RECT 344.270 3.670 347.110 4.280 ;
        RECT 347.950 3.670 350.790 4.280 ;
        RECT 351.630 3.670 354.470 4.280 ;
        RECT 355.310 3.670 358.150 4.280 ;
        RECT 358.990 3.670 361.830 4.280 ;
        RECT 362.670 3.670 365.510 4.280 ;
        RECT 366.350 3.670 369.190 4.280 ;
        RECT 370.030 3.670 372.870 4.280 ;
        RECT 373.710 3.670 376.550 4.280 ;
        RECT 377.390 3.670 380.230 4.280 ;
        RECT 381.070 3.670 383.910 4.280 ;
        RECT 384.750 3.670 387.590 4.280 ;
        RECT 388.430 3.670 391.270 4.280 ;
        RECT 392.110 3.670 394.950 4.280 ;
        RECT 395.790 3.670 398.630 4.280 ;
        RECT 399.470 3.670 402.310 4.280 ;
        RECT 403.150 3.670 405.990 4.280 ;
        RECT 406.830 3.670 409.670 4.280 ;
        RECT 410.510 3.670 413.350 4.280 ;
        RECT 414.190 3.670 417.030 4.280 ;
        RECT 417.870 3.670 420.710 4.280 ;
        RECT 421.550 3.670 424.390 4.280 ;
        RECT 425.230 3.670 428.070 4.280 ;
        RECT 428.910 3.670 431.750 4.280 ;
        RECT 432.590 3.670 435.430 4.280 ;
        RECT 436.270 3.670 439.110 4.280 ;
        RECT 439.950 3.670 442.790 4.280 ;
        RECT 443.630 3.670 446.470 4.280 ;
        RECT 447.310 3.670 450.150 4.280 ;
        RECT 450.990 3.670 453.830 4.280 ;
        RECT 454.670 3.670 457.510 4.280 ;
        RECT 458.350 3.670 461.190 4.280 ;
        RECT 462.030 3.670 464.870 4.280 ;
        RECT 465.710 3.670 468.550 4.280 ;
        RECT 469.390 3.670 472.230 4.280 ;
        RECT 473.070 3.670 475.910 4.280 ;
        RECT 476.750 3.670 479.590 4.280 ;
        RECT 480.430 3.670 483.270 4.280 ;
        RECT 484.110 3.670 499.930 4.280 ;
      LAYER met3 ;
        RECT 0.985 466.160 499.955 494.180 ;
        RECT 0.985 464.760 495.600 466.160 ;
        RECT 0.985 462.760 499.955 464.760 ;
        RECT 0.985 461.360 495.600 462.760 ;
        RECT 0.985 459.360 499.955 461.360 ;
        RECT 0.985 457.960 495.600 459.360 ;
        RECT 0.985 455.960 499.955 457.960 ;
        RECT 0.985 454.560 495.600 455.960 ;
        RECT 0.985 452.560 499.955 454.560 ;
        RECT 0.985 451.160 495.600 452.560 ;
        RECT 0.985 449.160 499.955 451.160 ;
        RECT 0.985 447.760 495.600 449.160 ;
        RECT 0.985 445.760 499.955 447.760 ;
        RECT 0.985 444.360 495.600 445.760 ;
        RECT 0.985 442.360 499.955 444.360 ;
        RECT 0.985 440.960 495.600 442.360 ;
        RECT 0.985 438.960 499.955 440.960 ;
        RECT 0.985 437.560 495.600 438.960 ;
        RECT 0.985 435.560 499.955 437.560 ;
        RECT 0.985 434.160 495.600 435.560 ;
        RECT 0.985 432.160 499.955 434.160 ;
        RECT 0.985 430.760 495.600 432.160 ;
        RECT 0.985 428.760 499.955 430.760 ;
        RECT 0.985 427.360 495.600 428.760 ;
        RECT 0.985 425.360 499.955 427.360 ;
        RECT 0.985 423.960 495.600 425.360 ;
        RECT 0.985 421.960 499.955 423.960 ;
        RECT 0.985 420.560 495.600 421.960 ;
        RECT 0.985 418.560 499.955 420.560 ;
        RECT 0.985 417.160 495.600 418.560 ;
        RECT 0.985 415.160 499.955 417.160 ;
        RECT 0.985 413.760 495.600 415.160 ;
        RECT 0.985 411.760 499.955 413.760 ;
        RECT 0.985 410.360 495.600 411.760 ;
        RECT 0.985 408.360 499.955 410.360 ;
        RECT 0.985 406.960 495.600 408.360 ;
        RECT 0.985 404.960 499.955 406.960 ;
        RECT 0.985 403.560 495.600 404.960 ;
        RECT 0.985 401.560 499.955 403.560 ;
        RECT 0.985 400.160 495.600 401.560 ;
        RECT 0.985 398.160 499.955 400.160 ;
        RECT 0.985 396.760 495.600 398.160 ;
        RECT 0.985 394.760 499.955 396.760 ;
        RECT 0.985 393.360 495.600 394.760 ;
        RECT 0.985 391.360 499.955 393.360 ;
        RECT 0.985 389.960 495.600 391.360 ;
        RECT 0.985 387.960 499.955 389.960 ;
        RECT 0.985 386.560 495.600 387.960 ;
        RECT 0.985 384.560 499.955 386.560 ;
        RECT 0.985 383.160 495.600 384.560 ;
        RECT 0.985 381.160 499.955 383.160 ;
        RECT 0.985 379.760 495.600 381.160 ;
        RECT 0.985 377.760 499.955 379.760 ;
        RECT 0.985 376.360 495.600 377.760 ;
        RECT 0.985 374.360 499.955 376.360 ;
        RECT 0.985 372.960 495.600 374.360 ;
        RECT 0.985 370.960 499.955 372.960 ;
        RECT 0.985 369.560 495.600 370.960 ;
        RECT 0.985 367.560 499.955 369.560 ;
        RECT 0.985 366.160 495.600 367.560 ;
        RECT 0.985 364.160 499.955 366.160 ;
        RECT 0.985 362.760 495.600 364.160 ;
        RECT 0.985 360.760 499.955 362.760 ;
        RECT 0.985 359.360 495.600 360.760 ;
        RECT 0.985 357.360 499.955 359.360 ;
        RECT 0.985 355.960 495.600 357.360 ;
        RECT 0.985 353.960 499.955 355.960 ;
        RECT 0.985 352.560 495.600 353.960 ;
        RECT 0.985 350.560 499.955 352.560 ;
        RECT 0.985 349.160 495.600 350.560 ;
        RECT 0.985 347.160 499.955 349.160 ;
        RECT 0.985 345.760 495.600 347.160 ;
        RECT 0.985 343.760 499.955 345.760 ;
        RECT 0.985 342.360 495.600 343.760 ;
        RECT 0.985 340.360 499.955 342.360 ;
        RECT 0.985 338.960 495.600 340.360 ;
        RECT 0.985 336.960 499.955 338.960 ;
        RECT 0.985 335.560 495.600 336.960 ;
        RECT 0.985 333.560 499.955 335.560 ;
        RECT 0.985 332.160 495.600 333.560 ;
        RECT 0.985 330.160 499.955 332.160 ;
        RECT 0.985 328.760 495.600 330.160 ;
        RECT 0.985 326.760 499.955 328.760 ;
        RECT 0.985 325.360 495.600 326.760 ;
        RECT 0.985 323.360 499.955 325.360 ;
        RECT 0.985 321.960 495.600 323.360 ;
        RECT 0.985 319.960 499.955 321.960 ;
        RECT 0.985 318.560 495.600 319.960 ;
        RECT 0.985 316.560 499.955 318.560 ;
        RECT 0.985 315.160 495.600 316.560 ;
        RECT 0.985 313.160 499.955 315.160 ;
        RECT 0.985 311.760 495.600 313.160 ;
        RECT 0.985 309.760 499.955 311.760 ;
        RECT 0.985 308.360 495.600 309.760 ;
        RECT 0.985 306.360 499.955 308.360 ;
        RECT 0.985 304.960 495.600 306.360 ;
        RECT 0.985 302.960 499.955 304.960 ;
        RECT 0.985 301.560 495.600 302.960 ;
        RECT 0.985 299.560 499.955 301.560 ;
        RECT 0.985 298.160 495.600 299.560 ;
        RECT 0.985 296.160 499.955 298.160 ;
        RECT 0.985 294.760 495.600 296.160 ;
        RECT 0.985 292.760 499.955 294.760 ;
        RECT 0.985 291.360 495.600 292.760 ;
        RECT 0.985 289.360 499.955 291.360 ;
        RECT 0.985 287.960 495.600 289.360 ;
        RECT 0.985 285.960 499.955 287.960 ;
        RECT 0.985 284.560 495.600 285.960 ;
        RECT 0.985 282.560 499.955 284.560 ;
        RECT 0.985 281.160 495.600 282.560 ;
        RECT 0.985 279.160 499.955 281.160 ;
        RECT 0.985 277.760 495.600 279.160 ;
        RECT 0.985 275.760 499.955 277.760 ;
        RECT 0.985 274.360 495.600 275.760 ;
        RECT 0.985 272.360 499.955 274.360 ;
        RECT 0.985 270.960 495.600 272.360 ;
        RECT 0.985 268.960 499.955 270.960 ;
        RECT 0.985 267.560 495.600 268.960 ;
        RECT 0.985 265.560 499.955 267.560 ;
        RECT 0.985 264.160 495.600 265.560 ;
        RECT 0.985 262.160 499.955 264.160 ;
        RECT 0.985 260.760 495.600 262.160 ;
        RECT 0.985 258.760 499.955 260.760 ;
        RECT 0.985 257.360 495.600 258.760 ;
        RECT 0.985 255.360 499.955 257.360 ;
        RECT 0.985 253.960 495.600 255.360 ;
        RECT 0.985 251.960 499.955 253.960 ;
        RECT 0.985 250.560 495.600 251.960 ;
        RECT 0.985 248.560 499.955 250.560 ;
        RECT 0.985 247.160 495.600 248.560 ;
        RECT 0.985 245.160 499.955 247.160 ;
        RECT 0.985 243.760 495.600 245.160 ;
        RECT 0.985 241.760 499.955 243.760 ;
        RECT 0.985 240.360 495.600 241.760 ;
        RECT 0.985 238.360 499.955 240.360 ;
        RECT 0.985 236.960 495.600 238.360 ;
        RECT 0.985 234.960 499.955 236.960 ;
        RECT 0.985 233.560 495.600 234.960 ;
        RECT 0.985 231.560 499.955 233.560 ;
        RECT 0.985 230.160 495.600 231.560 ;
        RECT 0.985 228.160 499.955 230.160 ;
        RECT 0.985 226.760 495.600 228.160 ;
        RECT 0.985 224.760 499.955 226.760 ;
        RECT 0.985 223.360 495.600 224.760 ;
        RECT 0.985 221.360 499.955 223.360 ;
        RECT 0.985 219.960 495.600 221.360 ;
        RECT 0.985 217.960 499.955 219.960 ;
        RECT 0.985 216.560 495.600 217.960 ;
        RECT 0.985 214.560 499.955 216.560 ;
        RECT 0.985 213.160 495.600 214.560 ;
        RECT 0.985 211.160 499.955 213.160 ;
        RECT 0.985 209.760 495.600 211.160 ;
        RECT 0.985 207.760 499.955 209.760 ;
        RECT 0.985 206.360 495.600 207.760 ;
        RECT 0.985 204.360 499.955 206.360 ;
        RECT 0.985 202.960 495.600 204.360 ;
        RECT 0.985 200.960 499.955 202.960 ;
        RECT 0.985 199.560 495.600 200.960 ;
        RECT 0.985 197.560 499.955 199.560 ;
        RECT 0.985 196.160 495.600 197.560 ;
        RECT 0.985 194.160 499.955 196.160 ;
        RECT 0.985 192.760 495.600 194.160 ;
        RECT 0.985 190.760 499.955 192.760 ;
        RECT 0.985 189.360 495.600 190.760 ;
        RECT 0.985 187.360 499.955 189.360 ;
        RECT 0.985 185.960 495.600 187.360 ;
        RECT 0.985 183.960 499.955 185.960 ;
        RECT 0.985 182.560 495.600 183.960 ;
        RECT 0.985 180.560 499.955 182.560 ;
        RECT 0.985 179.160 495.600 180.560 ;
        RECT 0.985 177.160 499.955 179.160 ;
        RECT 0.985 175.760 495.600 177.160 ;
        RECT 0.985 173.760 499.955 175.760 ;
        RECT 0.985 172.360 495.600 173.760 ;
        RECT 0.985 170.360 499.955 172.360 ;
        RECT 0.985 168.960 495.600 170.360 ;
        RECT 0.985 166.960 499.955 168.960 ;
        RECT 0.985 165.560 495.600 166.960 ;
        RECT 0.985 163.560 499.955 165.560 ;
        RECT 0.985 162.160 495.600 163.560 ;
        RECT 0.985 160.160 499.955 162.160 ;
        RECT 0.985 158.760 495.600 160.160 ;
        RECT 0.985 156.760 499.955 158.760 ;
        RECT 0.985 155.360 495.600 156.760 ;
        RECT 0.985 153.360 499.955 155.360 ;
        RECT 0.985 151.960 495.600 153.360 ;
        RECT 0.985 149.960 499.955 151.960 ;
        RECT 0.985 148.560 495.600 149.960 ;
        RECT 0.985 146.560 499.955 148.560 ;
        RECT 0.985 145.160 495.600 146.560 ;
        RECT 0.985 143.160 499.955 145.160 ;
        RECT 0.985 141.760 495.600 143.160 ;
        RECT 0.985 139.760 499.955 141.760 ;
        RECT 0.985 138.360 495.600 139.760 ;
        RECT 0.985 136.360 499.955 138.360 ;
        RECT 0.985 134.960 495.600 136.360 ;
        RECT 0.985 132.960 499.955 134.960 ;
        RECT 0.985 131.560 495.600 132.960 ;
        RECT 0.985 129.560 499.955 131.560 ;
        RECT 0.985 128.160 495.600 129.560 ;
        RECT 0.985 126.160 499.955 128.160 ;
        RECT 0.985 124.760 495.600 126.160 ;
        RECT 0.985 122.760 499.955 124.760 ;
        RECT 0.985 121.360 495.600 122.760 ;
        RECT 0.985 119.360 499.955 121.360 ;
        RECT 0.985 117.960 495.600 119.360 ;
        RECT 0.985 115.960 499.955 117.960 ;
        RECT 0.985 114.560 495.600 115.960 ;
        RECT 0.985 112.560 499.955 114.560 ;
        RECT 0.985 111.160 495.600 112.560 ;
        RECT 0.985 109.160 499.955 111.160 ;
        RECT 0.985 107.760 495.600 109.160 ;
        RECT 0.985 105.760 499.955 107.760 ;
        RECT 0.985 104.360 495.600 105.760 ;
        RECT 0.985 102.360 499.955 104.360 ;
        RECT 0.985 100.960 495.600 102.360 ;
        RECT 0.985 98.960 499.955 100.960 ;
        RECT 0.985 97.560 495.600 98.960 ;
        RECT 0.985 95.560 499.955 97.560 ;
        RECT 0.985 94.160 495.600 95.560 ;
        RECT 0.985 92.160 499.955 94.160 ;
        RECT 0.985 90.760 495.600 92.160 ;
        RECT 0.985 88.760 499.955 90.760 ;
        RECT 0.985 87.360 495.600 88.760 ;
        RECT 0.985 85.360 499.955 87.360 ;
        RECT 0.985 83.960 495.600 85.360 ;
        RECT 0.985 81.960 499.955 83.960 ;
        RECT 0.985 80.560 495.600 81.960 ;
        RECT 0.985 78.560 499.955 80.560 ;
        RECT 0.985 77.160 495.600 78.560 ;
        RECT 0.985 75.160 499.955 77.160 ;
        RECT 0.985 73.760 495.600 75.160 ;
        RECT 0.985 71.760 499.955 73.760 ;
        RECT 0.985 70.360 495.600 71.760 ;
        RECT 0.985 68.360 499.955 70.360 ;
        RECT 0.985 66.960 495.600 68.360 ;
        RECT 0.985 64.960 499.955 66.960 ;
        RECT 0.985 63.560 495.600 64.960 ;
        RECT 0.985 61.560 499.955 63.560 ;
        RECT 0.985 60.160 495.600 61.560 ;
        RECT 0.985 58.160 499.955 60.160 ;
        RECT 0.985 56.760 495.600 58.160 ;
        RECT 0.985 54.760 499.955 56.760 ;
        RECT 0.985 53.360 495.600 54.760 ;
        RECT 0.985 51.360 499.955 53.360 ;
        RECT 0.985 49.960 495.600 51.360 ;
        RECT 0.985 47.960 499.955 49.960 ;
        RECT 0.985 46.560 495.600 47.960 ;
        RECT 0.985 44.560 499.955 46.560 ;
        RECT 0.985 43.160 495.600 44.560 ;
        RECT 0.985 41.160 499.955 43.160 ;
        RECT 0.985 39.760 495.600 41.160 ;
        RECT 0.985 37.760 499.955 39.760 ;
        RECT 0.985 36.360 495.600 37.760 ;
        RECT 0.985 34.360 499.955 36.360 ;
        RECT 0.985 32.960 495.600 34.360 ;
        RECT 0.985 6.975 499.955 32.960 ;
      LAYER met4 ;
        RECT 2.135 487.520 492.825 494.185 ;
        RECT 2.135 10.240 8.570 487.520 ;
        RECT 12.470 10.240 98.570 487.520 ;
        RECT 102.470 10.240 188.570 487.520 ;
        RECT 192.470 10.240 278.570 487.520 ;
        RECT 282.470 10.240 368.570 487.520 ;
        RECT 372.470 10.240 458.570 487.520 ;
        RECT 462.470 10.240 492.825 487.520 ;
        RECT 2.135 6.975 492.825 10.240 ;
  END
END multiply_add_64x64
END LIBRARY

