VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiply_add_64x64
  CLASS BLOCK ;
  FOREIGN multiply_add_64x64 ;
  ORIGIN 0.000 0.000 ;
  SIZE 550.000 BY 550.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 98.970 10.640 102.070 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 10.640 282.070 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 10.640 462.070 538.800 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 8.970 10.640 12.070 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 10.640 192.070 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 10.640 372.070 538.800 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 17.720 550.000 18.320 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 58.520 550.000 59.120 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 62.600 550.000 63.200 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 66.680 550.000 67.280 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 70.760 550.000 71.360 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 74.840 550.000 75.440 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 78.920 550.000 79.520 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 83.000 550.000 83.600 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 87.080 550.000 87.680 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 91.160 550.000 91.760 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 95.240 550.000 95.840 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 21.800 550.000 22.400 ;
    END
  END a[1]
  PIN a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 99.320 550.000 99.920 ;
    END
  END a[20]
  PIN a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 103.400 550.000 104.000 ;
    END
  END a[21]
  PIN a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 107.480 550.000 108.080 ;
    END
  END a[22]
  PIN a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 111.560 550.000 112.160 ;
    END
  END a[23]
  PIN a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 115.640 550.000 116.240 ;
    END
  END a[24]
  PIN a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 119.720 550.000 120.320 ;
    END
  END a[25]
  PIN a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 123.800 550.000 124.400 ;
    END
  END a[26]
  PIN a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 127.880 550.000 128.480 ;
    END
  END a[27]
  PIN a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 131.960 550.000 132.560 ;
    END
  END a[28]
  PIN a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 136.040 550.000 136.640 ;
    END
  END a[29]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 25.880 550.000 26.480 ;
    END
  END a[2]
  PIN a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 140.120 550.000 140.720 ;
    END
  END a[30]
  PIN a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 144.200 550.000 144.800 ;
    END
  END a[31]
  PIN a[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 148.280 550.000 148.880 ;
    END
  END a[32]
  PIN a[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 152.360 550.000 152.960 ;
    END
  END a[33]
  PIN a[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 156.440 550.000 157.040 ;
    END
  END a[34]
  PIN a[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 160.520 550.000 161.120 ;
    END
  END a[35]
  PIN a[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 164.600 550.000 165.200 ;
    END
  END a[36]
  PIN a[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 168.680 550.000 169.280 ;
    END
  END a[37]
  PIN a[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 172.760 550.000 173.360 ;
    END
  END a[38]
  PIN a[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 176.840 550.000 177.440 ;
    END
  END a[39]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 29.960 550.000 30.560 ;
    END
  END a[3]
  PIN a[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 180.920 550.000 181.520 ;
    END
  END a[40]
  PIN a[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 185.000 550.000 185.600 ;
    END
  END a[41]
  PIN a[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 189.080 550.000 189.680 ;
    END
  END a[42]
  PIN a[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 193.160 550.000 193.760 ;
    END
  END a[43]
  PIN a[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 197.240 550.000 197.840 ;
    END
  END a[44]
  PIN a[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 201.320 550.000 201.920 ;
    END
  END a[45]
  PIN a[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 205.400 550.000 206.000 ;
    END
  END a[46]
  PIN a[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 209.480 550.000 210.080 ;
    END
  END a[47]
  PIN a[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 213.560 550.000 214.160 ;
    END
  END a[48]
  PIN a[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 217.640 550.000 218.240 ;
    END
  END a[49]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 34.040 550.000 34.640 ;
    END
  END a[4]
  PIN a[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 221.720 550.000 222.320 ;
    END
  END a[50]
  PIN a[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 225.800 550.000 226.400 ;
    END
  END a[51]
  PIN a[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 229.880 550.000 230.480 ;
    END
  END a[52]
  PIN a[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 233.960 550.000 234.560 ;
    END
  END a[53]
  PIN a[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 238.040 550.000 238.640 ;
    END
  END a[54]
  PIN a[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 242.120 550.000 242.720 ;
    END
  END a[55]
  PIN a[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 246.200 550.000 246.800 ;
    END
  END a[56]
  PIN a[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 250.280 550.000 250.880 ;
    END
  END a[57]
  PIN a[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 254.360 550.000 254.960 ;
    END
  END a[58]
  PIN a[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 258.440 550.000 259.040 ;
    END
  END a[59]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 38.120 550.000 38.720 ;
    END
  END a[5]
  PIN a[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 262.520 550.000 263.120 ;
    END
  END a[60]
  PIN a[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 266.600 550.000 267.200 ;
    END
  END a[61]
  PIN a[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 270.680 550.000 271.280 ;
    END
  END a[62]
  PIN a[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 274.760 550.000 275.360 ;
    END
  END a[63]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 42.200 550.000 42.800 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 46.280 550.000 46.880 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 50.360 550.000 50.960 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 54.440 550.000 55.040 ;
    END
  END a[9]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 278.840 550.000 279.440 ;
    END
  END b[0]
  PIN b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 319.640 550.000 320.240 ;
    END
  END b[10]
  PIN b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 323.720 550.000 324.320 ;
    END
  END b[11]
  PIN b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 327.800 550.000 328.400 ;
    END
  END b[12]
  PIN b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 331.880 550.000 332.480 ;
    END
  END b[13]
  PIN b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 335.960 550.000 336.560 ;
    END
  END b[14]
  PIN b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 340.040 550.000 340.640 ;
    END
  END b[15]
  PIN b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 344.120 550.000 344.720 ;
    END
  END b[16]
  PIN b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 348.200 550.000 348.800 ;
    END
  END b[17]
  PIN b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 352.280 550.000 352.880 ;
    END
  END b[18]
  PIN b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 356.360 550.000 356.960 ;
    END
  END b[19]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 282.920 550.000 283.520 ;
    END
  END b[1]
  PIN b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 360.440 550.000 361.040 ;
    END
  END b[20]
  PIN b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 364.520 550.000 365.120 ;
    END
  END b[21]
  PIN b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 368.600 550.000 369.200 ;
    END
  END b[22]
  PIN b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 372.680 550.000 373.280 ;
    END
  END b[23]
  PIN b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 376.760 550.000 377.360 ;
    END
  END b[24]
  PIN b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 380.840 550.000 381.440 ;
    END
  END b[25]
  PIN b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 384.920 550.000 385.520 ;
    END
  END b[26]
  PIN b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 389.000 550.000 389.600 ;
    END
  END b[27]
  PIN b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 393.080 550.000 393.680 ;
    END
  END b[28]
  PIN b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 397.160 550.000 397.760 ;
    END
  END b[29]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 287.000 550.000 287.600 ;
    END
  END b[2]
  PIN b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 401.240 550.000 401.840 ;
    END
  END b[30]
  PIN b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 405.320 550.000 405.920 ;
    END
  END b[31]
  PIN b[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 409.400 550.000 410.000 ;
    END
  END b[32]
  PIN b[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 413.480 550.000 414.080 ;
    END
  END b[33]
  PIN b[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 417.560 550.000 418.160 ;
    END
  END b[34]
  PIN b[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 421.640 550.000 422.240 ;
    END
  END b[35]
  PIN b[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 425.720 550.000 426.320 ;
    END
  END b[36]
  PIN b[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 429.800 550.000 430.400 ;
    END
  END b[37]
  PIN b[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 433.880 550.000 434.480 ;
    END
  END b[38]
  PIN b[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 437.960 550.000 438.560 ;
    END
  END b[39]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 291.080 550.000 291.680 ;
    END
  END b[3]
  PIN b[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 442.040 550.000 442.640 ;
    END
  END b[40]
  PIN b[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 446.120 550.000 446.720 ;
    END
  END b[41]
  PIN b[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 450.200 550.000 450.800 ;
    END
  END b[42]
  PIN b[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 454.280 550.000 454.880 ;
    END
  END b[43]
  PIN b[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 458.360 550.000 458.960 ;
    END
  END b[44]
  PIN b[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 462.440 550.000 463.040 ;
    END
  END b[45]
  PIN b[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 466.520 550.000 467.120 ;
    END
  END b[46]
  PIN b[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 470.600 550.000 471.200 ;
    END
  END b[47]
  PIN b[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 474.680 550.000 475.280 ;
    END
  END b[48]
  PIN b[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 478.760 550.000 479.360 ;
    END
  END b[49]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 295.160 550.000 295.760 ;
    END
  END b[4]
  PIN b[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 482.840 550.000 483.440 ;
    END
  END b[50]
  PIN b[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 486.920 550.000 487.520 ;
    END
  END b[51]
  PIN b[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 491.000 550.000 491.600 ;
    END
  END b[52]
  PIN b[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 495.080 550.000 495.680 ;
    END
  END b[53]
  PIN b[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 499.160 550.000 499.760 ;
    END
  END b[54]
  PIN b[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 503.240 550.000 503.840 ;
    END
  END b[55]
  PIN b[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 507.320 550.000 507.920 ;
    END
  END b[56]
  PIN b[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 511.400 550.000 512.000 ;
    END
  END b[57]
  PIN b[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 515.480 550.000 516.080 ;
    END
  END b[58]
  PIN b[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 519.560 550.000 520.160 ;
    END
  END b[59]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 299.240 550.000 299.840 ;
    END
  END b[5]
  PIN b[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 523.640 550.000 524.240 ;
    END
  END b[60]
  PIN b[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 527.720 550.000 528.320 ;
    END
  END b[61]
  PIN b[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 531.800 550.000 532.400 ;
    END
  END b[62]
  PIN b[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 535.880 550.000 536.480 ;
    END
  END b[63]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 303.320 550.000 303.920 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 307.400 550.000 308.000 ;
    END
  END b[7]
  PIN b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 311.480 550.000 312.080 ;
    END
  END b[8]
  PIN b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 315.560 550.000 316.160 ;
    END
  END b[9]
  PIN c[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END c[0]
  PIN c[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END c[100]
  PIN c[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END c[101]
  PIN c[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END c[102]
  PIN c[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END c[103]
  PIN c[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 4.000 ;
    END
  END c[104]
  PIN c[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END c[105]
  PIN c[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END c[106]
  PIN c[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 0.000 455.310 4.000 ;
    END
  END c[107]
  PIN c[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END c[108]
  PIN c[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 4.000 ;
    END
  END c[109]
  PIN c[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END c[10]
  PIN c[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END c[110]
  PIN c[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END c[111]
  PIN c[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 4.000 ;
    END
  END c[112]
  PIN c[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END c[113]
  PIN c[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END c[114]
  PIN c[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END c[115]
  PIN c[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END c[116]
  PIN c[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END c[117]
  PIN c[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END c[118]
  PIN c[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 4.000 ;
    END
  END c[119]
  PIN c[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END c[11]
  PIN c[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END c[120]
  PIN c[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 0.000 513.270 4.000 ;
    END
  END c[121]
  PIN c[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END c[122]
  PIN c[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END c[123]
  PIN c[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END c[124]
  PIN c[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END c[125]
  PIN c[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 4.000 ;
    END
  END c[126]
  PIN c[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END c[127]
  PIN c[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END c[12]
  PIN c[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END c[13]
  PIN c[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END c[14]
  PIN c[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END c[15]
  PIN c[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END c[16]
  PIN c[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END c[17]
  PIN c[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END c[18]
  PIN c[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END c[19]
  PIN c[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END c[1]
  PIN c[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END c[20]
  PIN c[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END c[21]
  PIN c[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END c[22]
  PIN c[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END c[23]
  PIN c[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END c[24]
  PIN c[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END c[25]
  PIN c[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END c[26]
  PIN c[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END c[27]
  PIN c[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END c[28]
  PIN c[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END c[29]
  PIN c[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END c[2]
  PIN c[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END c[30]
  PIN c[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END c[31]
  PIN c[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END c[32]
  PIN c[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END c[33]
  PIN c[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END c[34]
  PIN c[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END c[35]
  PIN c[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END c[36]
  PIN c[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END c[37]
  PIN c[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END c[38]
  PIN c[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END c[39]
  PIN c[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END c[3]
  PIN c[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END c[40]
  PIN c[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END c[41]
  PIN c[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END c[42]
  PIN c[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END c[43]
  PIN c[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END c[44]
  PIN c[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END c[45]
  PIN c[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END c[46]
  PIN c[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END c[47]
  PIN c[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END c[48]
  PIN c[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END c[49]
  PIN c[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END c[4]
  PIN c[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END c[50]
  PIN c[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END c[51]
  PIN c[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END c[52]
  PIN c[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END c[53]
  PIN c[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END c[54]
  PIN c[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END c[55]
  PIN c[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END c[56]
  PIN c[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END c[57]
  PIN c[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END c[58]
  PIN c[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END c[59]
  PIN c[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END c[5]
  PIN c[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END c[60]
  PIN c[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END c[61]
  PIN c[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END c[62]
  PIN c[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END c[63]
  PIN c[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END c[64]
  PIN c[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END c[65]
  PIN c[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END c[66]
  PIN c[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END c[67]
  PIN c[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END c[68]
  PIN c[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END c[69]
  PIN c[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END c[6]
  PIN c[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END c[70]
  PIN c[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END c[71]
  PIN c[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END c[72]
  PIN c[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END c[73]
  PIN c[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END c[74]
  PIN c[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END c[75]
  PIN c[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END c[76]
  PIN c[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END c[77]
  PIN c[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END c[78]
  PIN c[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END c[79]
  PIN c[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END c[7]
  PIN c[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END c[80]
  PIN c[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END c[81]
  PIN c[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END c[82]
  PIN c[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 4.000 ;
    END
  END c[83]
  PIN c[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END c[84]
  PIN c[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END c[85]
  PIN c[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END c[86]
  PIN c[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END c[87]
  PIN c[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END c[88]
  PIN c[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END c[89]
  PIN c[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END c[8]
  PIN c[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END c[90]
  PIN c[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 4.000 ;
    END
  END c[91]
  PIN c[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END c[92]
  PIN c[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END c[93]
  PIN c[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END c[94]
  PIN c[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 0.000 405.630 4.000 ;
    END
  END c[95]
  PIN c[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END c[96]
  PIN c[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END c[97]
  PIN c[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END c[98]
  PIN c[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END c[99]
  PIN c[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END c[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 13.640 550.000 14.240 ;
    END
  END clk
  PIN o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 546.000 10.030 550.000 ;
    END
  END o[0]
  PIN o[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 546.000 424.030 550.000 ;
    END
  END o[100]
  PIN o[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 546.000 428.170 550.000 ;
    END
  END o[101]
  PIN o[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 546.000 432.310 550.000 ;
    END
  END o[102]
  PIN o[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 546.000 436.450 550.000 ;
    END
  END o[103]
  PIN o[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 546.000 440.590 550.000 ;
    END
  END o[104]
  PIN o[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 546.000 444.730 550.000 ;
    END
  END o[105]
  PIN o[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 546.000 448.870 550.000 ;
    END
  END o[106]
  PIN o[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 546.000 453.010 550.000 ;
    END
  END o[107]
  PIN o[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 546.000 457.150 550.000 ;
    END
  END o[108]
  PIN o[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 546.000 461.290 550.000 ;
    END
  END o[109]
  PIN o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 546.000 51.430 550.000 ;
    END
  END o[10]
  PIN o[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 546.000 465.430 550.000 ;
    END
  END o[110]
  PIN o[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 546.000 469.570 550.000 ;
    END
  END o[111]
  PIN o[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 546.000 473.710 550.000 ;
    END
  END o[112]
  PIN o[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 546.000 477.850 550.000 ;
    END
  END o[113]
  PIN o[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 546.000 481.990 550.000 ;
    END
  END o[114]
  PIN o[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 546.000 486.130 550.000 ;
    END
  END o[115]
  PIN o[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 546.000 490.270 550.000 ;
    END
  END o[116]
  PIN o[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 546.000 494.410 550.000 ;
    END
  END o[117]
  PIN o[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 546.000 498.550 550.000 ;
    END
  END o[118]
  PIN o[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 546.000 502.690 550.000 ;
    END
  END o[119]
  PIN o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 546.000 55.570 550.000 ;
    END
  END o[11]
  PIN o[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 546.000 506.830 550.000 ;
    END
  END o[120]
  PIN o[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 546.000 510.970 550.000 ;
    END
  END o[121]
  PIN o[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 546.000 515.110 550.000 ;
    END
  END o[122]
  PIN o[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 546.000 519.250 550.000 ;
    END
  END o[123]
  PIN o[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 546.000 523.390 550.000 ;
    END
  END o[124]
  PIN o[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 546.000 527.530 550.000 ;
    END
  END o[125]
  PIN o[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 546.000 531.670 550.000 ;
    END
  END o[126]
  PIN o[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 546.000 535.810 550.000 ;
    END
  END o[127]
  PIN o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 546.000 59.710 550.000 ;
    END
  END o[12]
  PIN o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 546.000 63.850 550.000 ;
    END
  END o[13]
  PIN o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 546.000 67.990 550.000 ;
    END
  END o[14]
  PIN o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 546.000 72.130 550.000 ;
    END
  END o[15]
  PIN o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 546.000 76.270 550.000 ;
    END
  END o[16]
  PIN o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 546.000 80.410 550.000 ;
    END
  END o[17]
  PIN o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 546.000 84.550 550.000 ;
    END
  END o[18]
  PIN o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 546.000 88.690 550.000 ;
    END
  END o[19]
  PIN o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 546.000 14.170 550.000 ;
    END
  END o[1]
  PIN o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 546.000 92.830 550.000 ;
    END
  END o[20]
  PIN o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 546.000 96.970 550.000 ;
    END
  END o[21]
  PIN o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 546.000 101.110 550.000 ;
    END
  END o[22]
  PIN o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 546.000 105.250 550.000 ;
    END
  END o[23]
  PIN o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 546.000 109.390 550.000 ;
    END
  END o[24]
  PIN o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 546.000 113.530 550.000 ;
    END
  END o[25]
  PIN o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 546.000 117.670 550.000 ;
    END
  END o[26]
  PIN o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 546.000 121.810 550.000 ;
    END
  END o[27]
  PIN o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 546.000 125.950 550.000 ;
    END
  END o[28]
  PIN o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 546.000 130.090 550.000 ;
    END
  END o[29]
  PIN o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 546.000 18.310 550.000 ;
    END
  END o[2]
  PIN o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 546.000 134.230 550.000 ;
    END
  END o[30]
  PIN o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 546.000 138.370 550.000 ;
    END
  END o[31]
  PIN o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 546.000 142.510 550.000 ;
    END
  END o[32]
  PIN o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 546.000 146.650 550.000 ;
    END
  END o[33]
  PIN o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 546.000 150.790 550.000 ;
    END
  END o[34]
  PIN o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 546.000 154.930 550.000 ;
    END
  END o[35]
  PIN o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 546.000 159.070 550.000 ;
    END
  END o[36]
  PIN o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 546.000 163.210 550.000 ;
    END
  END o[37]
  PIN o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 546.000 167.350 550.000 ;
    END
  END o[38]
  PIN o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 546.000 171.490 550.000 ;
    END
  END o[39]
  PIN o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 546.000 22.450 550.000 ;
    END
  END o[3]
  PIN o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 546.000 175.630 550.000 ;
    END
  END o[40]
  PIN o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 546.000 179.770 550.000 ;
    END
  END o[41]
  PIN o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 546.000 183.910 550.000 ;
    END
  END o[42]
  PIN o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 546.000 188.050 550.000 ;
    END
  END o[43]
  PIN o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 546.000 192.190 550.000 ;
    END
  END o[44]
  PIN o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 546.000 196.330 550.000 ;
    END
  END o[45]
  PIN o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 546.000 200.470 550.000 ;
    END
  END o[46]
  PIN o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 546.000 204.610 550.000 ;
    END
  END o[47]
  PIN o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 546.000 208.750 550.000 ;
    END
  END o[48]
  PIN o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 546.000 212.890 550.000 ;
    END
  END o[49]
  PIN o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 546.000 26.590 550.000 ;
    END
  END o[4]
  PIN o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 546.000 217.030 550.000 ;
    END
  END o[50]
  PIN o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 546.000 221.170 550.000 ;
    END
  END o[51]
  PIN o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 546.000 225.310 550.000 ;
    END
  END o[52]
  PIN o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 546.000 229.450 550.000 ;
    END
  END o[53]
  PIN o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 546.000 233.590 550.000 ;
    END
  END o[54]
  PIN o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 546.000 237.730 550.000 ;
    END
  END o[55]
  PIN o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 546.000 241.870 550.000 ;
    END
  END o[56]
  PIN o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 546.000 246.010 550.000 ;
    END
  END o[57]
  PIN o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 546.000 250.150 550.000 ;
    END
  END o[58]
  PIN o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 546.000 254.290 550.000 ;
    END
  END o[59]
  PIN o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 546.000 30.730 550.000 ;
    END
  END o[5]
  PIN o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 546.000 258.430 550.000 ;
    END
  END o[60]
  PIN o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 546.000 262.570 550.000 ;
    END
  END o[61]
  PIN o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 546.000 266.710 550.000 ;
    END
  END o[62]
  PIN o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 546.000 270.850 550.000 ;
    END
  END o[63]
  PIN o[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 546.000 274.990 550.000 ;
    END
  END o[64]
  PIN o[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 546.000 279.130 550.000 ;
    END
  END o[65]
  PIN o[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 546.000 283.270 550.000 ;
    END
  END o[66]
  PIN o[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 546.000 287.410 550.000 ;
    END
  END o[67]
  PIN o[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 546.000 291.550 550.000 ;
    END
  END o[68]
  PIN o[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 546.000 295.690 550.000 ;
    END
  END o[69]
  PIN o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 546.000 34.870 550.000 ;
    END
  END o[6]
  PIN o[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 546.000 299.830 550.000 ;
    END
  END o[70]
  PIN o[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 546.000 303.970 550.000 ;
    END
  END o[71]
  PIN o[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 546.000 308.110 550.000 ;
    END
  END o[72]
  PIN o[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 546.000 312.250 550.000 ;
    END
  END o[73]
  PIN o[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 546.000 316.390 550.000 ;
    END
  END o[74]
  PIN o[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 546.000 320.530 550.000 ;
    END
  END o[75]
  PIN o[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 546.000 324.670 550.000 ;
    END
  END o[76]
  PIN o[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 546.000 328.810 550.000 ;
    END
  END o[77]
  PIN o[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 546.000 332.950 550.000 ;
    END
  END o[78]
  PIN o[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 546.000 337.090 550.000 ;
    END
  END o[79]
  PIN o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 546.000 39.010 550.000 ;
    END
  END o[7]
  PIN o[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 546.000 341.230 550.000 ;
    END
  END o[80]
  PIN o[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 546.000 345.370 550.000 ;
    END
  END o[81]
  PIN o[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 546.000 349.510 550.000 ;
    END
  END o[82]
  PIN o[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 546.000 353.650 550.000 ;
    END
  END o[83]
  PIN o[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 546.000 357.790 550.000 ;
    END
  END o[84]
  PIN o[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 546.000 361.930 550.000 ;
    END
  END o[85]
  PIN o[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 546.000 366.070 550.000 ;
    END
  END o[86]
  PIN o[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 546.000 370.210 550.000 ;
    END
  END o[87]
  PIN o[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 546.000 374.350 550.000 ;
    END
  END o[88]
  PIN o[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 546.000 378.490 550.000 ;
    END
  END o[89]
  PIN o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 546.000 43.150 550.000 ;
    END
  END o[8]
  PIN o[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 546.000 382.630 550.000 ;
    END
  END o[90]
  PIN o[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 546.000 386.770 550.000 ;
    END
  END o[91]
  PIN o[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 546.000 390.910 550.000 ;
    END
  END o[92]
  PIN o[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 546.000 395.050 550.000 ;
    END
  END o[93]
  PIN o[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 546.000 399.190 550.000 ;
    END
  END o[94]
  PIN o[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 546.000 403.330 550.000 ;
    END
  END o[95]
  PIN o[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 546.000 407.470 550.000 ;
    END
  END o[96]
  PIN o[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 546.000 411.610 550.000 ;
    END
  END o[97]
  PIN o[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 546.000 415.750 550.000 ;
    END
  END o[98]
  PIN o[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 546.000 419.890 550.000 ;
    END
  END o[99]
  PIN o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 546.000 47.290 550.000 ;
    END
  END o[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 546.000 539.950 550.000 ;
    END
  END rst
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 544.180 538.645 ;
      LAYER met1 ;
        RECT 0.990 9.220 550.000 538.800 ;
      LAYER met2 ;
        RECT 0.620 545.720 9.470 546.450 ;
        RECT 10.310 545.720 13.610 546.450 ;
        RECT 14.450 545.720 17.750 546.450 ;
        RECT 18.590 545.720 21.890 546.450 ;
        RECT 22.730 545.720 26.030 546.450 ;
        RECT 26.870 545.720 30.170 546.450 ;
        RECT 31.010 545.720 34.310 546.450 ;
        RECT 35.150 545.720 38.450 546.450 ;
        RECT 39.290 545.720 42.590 546.450 ;
        RECT 43.430 545.720 46.730 546.450 ;
        RECT 47.570 545.720 50.870 546.450 ;
        RECT 51.710 545.720 55.010 546.450 ;
        RECT 55.850 545.720 59.150 546.450 ;
        RECT 59.990 545.720 63.290 546.450 ;
        RECT 64.130 545.720 67.430 546.450 ;
        RECT 68.270 545.720 71.570 546.450 ;
        RECT 72.410 545.720 75.710 546.450 ;
        RECT 76.550 545.720 79.850 546.450 ;
        RECT 80.690 545.720 83.990 546.450 ;
        RECT 84.830 545.720 88.130 546.450 ;
        RECT 88.970 545.720 92.270 546.450 ;
        RECT 93.110 545.720 96.410 546.450 ;
        RECT 97.250 545.720 100.550 546.450 ;
        RECT 101.390 545.720 104.690 546.450 ;
        RECT 105.530 545.720 108.830 546.450 ;
        RECT 109.670 545.720 112.970 546.450 ;
        RECT 113.810 545.720 117.110 546.450 ;
        RECT 117.950 545.720 121.250 546.450 ;
        RECT 122.090 545.720 125.390 546.450 ;
        RECT 126.230 545.720 129.530 546.450 ;
        RECT 130.370 545.720 133.670 546.450 ;
        RECT 134.510 545.720 137.810 546.450 ;
        RECT 138.650 545.720 141.950 546.450 ;
        RECT 142.790 545.720 146.090 546.450 ;
        RECT 146.930 545.720 150.230 546.450 ;
        RECT 151.070 545.720 154.370 546.450 ;
        RECT 155.210 545.720 158.510 546.450 ;
        RECT 159.350 545.720 162.650 546.450 ;
        RECT 163.490 545.720 166.790 546.450 ;
        RECT 167.630 545.720 170.930 546.450 ;
        RECT 171.770 545.720 175.070 546.450 ;
        RECT 175.910 545.720 179.210 546.450 ;
        RECT 180.050 545.720 183.350 546.450 ;
        RECT 184.190 545.720 187.490 546.450 ;
        RECT 188.330 545.720 191.630 546.450 ;
        RECT 192.470 545.720 195.770 546.450 ;
        RECT 196.610 545.720 199.910 546.450 ;
        RECT 200.750 545.720 204.050 546.450 ;
        RECT 204.890 545.720 208.190 546.450 ;
        RECT 209.030 545.720 212.330 546.450 ;
        RECT 213.170 545.720 216.470 546.450 ;
        RECT 217.310 545.720 220.610 546.450 ;
        RECT 221.450 545.720 224.750 546.450 ;
        RECT 225.590 545.720 228.890 546.450 ;
        RECT 229.730 545.720 233.030 546.450 ;
        RECT 233.870 545.720 237.170 546.450 ;
        RECT 238.010 545.720 241.310 546.450 ;
        RECT 242.150 545.720 245.450 546.450 ;
        RECT 246.290 545.720 249.590 546.450 ;
        RECT 250.430 545.720 253.730 546.450 ;
        RECT 254.570 545.720 257.870 546.450 ;
        RECT 258.710 545.720 262.010 546.450 ;
        RECT 262.850 545.720 266.150 546.450 ;
        RECT 266.990 545.720 270.290 546.450 ;
        RECT 271.130 545.720 274.430 546.450 ;
        RECT 275.270 545.720 278.570 546.450 ;
        RECT 279.410 545.720 282.710 546.450 ;
        RECT 283.550 545.720 286.850 546.450 ;
        RECT 287.690 545.720 290.990 546.450 ;
        RECT 291.830 545.720 295.130 546.450 ;
        RECT 295.970 545.720 299.270 546.450 ;
        RECT 300.110 545.720 303.410 546.450 ;
        RECT 304.250 545.720 307.550 546.450 ;
        RECT 308.390 545.720 311.690 546.450 ;
        RECT 312.530 545.720 315.830 546.450 ;
        RECT 316.670 545.720 319.970 546.450 ;
        RECT 320.810 545.720 324.110 546.450 ;
        RECT 324.950 545.720 328.250 546.450 ;
        RECT 329.090 545.720 332.390 546.450 ;
        RECT 333.230 545.720 336.530 546.450 ;
        RECT 337.370 545.720 340.670 546.450 ;
        RECT 341.510 545.720 344.810 546.450 ;
        RECT 345.650 545.720 348.950 546.450 ;
        RECT 349.790 545.720 353.090 546.450 ;
        RECT 353.930 545.720 357.230 546.450 ;
        RECT 358.070 545.720 361.370 546.450 ;
        RECT 362.210 545.720 365.510 546.450 ;
        RECT 366.350 545.720 369.650 546.450 ;
        RECT 370.490 545.720 373.790 546.450 ;
        RECT 374.630 545.720 377.930 546.450 ;
        RECT 378.770 545.720 382.070 546.450 ;
        RECT 382.910 545.720 386.210 546.450 ;
        RECT 387.050 545.720 390.350 546.450 ;
        RECT 391.190 545.720 394.490 546.450 ;
        RECT 395.330 545.720 398.630 546.450 ;
        RECT 399.470 545.720 402.770 546.450 ;
        RECT 403.610 545.720 406.910 546.450 ;
        RECT 407.750 545.720 411.050 546.450 ;
        RECT 411.890 545.720 415.190 546.450 ;
        RECT 416.030 545.720 419.330 546.450 ;
        RECT 420.170 545.720 423.470 546.450 ;
        RECT 424.310 545.720 427.610 546.450 ;
        RECT 428.450 545.720 431.750 546.450 ;
        RECT 432.590 545.720 435.890 546.450 ;
        RECT 436.730 545.720 440.030 546.450 ;
        RECT 440.870 545.720 444.170 546.450 ;
        RECT 445.010 545.720 448.310 546.450 ;
        RECT 449.150 545.720 452.450 546.450 ;
        RECT 453.290 545.720 456.590 546.450 ;
        RECT 457.430 545.720 460.730 546.450 ;
        RECT 461.570 545.720 464.870 546.450 ;
        RECT 465.710 545.720 469.010 546.450 ;
        RECT 469.850 545.720 473.150 546.450 ;
        RECT 473.990 545.720 477.290 546.450 ;
        RECT 478.130 545.720 481.430 546.450 ;
        RECT 482.270 545.720 485.570 546.450 ;
        RECT 486.410 545.720 489.710 546.450 ;
        RECT 490.550 545.720 493.850 546.450 ;
        RECT 494.690 545.720 497.990 546.450 ;
        RECT 498.830 545.720 502.130 546.450 ;
        RECT 502.970 545.720 506.270 546.450 ;
        RECT 507.110 545.720 510.410 546.450 ;
        RECT 511.250 545.720 514.550 546.450 ;
        RECT 515.390 545.720 518.690 546.450 ;
        RECT 519.530 545.720 522.830 546.450 ;
        RECT 523.670 545.720 526.970 546.450 ;
        RECT 527.810 545.720 531.110 546.450 ;
        RECT 531.950 545.720 535.250 546.450 ;
        RECT 536.090 545.720 539.390 546.450 ;
        RECT 540.230 545.720 550.000 546.450 ;
        RECT 0.620 4.280 550.000 545.720 ;
        RECT 0.620 4.000 11.770 4.280 ;
        RECT 12.610 4.000 15.910 4.280 ;
        RECT 16.750 4.000 20.050 4.280 ;
        RECT 20.890 4.000 24.190 4.280 ;
        RECT 25.030 4.000 28.330 4.280 ;
        RECT 29.170 4.000 32.470 4.280 ;
        RECT 33.310 4.000 36.610 4.280 ;
        RECT 37.450 4.000 40.750 4.280 ;
        RECT 41.590 4.000 44.890 4.280 ;
        RECT 45.730 4.000 49.030 4.280 ;
        RECT 49.870 4.000 53.170 4.280 ;
        RECT 54.010 4.000 57.310 4.280 ;
        RECT 58.150 4.000 61.450 4.280 ;
        RECT 62.290 4.000 65.590 4.280 ;
        RECT 66.430 4.000 69.730 4.280 ;
        RECT 70.570 4.000 73.870 4.280 ;
        RECT 74.710 4.000 78.010 4.280 ;
        RECT 78.850 4.000 82.150 4.280 ;
        RECT 82.990 4.000 86.290 4.280 ;
        RECT 87.130 4.000 90.430 4.280 ;
        RECT 91.270 4.000 94.570 4.280 ;
        RECT 95.410 4.000 98.710 4.280 ;
        RECT 99.550 4.000 102.850 4.280 ;
        RECT 103.690 4.000 106.990 4.280 ;
        RECT 107.830 4.000 111.130 4.280 ;
        RECT 111.970 4.000 115.270 4.280 ;
        RECT 116.110 4.000 119.410 4.280 ;
        RECT 120.250 4.000 123.550 4.280 ;
        RECT 124.390 4.000 127.690 4.280 ;
        RECT 128.530 4.000 131.830 4.280 ;
        RECT 132.670 4.000 135.970 4.280 ;
        RECT 136.810 4.000 140.110 4.280 ;
        RECT 140.950 4.000 144.250 4.280 ;
        RECT 145.090 4.000 148.390 4.280 ;
        RECT 149.230 4.000 152.530 4.280 ;
        RECT 153.370 4.000 156.670 4.280 ;
        RECT 157.510 4.000 160.810 4.280 ;
        RECT 161.650 4.000 164.950 4.280 ;
        RECT 165.790 4.000 169.090 4.280 ;
        RECT 169.930 4.000 173.230 4.280 ;
        RECT 174.070 4.000 177.370 4.280 ;
        RECT 178.210 4.000 181.510 4.280 ;
        RECT 182.350 4.000 185.650 4.280 ;
        RECT 186.490 4.000 189.790 4.280 ;
        RECT 190.630 4.000 193.930 4.280 ;
        RECT 194.770 4.000 198.070 4.280 ;
        RECT 198.910 4.000 202.210 4.280 ;
        RECT 203.050 4.000 206.350 4.280 ;
        RECT 207.190 4.000 210.490 4.280 ;
        RECT 211.330 4.000 214.630 4.280 ;
        RECT 215.470 4.000 218.770 4.280 ;
        RECT 219.610 4.000 222.910 4.280 ;
        RECT 223.750 4.000 227.050 4.280 ;
        RECT 227.890 4.000 231.190 4.280 ;
        RECT 232.030 4.000 235.330 4.280 ;
        RECT 236.170 4.000 239.470 4.280 ;
        RECT 240.310 4.000 243.610 4.280 ;
        RECT 244.450 4.000 247.750 4.280 ;
        RECT 248.590 4.000 251.890 4.280 ;
        RECT 252.730 4.000 256.030 4.280 ;
        RECT 256.870 4.000 260.170 4.280 ;
        RECT 261.010 4.000 264.310 4.280 ;
        RECT 265.150 4.000 268.450 4.280 ;
        RECT 269.290 4.000 272.590 4.280 ;
        RECT 273.430 4.000 276.730 4.280 ;
        RECT 277.570 4.000 280.870 4.280 ;
        RECT 281.710 4.000 285.010 4.280 ;
        RECT 285.850 4.000 289.150 4.280 ;
        RECT 289.990 4.000 293.290 4.280 ;
        RECT 294.130 4.000 297.430 4.280 ;
        RECT 298.270 4.000 301.570 4.280 ;
        RECT 302.410 4.000 305.710 4.280 ;
        RECT 306.550 4.000 309.850 4.280 ;
        RECT 310.690 4.000 313.990 4.280 ;
        RECT 314.830 4.000 318.130 4.280 ;
        RECT 318.970 4.000 322.270 4.280 ;
        RECT 323.110 4.000 326.410 4.280 ;
        RECT 327.250 4.000 330.550 4.280 ;
        RECT 331.390 4.000 334.690 4.280 ;
        RECT 335.530 4.000 338.830 4.280 ;
        RECT 339.670 4.000 342.970 4.280 ;
        RECT 343.810 4.000 347.110 4.280 ;
        RECT 347.950 4.000 351.250 4.280 ;
        RECT 352.090 4.000 355.390 4.280 ;
        RECT 356.230 4.000 359.530 4.280 ;
        RECT 360.370 4.000 363.670 4.280 ;
        RECT 364.510 4.000 367.810 4.280 ;
        RECT 368.650 4.000 371.950 4.280 ;
        RECT 372.790 4.000 376.090 4.280 ;
        RECT 376.930 4.000 380.230 4.280 ;
        RECT 381.070 4.000 384.370 4.280 ;
        RECT 385.210 4.000 388.510 4.280 ;
        RECT 389.350 4.000 392.650 4.280 ;
        RECT 393.490 4.000 396.790 4.280 ;
        RECT 397.630 4.000 400.930 4.280 ;
        RECT 401.770 4.000 405.070 4.280 ;
        RECT 405.910 4.000 409.210 4.280 ;
        RECT 410.050 4.000 413.350 4.280 ;
        RECT 414.190 4.000 417.490 4.280 ;
        RECT 418.330 4.000 421.630 4.280 ;
        RECT 422.470 4.000 425.770 4.280 ;
        RECT 426.610 4.000 429.910 4.280 ;
        RECT 430.750 4.000 434.050 4.280 ;
        RECT 434.890 4.000 438.190 4.280 ;
        RECT 439.030 4.000 442.330 4.280 ;
        RECT 443.170 4.000 446.470 4.280 ;
        RECT 447.310 4.000 450.610 4.280 ;
        RECT 451.450 4.000 454.750 4.280 ;
        RECT 455.590 4.000 458.890 4.280 ;
        RECT 459.730 4.000 463.030 4.280 ;
        RECT 463.870 4.000 467.170 4.280 ;
        RECT 468.010 4.000 471.310 4.280 ;
        RECT 472.150 4.000 475.450 4.280 ;
        RECT 476.290 4.000 479.590 4.280 ;
        RECT 480.430 4.000 483.730 4.280 ;
        RECT 484.570 4.000 487.870 4.280 ;
        RECT 488.710 4.000 492.010 4.280 ;
        RECT 492.850 4.000 496.150 4.280 ;
        RECT 496.990 4.000 500.290 4.280 ;
        RECT 501.130 4.000 504.430 4.280 ;
        RECT 505.270 4.000 508.570 4.280 ;
        RECT 509.410 4.000 512.710 4.280 ;
        RECT 513.550 4.000 516.850 4.280 ;
        RECT 517.690 4.000 520.990 4.280 ;
        RECT 521.830 4.000 525.130 4.280 ;
        RECT 525.970 4.000 529.270 4.280 ;
        RECT 530.110 4.000 533.410 4.280 ;
        RECT 534.250 4.000 537.550 4.280 ;
        RECT 538.390 4.000 550.000 4.280 ;
      LAYER met3 ;
        RECT 1.905 536.880 549.635 538.725 ;
        RECT 1.905 535.480 545.600 536.880 ;
        RECT 1.905 532.800 549.635 535.480 ;
        RECT 1.905 531.400 545.600 532.800 ;
        RECT 1.905 528.720 549.635 531.400 ;
        RECT 1.905 527.320 545.600 528.720 ;
        RECT 1.905 524.640 549.635 527.320 ;
        RECT 1.905 523.240 545.600 524.640 ;
        RECT 1.905 520.560 549.635 523.240 ;
        RECT 1.905 519.160 545.600 520.560 ;
        RECT 1.905 516.480 549.635 519.160 ;
        RECT 1.905 515.080 545.600 516.480 ;
        RECT 1.905 512.400 549.635 515.080 ;
        RECT 1.905 511.000 545.600 512.400 ;
        RECT 1.905 508.320 549.635 511.000 ;
        RECT 1.905 506.920 545.600 508.320 ;
        RECT 1.905 504.240 549.635 506.920 ;
        RECT 1.905 502.840 545.600 504.240 ;
        RECT 1.905 500.160 549.635 502.840 ;
        RECT 1.905 498.760 545.600 500.160 ;
        RECT 1.905 496.080 549.635 498.760 ;
        RECT 1.905 494.680 545.600 496.080 ;
        RECT 1.905 492.000 549.635 494.680 ;
        RECT 1.905 490.600 545.600 492.000 ;
        RECT 1.905 487.920 549.635 490.600 ;
        RECT 1.905 486.520 545.600 487.920 ;
        RECT 1.905 483.840 549.635 486.520 ;
        RECT 1.905 482.440 545.600 483.840 ;
        RECT 1.905 479.760 549.635 482.440 ;
        RECT 1.905 478.360 545.600 479.760 ;
        RECT 1.905 475.680 549.635 478.360 ;
        RECT 1.905 474.280 545.600 475.680 ;
        RECT 1.905 471.600 549.635 474.280 ;
        RECT 1.905 470.200 545.600 471.600 ;
        RECT 1.905 467.520 549.635 470.200 ;
        RECT 1.905 466.120 545.600 467.520 ;
        RECT 1.905 463.440 549.635 466.120 ;
        RECT 1.905 462.040 545.600 463.440 ;
        RECT 1.905 459.360 549.635 462.040 ;
        RECT 1.905 457.960 545.600 459.360 ;
        RECT 1.905 455.280 549.635 457.960 ;
        RECT 1.905 453.880 545.600 455.280 ;
        RECT 1.905 451.200 549.635 453.880 ;
        RECT 1.905 449.800 545.600 451.200 ;
        RECT 1.905 447.120 549.635 449.800 ;
        RECT 1.905 445.720 545.600 447.120 ;
        RECT 1.905 443.040 549.635 445.720 ;
        RECT 1.905 441.640 545.600 443.040 ;
        RECT 1.905 438.960 549.635 441.640 ;
        RECT 1.905 437.560 545.600 438.960 ;
        RECT 1.905 434.880 549.635 437.560 ;
        RECT 1.905 433.480 545.600 434.880 ;
        RECT 1.905 430.800 549.635 433.480 ;
        RECT 1.905 429.400 545.600 430.800 ;
        RECT 1.905 426.720 549.635 429.400 ;
        RECT 1.905 425.320 545.600 426.720 ;
        RECT 1.905 422.640 549.635 425.320 ;
        RECT 1.905 421.240 545.600 422.640 ;
        RECT 1.905 418.560 549.635 421.240 ;
        RECT 1.905 417.160 545.600 418.560 ;
        RECT 1.905 414.480 549.635 417.160 ;
        RECT 1.905 413.080 545.600 414.480 ;
        RECT 1.905 410.400 549.635 413.080 ;
        RECT 1.905 409.000 545.600 410.400 ;
        RECT 1.905 406.320 549.635 409.000 ;
        RECT 1.905 404.920 545.600 406.320 ;
        RECT 1.905 402.240 549.635 404.920 ;
        RECT 1.905 400.840 545.600 402.240 ;
        RECT 1.905 398.160 549.635 400.840 ;
        RECT 1.905 396.760 545.600 398.160 ;
        RECT 1.905 394.080 549.635 396.760 ;
        RECT 1.905 392.680 545.600 394.080 ;
        RECT 1.905 390.000 549.635 392.680 ;
        RECT 1.905 388.600 545.600 390.000 ;
        RECT 1.905 385.920 549.635 388.600 ;
        RECT 1.905 384.520 545.600 385.920 ;
        RECT 1.905 381.840 549.635 384.520 ;
        RECT 1.905 380.440 545.600 381.840 ;
        RECT 1.905 377.760 549.635 380.440 ;
        RECT 1.905 376.360 545.600 377.760 ;
        RECT 1.905 373.680 549.635 376.360 ;
        RECT 1.905 372.280 545.600 373.680 ;
        RECT 1.905 369.600 549.635 372.280 ;
        RECT 1.905 368.200 545.600 369.600 ;
        RECT 1.905 365.520 549.635 368.200 ;
        RECT 1.905 364.120 545.600 365.520 ;
        RECT 1.905 361.440 549.635 364.120 ;
        RECT 1.905 360.040 545.600 361.440 ;
        RECT 1.905 357.360 549.635 360.040 ;
        RECT 1.905 355.960 545.600 357.360 ;
        RECT 1.905 353.280 549.635 355.960 ;
        RECT 1.905 351.880 545.600 353.280 ;
        RECT 1.905 349.200 549.635 351.880 ;
        RECT 1.905 347.800 545.600 349.200 ;
        RECT 1.905 345.120 549.635 347.800 ;
        RECT 1.905 343.720 545.600 345.120 ;
        RECT 1.905 341.040 549.635 343.720 ;
        RECT 1.905 339.640 545.600 341.040 ;
        RECT 1.905 336.960 549.635 339.640 ;
        RECT 1.905 335.560 545.600 336.960 ;
        RECT 1.905 332.880 549.635 335.560 ;
        RECT 1.905 331.480 545.600 332.880 ;
        RECT 1.905 328.800 549.635 331.480 ;
        RECT 1.905 327.400 545.600 328.800 ;
        RECT 1.905 324.720 549.635 327.400 ;
        RECT 1.905 323.320 545.600 324.720 ;
        RECT 1.905 320.640 549.635 323.320 ;
        RECT 1.905 319.240 545.600 320.640 ;
        RECT 1.905 316.560 549.635 319.240 ;
        RECT 1.905 315.160 545.600 316.560 ;
        RECT 1.905 312.480 549.635 315.160 ;
        RECT 1.905 311.080 545.600 312.480 ;
        RECT 1.905 308.400 549.635 311.080 ;
        RECT 1.905 307.000 545.600 308.400 ;
        RECT 1.905 304.320 549.635 307.000 ;
        RECT 1.905 302.920 545.600 304.320 ;
        RECT 1.905 300.240 549.635 302.920 ;
        RECT 1.905 298.840 545.600 300.240 ;
        RECT 1.905 296.160 549.635 298.840 ;
        RECT 1.905 294.760 545.600 296.160 ;
        RECT 1.905 292.080 549.635 294.760 ;
        RECT 1.905 290.680 545.600 292.080 ;
        RECT 1.905 288.000 549.635 290.680 ;
        RECT 1.905 286.600 545.600 288.000 ;
        RECT 1.905 283.920 549.635 286.600 ;
        RECT 1.905 282.520 545.600 283.920 ;
        RECT 1.905 279.840 549.635 282.520 ;
        RECT 1.905 278.440 545.600 279.840 ;
        RECT 1.905 275.760 549.635 278.440 ;
        RECT 1.905 274.360 545.600 275.760 ;
        RECT 1.905 271.680 549.635 274.360 ;
        RECT 1.905 270.280 545.600 271.680 ;
        RECT 1.905 267.600 549.635 270.280 ;
        RECT 1.905 266.200 545.600 267.600 ;
        RECT 1.905 263.520 549.635 266.200 ;
        RECT 1.905 262.120 545.600 263.520 ;
        RECT 1.905 259.440 549.635 262.120 ;
        RECT 1.905 258.040 545.600 259.440 ;
        RECT 1.905 255.360 549.635 258.040 ;
        RECT 1.905 253.960 545.600 255.360 ;
        RECT 1.905 251.280 549.635 253.960 ;
        RECT 1.905 249.880 545.600 251.280 ;
        RECT 1.905 247.200 549.635 249.880 ;
        RECT 1.905 245.800 545.600 247.200 ;
        RECT 1.905 243.120 549.635 245.800 ;
        RECT 1.905 241.720 545.600 243.120 ;
        RECT 1.905 239.040 549.635 241.720 ;
        RECT 1.905 237.640 545.600 239.040 ;
        RECT 1.905 234.960 549.635 237.640 ;
        RECT 1.905 233.560 545.600 234.960 ;
        RECT 1.905 230.880 549.635 233.560 ;
        RECT 1.905 229.480 545.600 230.880 ;
        RECT 1.905 226.800 549.635 229.480 ;
        RECT 1.905 225.400 545.600 226.800 ;
        RECT 1.905 222.720 549.635 225.400 ;
        RECT 1.905 221.320 545.600 222.720 ;
        RECT 1.905 218.640 549.635 221.320 ;
        RECT 1.905 217.240 545.600 218.640 ;
        RECT 1.905 214.560 549.635 217.240 ;
        RECT 1.905 213.160 545.600 214.560 ;
        RECT 1.905 210.480 549.635 213.160 ;
        RECT 1.905 209.080 545.600 210.480 ;
        RECT 1.905 206.400 549.635 209.080 ;
        RECT 1.905 205.000 545.600 206.400 ;
        RECT 1.905 202.320 549.635 205.000 ;
        RECT 1.905 200.920 545.600 202.320 ;
        RECT 1.905 198.240 549.635 200.920 ;
        RECT 1.905 196.840 545.600 198.240 ;
        RECT 1.905 194.160 549.635 196.840 ;
        RECT 1.905 192.760 545.600 194.160 ;
        RECT 1.905 190.080 549.635 192.760 ;
        RECT 1.905 188.680 545.600 190.080 ;
        RECT 1.905 186.000 549.635 188.680 ;
        RECT 1.905 184.600 545.600 186.000 ;
        RECT 1.905 181.920 549.635 184.600 ;
        RECT 1.905 180.520 545.600 181.920 ;
        RECT 1.905 177.840 549.635 180.520 ;
        RECT 1.905 176.440 545.600 177.840 ;
        RECT 1.905 173.760 549.635 176.440 ;
        RECT 1.905 172.360 545.600 173.760 ;
        RECT 1.905 169.680 549.635 172.360 ;
        RECT 1.905 168.280 545.600 169.680 ;
        RECT 1.905 165.600 549.635 168.280 ;
        RECT 1.905 164.200 545.600 165.600 ;
        RECT 1.905 161.520 549.635 164.200 ;
        RECT 1.905 160.120 545.600 161.520 ;
        RECT 1.905 157.440 549.635 160.120 ;
        RECT 1.905 156.040 545.600 157.440 ;
        RECT 1.905 153.360 549.635 156.040 ;
        RECT 1.905 151.960 545.600 153.360 ;
        RECT 1.905 149.280 549.635 151.960 ;
        RECT 1.905 147.880 545.600 149.280 ;
        RECT 1.905 145.200 549.635 147.880 ;
        RECT 1.905 143.800 545.600 145.200 ;
        RECT 1.905 141.120 549.635 143.800 ;
        RECT 1.905 139.720 545.600 141.120 ;
        RECT 1.905 137.040 549.635 139.720 ;
        RECT 1.905 135.640 545.600 137.040 ;
        RECT 1.905 132.960 549.635 135.640 ;
        RECT 1.905 131.560 545.600 132.960 ;
        RECT 1.905 128.880 549.635 131.560 ;
        RECT 1.905 127.480 545.600 128.880 ;
        RECT 1.905 124.800 549.635 127.480 ;
        RECT 1.905 123.400 545.600 124.800 ;
        RECT 1.905 120.720 549.635 123.400 ;
        RECT 1.905 119.320 545.600 120.720 ;
        RECT 1.905 116.640 549.635 119.320 ;
        RECT 1.905 115.240 545.600 116.640 ;
        RECT 1.905 112.560 549.635 115.240 ;
        RECT 1.905 111.160 545.600 112.560 ;
        RECT 1.905 108.480 549.635 111.160 ;
        RECT 1.905 107.080 545.600 108.480 ;
        RECT 1.905 104.400 549.635 107.080 ;
        RECT 1.905 103.000 545.600 104.400 ;
        RECT 1.905 100.320 549.635 103.000 ;
        RECT 1.905 98.920 545.600 100.320 ;
        RECT 1.905 96.240 549.635 98.920 ;
        RECT 1.905 94.840 545.600 96.240 ;
        RECT 1.905 92.160 549.635 94.840 ;
        RECT 1.905 90.760 545.600 92.160 ;
        RECT 1.905 88.080 549.635 90.760 ;
        RECT 1.905 86.680 545.600 88.080 ;
        RECT 1.905 84.000 549.635 86.680 ;
        RECT 1.905 82.600 545.600 84.000 ;
        RECT 1.905 79.920 549.635 82.600 ;
        RECT 1.905 78.520 545.600 79.920 ;
        RECT 1.905 75.840 549.635 78.520 ;
        RECT 1.905 74.440 545.600 75.840 ;
        RECT 1.905 71.760 549.635 74.440 ;
        RECT 1.905 70.360 545.600 71.760 ;
        RECT 1.905 67.680 549.635 70.360 ;
        RECT 1.905 66.280 545.600 67.680 ;
        RECT 1.905 63.600 549.635 66.280 ;
        RECT 1.905 62.200 545.600 63.600 ;
        RECT 1.905 59.520 549.635 62.200 ;
        RECT 1.905 58.120 545.600 59.520 ;
        RECT 1.905 55.440 549.635 58.120 ;
        RECT 1.905 54.040 545.600 55.440 ;
        RECT 1.905 51.360 549.635 54.040 ;
        RECT 1.905 49.960 545.600 51.360 ;
        RECT 1.905 47.280 549.635 49.960 ;
        RECT 1.905 45.880 545.600 47.280 ;
        RECT 1.905 43.200 549.635 45.880 ;
        RECT 1.905 41.800 545.600 43.200 ;
        RECT 1.905 39.120 549.635 41.800 ;
        RECT 1.905 37.720 545.600 39.120 ;
        RECT 1.905 35.040 549.635 37.720 ;
        RECT 1.905 33.640 545.600 35.040 ;
        RECT 1.905 30.960 549.635 33.640 ;
        RECT 1.905 29.560 545.600 30.960 ;
        RECT 1.905 26.880 549.635 29.560 ;
        RECT 1.905 25.480 545.600 26.880 ;
        RECT 1.905 22.800 549.635 25.480 ;
        RECT 1.905 21.400 545.600 22.800 ;
        RECT 1.905 18.720 549.635 21.400 ;
        RECT 1.905 17.320 545.600 18.720 ;
        RECT 1.905 14.640 549.635 17.320 ;
        RECT 1.905 13.240 545.600 14.640 ;
        RECT 1.905 10.715 549.635 13.240 ;
      LAYER met4 ;
        RECT 2.135 13.095 8.570 536.345 ;
        RECT 12.470 13.095 98.570 536.345 ;
        RECT 102.470 13.095 188.570 536.345 ;
        RECT 192.470 13.095 278.570 536.345 ;
        RECT 282.470 13.095 368.570 536.345 ;
        RECT 372.470 13.095 458.570 536.345 ;
        RECT 462.470 13.095 547.105 536.345 ;
  END
END multiply_add_64x64
END LIBRARY

