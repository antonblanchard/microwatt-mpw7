magic
tech sky130A
magscale 1 2
timestamp 1657540616
<< obsli1 >>
rect 1104 2159 228896 227409
<< obsm1 >>
rect 566 484 228896 227440
<< metal2 >>
rect 4250 229200 4306 230000
rect 11886 229200 11942 230000
rect 19522 229200 19578 230000
rect 27158 229200 27214 230000
rect 34794 229200 34850 230000
rect 42430 229200 42486 230000
rect 50066 229200 50122 230000
rect 57702 229200 57758 230000
rect 65338 229200 65394 230000
rect 72974 229200 73030 230000
rect 80610 229200 80666 230000
rect 88246 229200 88302 230000
rect 95882 229200 95938 230000
rect 103518 229200 103574 230000
rect 111154 229200 111210 230000
rect 118790 229200 118846 230000
rect 126426 229200 126482 230000
rect 134062 229200 134118 230000
rect 141698 229200 141754 230000
rect 149334 229200 149390 230000
rect 156970 229200 157026 230000
rect 164606 229200 164662 230000
rect 172242 229200 172298 230000
rect 179878 229200 179934 230000
rect 187514 229200 187570 230000
rect 195150 229200 195206 230000
rect 202786 229200 202842 230000
rect 210422 229200 210478 230000
rect 218058 229200 218114 230000
rect 225694 229200 225750 230000
rect 3974 0 4030 800
rect 5722 0 5778 800
rect 7470 0 7526 800
rect 9218 0 9274 800
rect 10966 0 11022 800
rect 12714 0 12770 800
rect 14462 0 14518 800
rect 16210 0 16266 800
rect 17958 0 18014 800
rect 19706 0 19762 800
rect 21454 0 21510 800
rect 23202 0 23258 800
rect 24950 0 25006 800
rect 26698 0 26754 800
rect 28446 0 28502 800
rect 30194 0 30250 800
rect 31942 0 31998 800
rect 33690 0 33746 800
rect 35438 0 35494 800
rect 37186 0 37242 800
rect 38934 0 38990 800
rect 40682 0 40738 800
rect 42430 0 42486 800
rect 44178 0 44234 800
rect 45926 0 45982 800
rect 47674 0 47730 800
rect 49422 0 49478 800
rect 51170 0 51226 800
rect 52918 0 52974 800
rect 54666 0 54722 800
rect 56414 0 56470 800
rect 58162 0 58218 800
rect 59910 0 59966 800
rect 61658 0 61714 800
rect 63406 0 63462 800
rect 65154 0 65210 800
rect 66902 0 66958 800
rect 68650 0 68706 800
rect 70398 0 70454 800
rect 72146 0 72202 800
rect 73894 0 73950 800
rect 75642 0 75698 800
rect 77390 0 77446 800
rect 79138 0 79194 800
rect 80886 0 80942 800
rect 82634 0 82690 800
rect 84382 0 84438 800
rect 86130 0 86186 800
rect 87878 0 87934 800
rect 89626 0 89682 800
rect 91374 0 91430 800
rect 93122 0 93178 800
rect 94870 0 94926 800
rect 96618 0 96674 800
rect 98366 0 98422 800
rect 100114 0 100170 800
rect 101862 0 101918 800
rect 103610 0 103666 800
rect 105358 0 105414 800
rect 107106 0 107162 800
rect 108854 0 108910 800
rect 110602 0 110658 800
rect 112350 0 112406 800
rect 114098 0 114154 800
rect 115846 0 115902 800
rect 117594 0 117650 800
rect 119342 0 119398 800
rect 121090 0 121146 800
rect 122838 0 122894 800
rect 124586 0 124642 800
rect 126334 0 126390 800
rect 128082 0 128138 800
rect 129830 0 129886 800
rect 131578 0 131634 800
rect 133326 0 133382 800
rect 135074 0 135130 800
rect 136822 0 136878 800
rect 138570 0 138626 800
rect 140318 0 140374 800
rect 142066 0 142122 800
rect 143814 0 143870 800
rect 145562 0 145618 800
rect 147310 0 147366 800
rect 149058 0 149114 800
rect 150806 0 150862 800
rect 152554 0 152610 800
rect 154302 0 154358 800
rect 156050 0 156106 800
rect 157798 0 157854 800
rect 159546 0 159602 800
rect 161294 0 161350 800
rect 163042 0 163098 800
rect 164790 0 164846 800
rect 166538 0 166594 800
rect 168286 0 168342 800
rect 170034 0 170090 800
rect 171782 0 171838 800
rect 173530 0 173586 800
rect 175278 0 175334 800
rect 177026 0 177082 800
rect 178774 0 178830 800
rect 180522 0 180578 800
rect 182270 0 182326 800
rect 184018 0 184074 800
rect 185766 0 185822 800
rect 187514 0 187570 800
rect 189262 0 189318 800
rect 191010 0 191066 800
rect 192758 0 192814 800
rect 194506 0 194562 800
rect 196254 0 196310 800
rect 198002 0 198058 800
rect 199750 0 199806 800
rect 201498 0 201554 800
rect 203246 0 203302 800
rect 204994 0 205050 800
rect 206742 0 206798 800
rect 208490 0 208546 800
rect 210238 0 210294 800
rect 211986 0 212042 800
rect 213734 0 213790 800
rect 215482 0 215538 800
rect 217230 0 217286 800
rect 218978 0 219034 800
rect 220726 0 220782 800
rect 222474 0 222530 800
rect 224222 0 224278 800
rect 225970 0 226026 800
<< obsm2 >>
rect 572 229144 4194 229200
rect 4362 229144 11830 229200
rect 11998 229144 19466 229200
rect 19634 229144 27102 229200
rect 27270 229144 34738 229200
rect 34906 229144 42374 229200
rect 42542 229144 50010 229200
rect 50178 229144 57646 229200
rect 57814 229144 65282 229200
rect 65450 229144 72918 229200
rect 73086 229144 80554 229200
rect 80722 229144 88190 229200
rect 88358 229144 95826 229200
rect 95994 229144 103462 229200
rect 103630 229144 111098 229200
rect 111266 229144 118734 229200
rect 118902 229144 126370 229200
rect 126538 229144 134006 229200
rect 134174 229144 141642 229200
rect 141810 229144 149278 229200
rect 149446 229144 156914 229200
rect 157082 229144 164550 229200
rect 164718 229144 172186 229200
rect 172354 229144 179822 229200
rect 179990 229144 187458 229200
rect 187626 229144 195094 229200
rect 195262 229144 202730 229200
rect 202898 229144 210366 229200
rect 210534 229144 218002 229200
rect 218170 229144 225638 229200
rect 225806 229144 228232 229200
rect 572 856 228232 229144
rect 572 478 3918 856
rect 4086 478 5666 856
rect 5834 478 7414 856
rect 7582 478 9162 856
rect 9330 478 10910 856
rect 11078 478 12658 856
rect 12826 478 14406 856
rect 14574 478 16154 856
rect 16322 478 17902 856
rect 18070 478 19650 856
rect 19818 478 21398 856
rect 21566 478 23146 856
rect 23314 478 24894 856
rect 25062 478 26642 856
rect 26810 478 28390 856
rect 28558 478 30138 856
rect 30306 478 31886 856
rect 32054 478 33634 856
rect 33802 478 35382 856
rect 35550 478 37130 856
rect 37298 478 38878 856
rect 39046 478 40626 856
rect 40794 478 42374 856
rect 42542 478 44122 856
rect 44290 478 45870 856
rect 46038 478 47618 856
rect 47786 478 49366 856
rect 49534 478 51114 856
rect 51282 478 52862 856
rect 53030 478 54610 856
rect 54778 478 56358 856
rect 56526 478 58106 856
rect 58274 478 59854 856
rect 60022 478 61602 856
rect 61770 478 63350 856
rect 63518 478 65098 856
rect 65266 478 66846 856
rect 67014 478 68594 856
rect 68762 478 70342 856
rect 70510 478 72090 856
rect 72258 478 73838 856
rect 74006 478 75586 856
rect 75754 478 77334 856
rect 77502 478 79082 856
rect 79250 478 80830 856
rect 80998 478 82578 856
rect 82746 478 84326 856
rect 84494 478 86074 856
rect 86242 478 87822 856
rect 87990 478 89570 856
rect 89738 478 91318 856
rect 91486 478 93066 856
rect 93234 478 94814 856
rect 94982 478 96562 856
rect 96730 478 98310 856
rect 98478 478 100058 856
rect 100226 478 101806 856
rect 101974 478 103554 856
rect 103722 478 105302 856
rect 105470 478 107050 856
rect 107218 478 108798 856
rect 108966 478 110546 856
rect 110714 478 112294 856
rect 112462 478 114042 856
rect 114210 478 115790 856
rect 115958 478 117538 856
rect 117706 478 119286 856
rect 119454 478 121034 856
rect 121202 478 122782 856
rect 122950 478 124530 856
rect 124698 478 126278 856
rect 126446 478 128026 856
rect 128194 478 129774 856
rect 129942 478 131522 856
rect 131690 478 133270 856
rect 133438 478 135018 856
rect 135186 478 136766 856
rect 136934 478 138514 856
rect 138682 478 140262 856
rect 140430 478 142010 856
rect 142178 478 143758 856
rect 143926 478 145506 856
rect 145674 478 147254 856
rect 147422 478 149002 856
rect 149170 478 150750 856
rect 150918 478 152498 856
rect 152666 478 154246 856
rect 154414 478 155994 856
rect 156162 478 157742 856
rect 157910 478 159490 856
rect 159658 478 161238 856
rect 161406 478 162986 856
rect 163154 478 164734 856
rect 164902 478 166482 856
rect 166650 478 168230 856
rect 168398 478 169978 856
rect 170146 478 171726 856
rect 171894 478 173474 856
rect 173642 478 175222 856
rect 175390 478 176970 856
rect 177138 478 178718 856
rect 178886 478 180466 856
rect 180634 478 182214 856
rect 182382 478 183962 856
rect 184130 478 185710 856
rect 185878 478 187458 856
rect 187626 478 189206 856
rect 189374 478 190954 856
rect 191122 478 192702 856
rect 192870 478 194450 856
rect 194618 478 196198 856
rect 196366 478 197946 856
rect 198114 478 199694 856
rect 199862 478 201442 856
rect 201610 478 203190 856
rect 203358 478 204938 856
rect 205106 478 206686 856
rect 206854 478 208434 856
rect 208602 478 210182 856
rect 210350 478 211930 856
rect 212098 478 213678 856
rect 213846 478 215426 856
rect 215594 478 217174 856
rect 217342 478 218922 856
rect 219090 478 220670 856
rect 220838 478 222418 856
rect 222586 478 224166 856
rect 224334 478 225914 856
rect 226082 478 228232 856
<< metal3 >>
rect 0 227128 800 227248
rect 0 225360 800 225480
rect 0 223592 800 223712
rect 0 221824 800 221944
rect 0 220056 800 220176
rect 0 218288 800 218408
rect 0 216520 800 216640
rect 0 214752 800 214872
rect 0 212984 800 213104
rect 0 211216 800 211336
rect 0 209448 800 209568
rect 0 207680 800 207800
rect 0 205912 800 206032
rect 0 204144 800 204264
rect 0 202376 800 202496
rect 0 200608 800 200728
rect 0 198840 800 198960
rect 0 197072 800 197192
rect 0 195304 800 195424
rect 0 193536 800 193656
rect 0 191768 800 191888
rect 0 190000 800 190120
rect 0 188232 800 188352
rect 0 186464 800 186584
rect 0 184696 800 184816
rect 0 182928 800 183048
rect 0 181160 800 181280
rect 0 179392 800 179512
rect 0 177624 800 177744
rect 0 175856 800 175976
rect 0 174088 800 174208
rect 0 172320 800 172440
rect 0 170552 800 170672
rect 0 168784 800 168904
rect 0 167016 800 167136
rect 0 165248 800 165368
rect 0 163480 800 163600
rect 0 161712 800 161832
rect 0 159944 800 160064
rect 0 158176 800 158296
rect 0 156408 800 156528
rect 0 154640 800 154760
rect 0 152872 800 152992
rect 0 151104 800 151224
rect 0 149336 800 149456
rect 0 147568 800 147688
rect 0 145800 800 145920
rect 0 144032 800 144152
rect 0 142264 800 142384
rect 0 140496 800 140616
rect 0 138728 800 138848
rect 0 136960 800 137080
rect 0 135192 800 135312
rect 0 133424 800 133544
rect 0 131656 800 131776
rect 0 129888 800 130008
rect 0 128120 800 128240
rect 0 126352 800 126472
rect 0 124584 800 124704
rect 0 122816 800 122936
rect 0 121048 800 121168
rect 0 119280 800 119400
rect 0 117512 800 117632
rect 0 115744 800 115864
rect 0 113976 800 114096
rect 0 112208 800 112328
rect 0 110440 800 110560
rect 0 108672 800 108792
rect 0 106904 800 107024
rect 0 105136 800 105256
rect 0 103368 800 103488
rect 0 101600 800 101720
rect 0 99832 800 99952
rect 0 98064 800 98184
rect 0 96296 800 96416
rect 0 94528 800 94648
rect 0 92760 800 92880
rect 0 90992 800 91112
rect 0 89224 800 89344
rect 0 87456 800 87576
rect 0 85688 800 85808
rect 0 83920 800 84040
rect 0 82152 800 82272
rect 0 80384 800 80504
rect 0 78616 800 78736
rect 0 76848 800 76968
rect 0 75080 800 75200
rect 0 73312 800 73432
rect 0 71544 800 71664
rect 0 69776 800 69896
rect 0 68008 800 68128
rect 0 66240 800 66360
rect 0 64472 800 64592
rect 0 62704 800 62824
rect 0 60936 800 61056
rect 0 59168 800 59288
rect 0 57400 800 57520
rect 0 55632 800 55752
rect 0 53864 800 53984
rect 0 52096 800 52216
rect 0 50328 800 50448
rect 0 48560 800 48680
rect 0 46792 800 46912
rect 0 45024 800 45144
rect 0 43256 800 43376
rect 0 41488 800 41608
rect 0 39720 800 39840
rect 0 37952 800 38072
rect 0 36184 800 36304
rect 0 34416 800 34536
rect 0 32648 800 32768
rect 0 30880 800 31000
rect 0 29112 800 29232
rect 0 27344 800 27464
rect 0 25576 800 25696
rect 0 23808 800 23928
rect 0 22040 800 22160
rect 0 20272 800 20392
rect 0 18504 800 18624
rect 0 16736 800 16856
rect 0 14968 800 15088
rect 0 13200 800 13320
rect 0 11432 800 11552
rect 0 9664 800 9784
rect 0 7896 800 8016
rect 0 6128 800 6248
rect 0 4360 800 4480
rect 0 2592 800 2712
<< obsm3 >>
rect 749 227328 227319 227425
rect 880 227048 227319 227328
rect 749 225560 227319 227048
rect 880 225280 227319 225560
rect 749 223792 227319 225280
rect 880 223512 227319 223792
rect 749 222024 227319 223512
rect 880 221744 227319 222024
rect 749 220256 227319 221744
rect 880 219976 227319 220256
rect 749 218488 227319 219976
rect 880 218208 227319 218488
rect 749 216720 227319 218208
rect 880 216440 227319 216720
rect 749 214952 227319 216440
rect 880 214672 227319 214952
rect 749 213184 227319 214672
rect 880 212904 227319 213184
rect 749 211416 227319 212904
rect 880 211136 227319 211416
rect 749 209648 227319 211136
rect 880 209368 227319 209648
rect 749 207880 227319 209368
rect 880 207600 227319 207880
rect 749 206112 227319 207600
rect 880 205832 227319 206112
rect 749 204344 227319 205832
rect 880 204064 227319 204344
rect 749 202576 227319 204064
rect 880 202296 227319 202576
rect 749 200808 227319 202296
rect 880 200528 227319 200808
rect 749 199040 227319 200528
rect 880 198760 227319 199040
rect 749 197272 227319 198760
rect 880 196992 227319 197272
rect 749 195504 227319 196992
rect 880 195224 227319 195504
rect 749 193736 227319 195224
rect 880 193456 227319 193736
rect 749 191968 227319 193456
rect 880 191688 227319 191968
rect 749 190200 227319 191688
rect 880 189920 227319 190200
rect 749 188432 227319 189920
rect 880 188152 227319 188432
rect 749 186664 227319 188152
rect 880 186384 227319 186664
rect 749 184896 227319 186384
rect 880 184616 227319 184896
rect 749 183128 227319 184616
rect 880 182848 227319 183128
rect 749 181360 227319 182848
rect 880 181080 227319 181360
rect 749 179592 227319 181080
rect 880 179312 227319 179592
rect 749 177824 227319 179312
rect 880 177544 227319 177824
rect 749 176056 227319 177544
rect 880 175776 227319 176056
rect 749 174288 227319 175776
rect 880 174008 227319 174288
rect 749 172520 227319 174008
rect 880 172240 227319 172520
rect 749 170752 227319 172240
rect 880 170472 227319 170752
rect 749 168984 227319 170472
rect 880 168704 227319 168984
rect 749 167216 227319 168704
rect 880 166936 227319 167216
rect 749 165448 227319 166936
rect 880 165168 227319 165448
rect 749 163680 227319 165168
rect 880 163400 227319 163680
rect 749 161912 227319 163400
rect 880 161632 227319 161912
rect 749 160144 227319 161632
rect 880 159864 227319 160144
rect 749 158376 227319 159864
rect 880 158096 227319 158376
rect 749 156608 227319 158096
rect 880 156328 227319 156608
rect 749 154840 227319 156328
rect 880 154560 227319 154840
rect 749 153072 227319 154560
rect 880 152792 227319 153072
rect 749 151304 227319 152792
rect 880 151024 227319 151304
rect 749 149536 227319 151024
rect 880 149256 227319 149536
rect 749 147768 227319 149256
rect 880 147488 227319 147768
rect 749 146000 227319 147488
rect 880 145720 227319 146000
rect 749 144232 227319 145720
rect 880 143952 227319 144232
rect 749 142464 227319 143952
rect 880 142184 227319 142464
rect 749 140696 227319 142184
rect 880 140416 227319 140696
rect 749 138928 227319 140416
rect 880 138648 227319 138928
rect 749 137160 227319 138648
rect 880 136880 227319 137160
rect 749 135392 227319 136880
rect 880 135112 227319 135392
rect 749 133624 227319 135112
rect 880 133344 227319 133624
rect 749 131856 227319 133344
rect 880 131576 227319 131856
rect 749 130088 227319 131576
rect 880 129808 227319 130088
rect 749 128320 227319 129808
rect 880 128040 227319 128320
rect 749 126552 227319 128040
rect 880 126272 227319 126552
rect 749 124784 227319 126272
rect 880 124504 227319 124784
rect 749 123016 227319 124504
rect 880 122736 227319 123016
rect 749 121248 227319 122736
rect 880 120968 227319 121248
rect 749 119480 227319 120968
rect 880 119200 227319 119480
rect 749 117712 227319 119200
rect 880 117432 227319 117712
rect 749 115944 227319 117432
rect 880 115664 227319 115944
rect 749 114176 227319 115664
rect 880 113896 227319 114176
rect 749 112408 227319 113896
rect 880 112128 227319 112408
rect 749 110640 227319 112128
rect 880 110360 227319 110640
rect 749 108872 227319 110360
rect 880 108592 227319 108872
rect 749 107104 227319 108592
rect 880 106824 227319 107104
rect 749 105336 227319 106824
rect 880 105056 227319 105336
rect 749 103568 227319 105056
rect 880 103288 227319 103568
rect 749 101800 227319 103288
rect 880 101520 227319 101800
rect 749 100032 227319 101520
rect 880 99752 227319 100032
rect 749 98264 227319 99752
rect 880 97984 227319 98264
rect 749 96496 227319 97984
rect 880 96216 227319 96496
rect 749 94728 227319 96216
rect 880 94448 227319 94728
rect 749 92960 227319 94448
rect 880 92680 227319 92960
rect 749 91192 227319 92680
rect 880 90912 227319 91192
rect 749 89424 227319 90912
rect 880 89144 227319 89424
rect 749 87656 227319 89144
rect 880 87376 227319 87656
rect 749 85888 227319 87376
rect 880 85608 227319 85888
rect 749 84120 227319 85608
rect 880 83840 227319 84120
rect 749 82352 227319 83840
rect 880 82072 227319 82352
rect 749 80584 227319 82072
rect 880 80304 227319 80584
rect 749 78816 227319 80304
rect 880 78536 227319 78816
rect 749 77048 227319 78536
rect 880 76768 227319 77048
rect 749 75280 227319 76768
rect 880 75000 227319 75280
rect 749 73512 227319 75000
rect 880 73232 227319 73512
rect 749 71744 227319 73232
rect 880 71464 227319 71744
rect 749 69976 227319 71464
rect 880 69696 227319 69976
rect 749 68208 227319 69696
rect 880 67928 227319 68208
rect 749 66440 227319 67928
rect 880 66160 227319 66440
rect 749 64672 227319 66160
rect 880 64392 227319 64672
rect 749 62904 227319 64392
rect 880 62624 227319 62904
rect 749 61136 227319 62624
rect 880 60856 227319 61136
rect 749 59368 227319 60856
rect 880 59088 227319 59368
rect 749 57600 227319 59088
rect 880 57320 227319 57600
rect 749 55832 227319 57320
rect 880 55552 227319 55832
rect 749 54064 227319 55552
rect 880 53784 227319 54064
rect 749 52296 227319 53784
rect 880 52016 227319 52296
rect 749 50528 227319 52016
rect 880 50248 227319 50528
rect 749 48760 227319 50248
rect 880 48480 227319 48760
rect 749 46992 227319 48480
rect 880 46712 227319 46992
rect 749 45224 227319 46712
rect 880 44944 227319 45224
rect 749 43456 227319 44944
rect 880 43176 227319 43456
rect 749 41688 227319 43176
rect 880 41408 227319 41688
rect 749 39920 227319 41408
rect 880 39640 227319 39920
rect 749 38152 227319 39640
rect 880 37872 227319 38152
rect 749 36384 227319 37872
rect 880 36104 227319 36384
rect 749 34616 227319 36104
rect 880 34336 227319 34616
rect 749 32848 227319 34336
rect 880 32568 227319 32848
rect 749 31080 227319 32568
rect 880 30800 227319 31080
rect 749 29312 227319 30800
rect 880 29032 227319 29312
rect 749 27544 227319 29032
rect 880 27264 227319 27544
rect 749 25776 227319 27264
rect 880 25496 227319 25776
rect 749 24008 227319 25496
rect 880 23728 227319 24008
rect 749 22240 227319 23728
rect 880 21960 227319 22240
rect 749 20472 227319 21960
rect 880 20192 227319 20472
rect 749 18704 227319 20192
rect 880 18424 227319 18704
rect 749 16936 227319 18424
rect 880 16656 227319 16936
rect 749 15168 227319 16656
rect 880 14888 227319 15168
rect 749 13400 227319 14888
rect 880 13120 227319 13400
rect 749 11632 227319 13120
rect 880 11352 227319 11632
rect 749 9864 227319 11352
rect 880 9584 227319 9864
rect 749 8096 227319 9584
rect 880 7816 227319 8096
rect 749 6328 227319 7816
rect 880 6048 227319 6328
rect 749 4560 227319 6048
rect 880 4280 227319 4560
rect 749 2792 227319 4280
rect 880 2512 227319 2792
rect 749 1395 227319 2512
<< metal4 >>
rect 1794 2128 2414 227440
rect 19794 2128 20414 227440
rect 37794 2128 38414 227440
rect 55794 2128 56414 227440
rect 73794 2128 74414 227440
rect 91794 2128 92414 227440
rect 109794 2128 110414 227440
rect 127794 2128 128414 227440
rect 145794 2128 146414 227440
rect 163794 2128 164414 227440
rect 181794 2128 182414 227440
rect 199794 2128 200414 227440
rect 217794 2128 218414 227440
<< obsm4 >>
rect 979 3979 1714 227221
rect 2494 3979 19714 227221
rect 20494 3979 37714 227221
rect 38494 3979 55714 227221
rect 56494 3979 73714 227221
rect 74494 3979 91714 227221
rect 92494 3979 109714 227221
rect 110494 3979 127714 227221
rect 128494 3979 145714 227221
rect 146494 3979 163714 227221
rect 164494 3979 181714 227221
rect 182494 3979 199714 227221
rect 200494 3979 217714 227221
rect 218494 3979 224237 227221
<< labels >>
rlabel metal2 s 4250 229200 4306 230000 6 CLK
port 1 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 D1[0]
port 2 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 D1[10]
port 3 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 D1[11]
port 4 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 D1[12]
port 5 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 D1[13]
port 6 nsew signal output
rlabel metal3 s 0 27344 800 27464 6 D1[14]
port 7 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 D1[15]
port 8 nsew signal output
rlabel metal3 s 0 30880 800 31000 6 D1[16]
port 9 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 D1[17]
port 10 nsew signal output
rlabel metal3 s 0 34416 800 34536 6 D1[18]
port 11 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 D1[19]
port 12 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 D1[1]
port 13 nsew signal output
rlabel metal3 s 0 37952 800 38072 6 D1[20]
port 14 nsew signal output
rlabel metal3 s 0 39720 800 39840 6 D1[21]
port 15 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 D1[22]
port 16 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 D1[23]
port 17 nsew signal output
rlabel metal3 s 0 45024 800 45144 6 D1[24]
port 18 nsew signal output
rlabel metal3 s 0 46792 800 46912 6 D1[25]
port 19 nsew signal output
rlabel metal3 s 0 48560 800 48680 6 D1[26]
port 20 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 D1[27]
port 21 nsew signal output
rlabel metal3 s 0 52096 800 52216 6 D1[28]
port 22 nsew signal output
rlabel metal3 s 0 53864 800 53984 6 D1[29]
port 23 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 D1[2]
port 24 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 D1[30]
port 25 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 D1[31]
port 26 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 D1[32]
port 27 nsew signal output
rlabel metal3 s 0 60936 800 61056 6 D1[33]
port 28 nsew signal output
rlabel metal3 s 0 62704 800 62824 6 D1[34]
port 29 nsew signal output
rlabel metal3 s 0 64472 800 64592 6 D1[35]
port 30 nsew signal output
rlabel metal3 s 0 66240 800 66360 6 D1[36]
port 31 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 D1[37]
port 32 nsew signal output
rlabel metal3 s 0 69776 800 69896 6 D1[38]
port 33 nsew signal output
rlabel metal3 s 0 71544 800 71664 6 D1[39]
port 34 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 D1[3]
port 35 nsew signal output
rlabel metal3 s 0 73312 800 73432 6 D1[40]
port 36 nsew signal output
rlabel metal3 s 0 75080 800 75200 6 D1[41]
port 37 nsew signal output
rlabel metal3 s 0 76848 800 76968 6 D1[42]
port 38 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 D1[43]
port 39 nsew signal output
rlabel metal3 s 0 80384 800 80504 6 D1[44]
port 40 nsew signal output
rlabel metal3 s 0 82152 800 82272 6 D1[45]
port 41 nsew signal output
rlabel metal3 s 0 83920 800 84040 6 D1[46]
port 42 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 D1[47]
port 43 nsew signal output
rlabel metal3 s 0 87456 800 87576 6 D1[48]
port 44 nsew signal output
rlabel metal3 s 0 89224 800 89344 6 D1[49]
port 45 nsew signal output
rlabel metal3 s 0 9664 800 9784 6 D1[4]
port 46 nsew signal output
rlabel metal3 s 0 90992 800 91112 6 D1[50]
port 47 nsew signal output
rlabel metal3 s 0 92760 800 92880 6 D1[51]
port 48 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 D1[52]
port 49 nsew signal output
rlabel metal3 s 0 96296 800 96416 6 D1[53]
port 50 nsew signal output
rlabel metal3 s 0 98064 800 98184 6 D1[54]
port 51 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 D1[55]
port 52 nsew signal output
rlabel metal3 s 0 101600 800 101720 6 D1[56]
port 53 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 D1[57]
port 54 nsew signal output
rlabel metal3 s 0 105136 800 105256 6 D1[58]
port 55 nsew signal output
rlabel metal3 s 0 106904 800 107024 6 D1[59]
port 56 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 D1[5]
port 57 nsew signal output
rlabel metal3 s 0 108672 800 108792 6 D1[60]
port 58 nsew signal output
rlabel metal3 s 0 110440 800 110560 6 D1[61]
port 59 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 D1[62]
port 60 nsew signal output
rlabel metal3 s 0 113976 800 114096 6 D1[63]
port 61 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 D1[6]
port 62 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 D1[7]
port 63 nsew signal output
rlabel metal3 s 0 16736 800 16856 6 D1[8]
port 64 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 D1[9]
port 65 nsew signal output
rlabel metal3 s 0 115744 800 115864 6 D2[0]
port 66 nsew signal output
rlabel metal3 s 0 133424 800 133544 6 D2[10]
port 67 nsew signal output
rlabel metal3 s 0 135192 800 135312 6 D2[11]
port 68 nsew signal output
rlabel metal3 s 0 136960 800 137080 6 D2[12]
port 69 nsew signal output
rlabel metal3 s 0 138728 800 138848 6 D2[13]
port 70 nsew signal output
rlabel metal3 s 0 140496 800 140616 6 D2[14]
port 71 nsew signal output
rlabel metal3 s 0 142264 800 142384 6 D2[15]
port 72 nsew signal output
rlabel metal3 s 0 144032 800 144152 6 D2[16]
port 73 nsew signal output
rlabel metal3 s 0 145800 800 145920 6 D2[17]
port 74 nsew signal output
rlabel metal3 s 0 147568 800 147688 6 D2[18]
port 75 nsew signal output
rlabel metal3 s 0 149336 800 149456 6 D2[19]
port 76 nsew signal output
rlabel metal3 s 0 117512 800 117632 6 D2[1]
port 77 nsew signal output
rlabel metal3 s 0 151104 800 151224 6 D2[20]
port 78 nsew signal output
rlabel metal3 s 0 152872 800 152992 6 D2[21]
port 79 nsew signal output
rlabel metal3 s 0 154640 800 154760 6 D2[22]
port 80 nsew signal output
rlabel metal3 s 0 156408 800 156528 6 D2[23]
port 81 nsew signal output
rlabel metal3 s 0 158176 800 158296 6 D2[24]
port 82 nsew signal output
rlabel metal3 s 0 159944 800 160064 6 D2[25]
port 83 nsew signal output
rlabel metal3 s 0 161712 800 161832 6 D2[26]
port 84 nsew signal output
rlabel metal3 s 0 163480 800 163600 6 D2[27]
port 85 nsew signal output
rlabel metal3 s 0 165248 800 165368 6 D2[28]
port 86 nsew signal output
rlabel metal3 s 0 167016 800 167136 6 D2[29]
port 87 nsew signal output
rlabel metal3 s 0 119280 800 119400 6 D2[2]
port 88 nsew signal output
rlabel metal3 s 0 168784 800 168904 6 D2[30]
port 89 nsew signal output
rlabel metal3 s 0 170552 800 170672 6 D2[31]
port 90 nsew signal output
rlabel metal3 s 0 172320 800 172440 6 D2[32]
port 91 nsew signal output
rlabel metal3 s 0 174088 800 174208 6 D2[33]
port 92 nsew signal output
rlabel metal3 s 0 175856 800 175976 6 D2[34]
port 93 nsew signal output
rlabel metal3 s 0 177624 800 177744 6 D2[35]
port 94 nsew signal output
rlabel metal3 s 0 179392 800 179512 6 D2[36]
port 95 nsew signal output
rlabel metal3 s 0 181160 800 181280 6 D2[37]
port 96 nsew signal output
rlabel metal3 s 0 182928 800 183048 6 D2[38]
port 97 nsew signal output
rlabel metal3 s 0 184696 800 184816 6 D2[39]
port 98 nsew signal output
rlabel metal3 s 0 121048 800 121168 6 D2[3]
port 99 nsew signal output
rlabel metal3 s 0 186464 800 186584 6 D2[40]
port 100 nsew signal output
rlabel metal3 s 0 188232 800 188352 6 D2[41]
port 101 nsew signal output
rlabel metal3 s 0 190000 800 190120 6 D2[42]
port 102 nsew signal output
rlabel metal3 s 0 191768 800 191888 6 D2[43]
port 103 nsew signal output
rlabel metal3 s 0 193536 800 193656 6 D2[44]
port 104 nsew signal output
rlabel metal3 s 0 195304 800 195424 6 D2[45]
port 105 nsew signal output
rlabel metal3 s 0 197072 800 197192 6 D2[46]
port 106 nsew signal output
rlabel metal3 s 0 198840 800 198960 6 D2[47]
port 107 nsew signal output
rlabel metal3 s 0 200608 800 200728 6 D2[48]
port 108 nsew signal output
rlabel metal3 s 0 202376 800 202496 6 D2[49]
port 109 nsew signal output
rlabel metal3 s 0 122816 800 122936 6 D2[4]
port 110 nsew signal output
rlabel metal3 s 0 204144 800 204264 6 D2[50]
port 111 nsew signal output
rlabel metal3 s 0 205912 800 206032 6 D2[51]
port 112 nsew signal output
rlabel metal3 s 0 207680 800 207800 6 D2[52]
port 113 nsew signal output
rlabel metal3 s 0 209448 800 209568 6 D2[53]
port 114 nsew signal output
rlabel metal3 s 0 211216 800 211336 6 D2[54]
port 115 nsew signal output
rlabel metal3 s 0 212984 800 213104 6 D2[55]
port 116 nsew signal output
rlabel metal3 s 0 214752 800 214872 6 D2[56]
port 117 nsew signal output
rlabel metal3 s 0 216520 800 216640 6 D2[57]
port 118 nsew signal output
rlabel metal3 s 0 218288 800 218408 6 D2[58]
port 119 nsew signal output
rlabel metal3 s 0 220056 800 220176 6 D2[59]
port 120 nsew signal output
rlabel metal3 s 0 124584 800 124704 6 D2[5]
port 121 nsew signal output
rlabel metal3 s 0 221824 800 221944 6 D2[60]
port 122 nsew signal output
rlabel metal3 s 0 223592 800 223712 6 D2[61]
port 123 nsew signal output
rlabel metal3 s 0 225360 800 225480 6 D2[62]
port 124 nsew signal output
rlabel metal3 s 0 227128 800 227248 6 D2[63]
port 125 nsew signal output
rlabel metal3 s 0 126352 800 126472 6 D2[6]
port 126 nsew signal output
rlabel metal3 s 0 128120 800 128240 6 D2[7]
port 127 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 D2[8]
port 128 nsew signal output
rlabel metal3 s 0 131656 800 131776 6 D2[9]
port 129 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 D3[0]
port 130 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 D3[10]
port 131 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 D3[11]
port 132 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 D3[12]
port 133 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 D3[13]
port 134 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 D3[14]
port 135 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 D3[15]
port 136 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 D3[16]
port 137 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 D3[17]
port 138 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 D3[18]
port 139 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 D3[19]
port 140 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 D3[1]
port 141 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 D3[20]
port 142 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 D3[21]
port 143 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 D3[22]
port 144 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 D3[23]
port 145 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 D3[24]
port 146 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 D3[25]
port 147 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 D3[26]
port 148 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 D3[27]
port 149 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 D3[28]
port 150 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 D3[29]
port 151 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 D3[2]
port 152 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 D3[30]
port 153 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 D3[31]
port 154 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 D3[32]
port 155 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 D3[33]
port 156 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 D3[34]
port 157 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 D3[35]
port 158 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 D3[36]
port 159 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 D3[37]
port 160 nsew signal output
rlabel metal2 s 70398 0 70454 800 6 D3[38]
port 161 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 D3[39]
port 162 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 D3[3]
port 163 nsew signal output
rlabel metal2 s 73894 0 73950 800 6 D3[40]
port 164 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 D3[41]
port 165 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 D3[42]
port 166 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 D3[43]
port 167 nsew signal output
rlabel metal2 s 80886 0 80942 800 6 D3[44]
port 168 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 D3[45]
port 169 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 D3[46]
port 170 nsew signal output
rlabel metal2 s 86130 0 86186 800 6 D3[47]
port 171 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 D3[48]
port 172 nsew signal output
rlabel metal2 s 89626 0 89682 800 6 D3[49]
port 173 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 D3[4]
port 174 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 D3[50]
port 175 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 D3[51]
port 176 nsew signal output
rlabel metal2 s 94870 0 94926 800 6 D3[52]
port 177 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 D3[53]
port 178 nsew signal output
rlabel metal2 s 98366 0 98422 800 6 D3[54]
port 179 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 D3[55]
port 180 nsew signal output
rlabel metal2 s 101862 0 101918 800 6 D3[56]
port 181 nsew signal output
rlabel metal2 s 103610 0 103666 800 6 D3[57]
port 182 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 D3[58]
port 183 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 D3[59]
port 184 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 D3[5]
port 185 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 D3[60]
port 186 nsew signal output
rlabel metal2 s 110602 0 110658 800 6 D3[61]
port 187 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 D3[62]
port 188 nsew signal output
rlabel metal2 s 114098 0 114154 800 6 D3[63]
port 189 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 D3[6]
port 190 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 D3[7]
port 191 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 D3[8]
port 192 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 D3[9]
port 193 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 DW[0]
port 194 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 DW[10]
port 195 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 DW[11]
port 196 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 DW[12]
port 197 nsew signal input
rlabel metal2 s 138570 0 138626 800 6 DW[13]
port 198 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 DW[14]
port 199 nsew signal input
rlabel metal2 s 142066 0 142122 800 6 DW[15]
port 200 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 DW[16]
port 201 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 DW[17]
port 202 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 DW[18]
port 203 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 DW[19]
port 204 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 DW[1]
port 205 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 DW[20]
port 206 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 DW[21]
port 207 nsew signal input
rlabel metal2 s 154302 0 154358 800 6 DW[22]
port 208 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 DW[23]
port 209 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 DW[24]
port 210 nsew signal input
rlabel metal2 s 159546 0 159602 800 6 DW[25]
port 211 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 DW[26]
port 212 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 DW[27]
port 213 nsew signal input
rlabel metal2 s 164790 0 164846 800 6 DW[28]
port 214 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 DW[29]
port 215 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 DW[2]
port 216 nsew signal input
rlabel metal2 s 168286 0 168342 800 6 DW[30]
port 217 nsew signal input
rlabel metal2 s 170034 0 170090 800 6 DW[31]
port 218 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 DW[32]
port 219 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 DW[33]
port 220 nsew signal input
rlabel metal2 s 175278 0 175334 800 6 DW[34]
port 221 nsew signal input
rlabel metal2 s 177026 0 177082 800 6 DW[35]
port 222 nsew signal input
rlabel metal2 s 178774 0 178830 800 6 DW[36]
port 223 nsew signal input
rlabel metal2 s 180522 0 180578 800 6 DW[37]
port 224 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 DW[38]
port 225 nsew signal input
rlabel metal2 s 184018 0 184074 800 6 DW[39]
port 226 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 DW[3]
port 227 nsew signal input
rlabel metal2 s 185766 0 185822 800 6 DW[40]
port 228 nsew signal input
rlabel metal2 s 187514 0 187570 800 6 DW[41]
port 229 nsew signal input
rlabel metal2 s 189262 0 189318 800 6 DW[42]
port 230 nsew signal input
rlabel metal2 s 191010 0 191066 800 6 DW[43]
port 231 nsew signal input
rlabel metal2 s 192758 0 192814 800 6 DW[44]
port 232 nsew signal input
rlabel metal2 s 194506 0 194562 800 6 DW[45]
port 233 nsew signal input
rlabel metal2 s 196254 0 196310 800 6 DW[46]
port 234 nsew signal input
rlabel metal2 s 198002 0 198058 800 6 DW[47]
port 235 nsew signal input
rlabel metal2 s 199750 0 199806 800 6 DW[48]
port 236 nsew signal input
rlabel metal2 s 201498 0 201554 800 6 DW[49]
port 237 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 DW[4]
port 238 nsew signal input
rlabel metal2 s 203246 0 203302 800 6 DW[50]
port 239 nsew signal input
rlabel metal2 s 204994 0 205050 800 6 DW[51]
port 240 nsew signal input
rlabel metal2 s 206742 0 206798 800 6 DW[52]
port 241 nsew signal input
rlabel metal2 s 208490 0 208546 800 6 DW[53]
port 242 nsew signal input
rlabel metal2 s 210238 0 210294 800 6 DW[54]
port 243 nsew signal input
rlabel metal2 s 211986 0 212042 800 6 DW[55]
port 244 nsew signal input
rlabel metal2 s 213734 0 213790 800 6 DW[56]
port 245 nsew signal input
rlabel metal2 s 215482 0 215538 800 6 DW[57]
port 246 nsew signal input
rlabel metal2 s 217230 0 217286 800 6 DW[58]
port 247 nsew signal input
rlabel metal2 s 218978 0 219034 800 6 DW[59]
port 248 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 DW[5]
port 249 nsew signal input
rlabel metal2 s 220726 0 220782 800 6 DW[60]
port 250 nsew signal input
rlabel metal2 s 222474 0 222530 800 6 DW[61]
port 251 nsew signal input
rlabel metal2 s 224222 0 224278 800 6 DW[62]
port 252 nsew signal input
rlabel metal2 s 225970 0 226026 800 6 DW[63]
port 253 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 DW[6]
port 254 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 DW[7]
port 255 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 DW[8]
port 256 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 DW[9]
port 257 nsew signal input
rlabel metal2 s 19522 229200 19578 230000 6 R1[0]
port 258 nsew signal input
rlabel metal2 s 27158 229200 27214 230000 6 R1[1]
port 259 nsew signal input
rlabel metal2 s 34794 229200 34850 230000 6 R1[2]
port 260 nsew signal input
rlabel metal2 s 42430 229200 42486 230000 6 R1[3]
port 261 nsew signal input
rlabel metal2 s 50066 229200 50122 230000 6 R1[4]
port 262 nsew signal input
rlabel metal2 s 57702 229200 57758 230000 6 R1[5]
port 263 nsew signal input
rlabel metal2 s 65338 229200 65394 230000 6 R1[6]
port 264 nsew signal input
rlabel metal2 s 72974 229200 73030 230000 6 R2[0]
port 265 nsew signal input
rlabel metal2 s 80610 229200 80666 230000 6 R2[1]
port 266 nsew signal input
rlabel metal2 s 88246 229200 88302 230000 6 R2[2]
port 267 nsew signal input
rlabel metal2 s 95882 229200 95938 230000 6 R2[3]
port 268 nsew signal input
rlabel metal2 s 103518 229200 103574 230000 6 R2[4]
port 269 nsew signal input
rlabel metal2 s 111154 229200 111210 230000 6 R2[5]
port 270 nsew signal input
rlabel metal2 s 118790 229200 118846 230000 6 R2[6]
port 271 nsew signal input
rlabel metal2 s 126426 229200 126482 230000 6 R3[0]
port 272 nsew signal input
rlabel metal2 s 134062 229200 134118 230000 6 R3[1]
port 273 nsew signal input
rlabel metal2 s 141698 229200 141754 230000 6 R3[2]
port 274 nsew signal input
rlabel metal2 s 149334 229200 149390 230000 6 R3[3]
port 275 nsew signal input
rlabel metal2 s 156970 229200 157026 230000 6 R3[4]
port 276 nsew signal input
rlabel metal2 s 164606 229200 164662 230000 6 R3[5]
port 277 nsew signal input
rlabel metal2 s 172242 229200 172298 230000 6 R3[6]
port 278 nsew signal input
rlabel metal2 s 179878 229200 179934 230000 6 RW[0]
port 279 nsew signal input
rlabel metal2 s 187514 229200 187570 230000 6 RW[1]
port 280 nsew signal input
rlabel metal2 s 195150 229200 195206 230000 6 RW[2]
port 281 nsew signal input
rlabel metal2 s 202786 229200 202842 230000 6 RW[3]
port 282 nsew signal input
rlabel metal2 s 210422 229200 210478 230000 6 RW[4]
port 283 nsew signal input
rlabel metal2 s 218058 229200 218114 230000 6 RW[5]
port 284 nsew signal input
rlabel metal2 s 225694 229200 225750 230000 6 RW[6]
port 285 nsew signal input
rlabel metal4 s 19794 2128 20414 227440 6 VGND
port 286 nsew ground bidirectional
rlabel metal4 s 55794 2128 56414 227440 6 VGND
port 286 nsew ground bidirectional
rlabel metal4 s 91794 2128 92414 227440 6 VGND
port 286 nsew ground bidirectional
rlabel metal4 s 127794 2128 128414 227440 6 VGND
port 286 nsew ground bidirectional
rlabel metal4 s 163794 2128 164414 227440 6 VGND
port 286 nsew ground bidirectional
rlabel metal4 s 199794 2128 200414 227440 6 VGND
port 286 nsew ground bidirectional
rlabel metal4 s 1794 2128 2414 227440 6 VPWR
port 287 nsew power bidirectional
rlabel metal4 s 37794 2128 38414 227440 6 VPWR
port 287 nsew power bidirectional
rlabel metal4 s 73794 2128 74414 227440 6 VPWR
port 287 nsew power bidirectional
rlabel metal4 s 109794 2128 110414 227440 6 VPWR
port 287 nsew power bidirectional
rlabel metal4 s 145794 2128 146414 227440 6 VPWR
port 287 nsew power bidirectional
rlabel metal4 s 181794 2128 182414 227440 6 VPWR
port 287 nsew power bidirectional
rlabel metal4 s 217794 2128 218414 227440 6 VPWR
port 287 nsew power bidirectional
rlabel metal2 s 11886 229200 11942 230000 6 WE
port 288 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 230000 230000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 123319116
string GDS_FILE /scratch/mpw7/caravel_user_project/openlane/Microwatt_FP_DFFRFile/runs/22_07_11_21_36/results/signoff/Microwatt_FP_DFFRFile.magic.gds
string GDS_START 583198
<< end >>

