magic
tech sky130B
magscale 1 2
timestamp 1662419477
<< obsli1 >>
rect 1104 2159 138828 137649
<< obsm1 >>
rect 474 824 139734 137680
<< metal2 >>
rect 3238 139200 3294 140000
rect 8574 139200 8630 140000
rect 13910 139200 13966 140000
rect 19246 139200 19302 140000
rect 24582 139200 24638 140000
rect 29918 139200 29974 140000
rect 35254 139200 35310 140000
rect 40590 139200 40646 140000
rect 45926 139200 45982 140000
rect 51262 139200 51318 140000
rect 56598 139200 56654 140000
rect 61934 139200 61990 140000
rect 67270 139200 67326 140000
rect 72606 139200 72662 140000
rect 77942 139200 77998 140000
rect 83278 139200 83334 140000
rect 88614 139200 88670 140000
rect 93950 139200 94006 140000
rect 99286 139200 99342 140000
rect 104622 139200 104678 140000
rect 109958 139200 110014 140000
rect 115294 139200 115350 140000
rect 120630 139200 120686 140000
rect 125966 139200 126022 140000
rect 131302 139200 131358 140000
rect 136638 139200 136694 140000
rect 5722 0 5778 800
rect 6734 0 6790 800
rect 7746 0 7802 800
rect 8758 0 8814 800
rect 9770 0 9826 800
rect 10782 0 10838 800
rect 11794 0 11850 800
rect 12806 0 12862 800
rect 13818 0 13874 800
rect 14830 0 14886 800
rect 15842 0 15898 800
rect 16854 0 16910 800
rect 17866 0 17922 800
rect 18878 0 18934 800
rect 19890 0 19946 800
rect 20902 0 20958 800
rect 21914 0 21970 800
rect 22926 0 22982 800
rect 23938 0 23994 800
rect 24950 0 25006 800
rect 25962 0 26018 800
rect 26974 0 27030 800
rect 27986 0 28042 800
rect 28998 0 29054 800
rect 30010 0 30066 800
rect 31022 0 31078 800
rect 32034 0 32090 800
rect 33046 0 33102 800
rect 34058 0 34114 800
rect 35070 0 35126 800
rect 36082 0 36138 800
rect 37094 0 37150 800
rect 38106 0 38162 800
rect 39118 0 39174 800
rect 40130 0 40186 800
rect 41142 0 41198 800
rect 42154 0 42210 800
rect 43166 0 43222 800
rect 44178 0 44234 800
rect 45190 0 45246 800
rect 46202 0 46258 800
rect 47214 0 47270 800
rect 48226 0 48282 800
rect 49238 0 49294 800
rect 50250 0 50306 800
rect 51262 0 51318 800
rect 52274 0 52330 800
rect 53286 0 53342 800
rect 54298 0 54354 800
rect 55310 0 55366 800
rect 56322 0 56378 800
rect 57334 0 57390 800
rect 58346 0 58402 800
rect 59358 0 59414 800
rect 60370 0 60426 800
rect 61382 0 61438 800
rect 62394 0 62450 800
rect 63406 0 63462 800
rect 64418 0 64474 800
rect 65430 0 65486 800
rect 66442 0 66498 800
rect 67454 0 67510 800
rect 68466 0 68522 800
rect 69478 0 69534 800
rect 70490 0 70546 800
rect 71502 0 71558 800
rect 72514 0 72570 800
rect 73526 0 73582 800
rect 74538 0 74594 800
rect 75550 0 75606 800
rect 76562 0 76618 800
rect 77574 0 77630 800
rect 78586 0 78642 800
rect 79598 0 79654 800
rect 80610 0 80666 800
rect 81622 0 81678 800
rect 82634 0 82690 800
rect 83646 0 83702 800
rect 84658 0 84714 800
rect 85670 0 85726 800
rect 86682 0 86738 800
rect 87694 0 87750 800
rect 88706 0 88762 800
rect 89718 0 89774 800
rect 90730 0 90786 800
rect 91742 0 91798 800
rect 92754 0 92810 800
rect 93766 0 93822 800
rect 94778 0 94834 800
rect 95790 0 95846 800
rect 96802 0 96858 800
rect 97814 0 97870 800
rect 98826 0 98882 800
rect 99838 0 99894 800
rect 100850 0 100906 800
rect 101862 0 101918 800
rect 102874 0 102930 800
rect 103886 0 103942 800
rect 104898 0 104954 800
rect 105910 0 105966 800
rect 106922 0 106978 800
rect 107934 0 107990 800
rect 108946 0 109002 800
rect 109958 0 110014 800
rect 110970 0 111026 800
rect 111982 0 112038 800
rect 112994 0 113050 800
rect 114006 0 114062 800
rect 115018 0 115074 800
rect 116030 0 116086 800
rect 117042 0 117098 800
rect 118054 0 118110 800
rect 119066 0 119122 800
rect 120078 0 120134 800
rect 121090 0 121146 800
rect 122102 0 122158 800
rect 123114 0 123170 800
rect 124126 0 124182 800
rect 125138 0 125194 800
rect 126150 0 126206 800
rect 127162 0 127218 800
rect 128174 0 128230 800
rect 129186 0 129242 800
rect 130198 0 130254 800
rect 131210 0 131266 800
rect 132222 0 132278 800
rect 133234 0 133290 800
rect 134246 0 134302 800
<< obsm2 >>
rect 480 139144 3182 139346
rect 3350 139144 8518 139346
rect 8686 139144 13854 139346
rect 14022 139144 19190 139346
rect 19358 139144 24526 139346
rect 24694 139144 29862 139346
rect 30030 139144 35198 139346
rect 35366 139144 40534 139346
rect 40702 139144 45870 139346
rect 46038 139144 51206 139346
rect 51374 139144 56542 139346
rect 56710 139144 61878 139346
rect 62046 139144 67214 139346
rect 67382 139144 72550 139346
rect 72718 139144 77886 139346
rect 78054 139144 83222 139346
rect 83390 139144 88558 139346
rect 88726 139144 93894 139346
rect 94062 139144 99230 139346
rect 99398 139144 104566 139346
rect 104734 139144 109902 139346
rect 110070 139144 115238 139346
rect 115406 139144 120574 139346
rect 120742 139144 125910 139346
rect 126078 139144 131246 139346
rect 131414 139144 136582 139346
rect 136750 139144 139728 139346
rect 480 856 139728 139144
rect 480 734 5666 856
rect 5834 734 6678 856
rect 6846 734 7690 856
rect 7858 734 8702 856
rect 8870 734 9714 856
rect 9882 734 10726 856
rect 10894 734 11738 856
rect 11906 734 12750 856
rect 12918 734 13762 856
rect 13930 734 14774 856
rect 14942 734 15786 856
rect 15954 734 16798 856
rect 16966 734 17810 856
rect 17978 734 18822 856
rect 18990 734 19834 856
rect 20002 734 20846 856
rect 21014 734 21858 856
rect 22026 734 22870 856
rect 23038 734 23882 856
rect 24050 734 24894 856
rect 25062 734 25906 856
rect 26074 734 26918 856
rect 27086 734 27930 856
rect 28098 734 28942 856
rect 29110 734 29954 856
rect 30122 734 30966 856
rect 31134 734 31978 856
rect 32146 734 32990 856
rect 33158 734 34002 856
rect 34170 734 35014 856
rect 35182 734 36026 856
rect 36194 734 37038 856
rect 37206 734 38050 856
rect 38218 734 39062 856
rect 39230 734 40074 856
rect 40242 734 41086 856
rect 41254 734 42098 856
rect 42266 734 43110 856
rect 43278 734 44122 856
rect 44290 734 45134 856
rect 45302 734 46146 856
rect 46314 734 47158 856
rect 47326 734 48170 856
rect 48338 734 49182 856
rect 49350 734 50194 856
rect 50362 734 51206 856
rect 51374 734 52218 856
rect 52386 734 53230 856
rect 53398 734 54242 856
rect 54410 734 55254 856
rect 55422 734 56266 856
rect 56434 734 57278 856
rect 57446 734 58290 856
rect 58458 734 59302 856
rect 59470 734 60314 856
rect 60482 734 61326 856
rect 61494 734 62338 856
rect 62506 734 63350 856
rect 63518 734 64362 856
rect 64530 734 65374 856
rect 65542 734 66386 856
rect 66554 734 67398 856
rect 67566 734 68410 856
rect 68578 734 69422 856
rect 69590 734 70434 856
rect 70602 734 71446 856
rect 71614 734 72458 856
rect 72626 734 73470 856
rect 73638 734 74482 856
rect 74650 734 75494 856
rect 75662 734 76506 856
rect 76674 734 77518 856
rect 77686 734 78530 856
rect 78698 734 79542 856
rect 79710 734 80554 856
rect 80722 734 81566 856
rect 81734 734 82578 856
rect 82746 734 83590 856
rect 83758 734 84602 856
rect 84770 734 85614 856
rect 85782 734 86626 856
rect 86794 734 87638 856
rect 87806 734 88650 856
rect 88818 734 89662 856
rect 89830 734 90674 856
rect 90842 734 91686 856
rect 91854 734 92698 856
rect 92866 734 93710 856
rect 93878 734 94722 856
rect 94890 734 95734 856
rect 95902 734 96746 856
rect 96914 734 97758 856
rect 97926 734 98770 856
rect 98938 734 99782 856
rect 99950 734 100794 856
rect 100962 734 101806 856
rect 101974 734 102818 856
rect 102986 734 103830 856
rect 103998 734 104842 856
rect 105010 734 105854 856
rect 106022 734 106866 856
rect 107034 734 107878 856
rect 108046 734 108890 856
rect 109058 734 109902 856
rect 110070 734 110914 856
rect 111082 734 111926 856
rect 112094 734 112938 856
rect 113106 734 113950 856
rect 114118 734 114962 856
rect 115130 734 115974 856
rect 116142 734 116986 856
rect 117154 734 117998 856
rect 118166 734 119010 856
rect 119178 734 120022 856
rect 120190 734 121034 856
rect 121202 734 122046 856
rect 122214 734 123058 856
rect 123226 734 124070 856
rect 124238 734 125082 856
rect 125250 734 126094 856
rect 126262 734 127106 856
rect 127274 734 128118 856
rect 128286 734 129130 856
rect 129298 734 130142 856
rect 130310 734 131154 856
rect 131322 734 132166 856
rect 132334 734 133178 856
rect 133346 734 134190 856
rect 134358 734 139728 856
<< metal3 >>
rect 0 139000 800 139120
rect 0 137912 800 138032
rect 0 136824 800 136944
rect 0 135736 800 135856
rect 0 134648 800 134768
rect 0 133560 800 133680
rect 0 132472 800 132592
rect 0 131384 800 131504
rect 0 130296 800 130416
rect 0 129208 800 129328
rect 0 128120 800 128240
rect 0 127032 800 127152
rect 0 125944 800 126064
rect 0 124856 800 124976
rect 0 123768 800 123888
rect 0 122680 800 122800
rect 0 121592 800 121712
rect 0 120504 800 120624
rect 0 119416 800 119536
rect 0 118328 800 118448
rect 0 117240 800 117360
rect 0 116152 800 116272
rect 0 115064 800 115184
rect 0 113976 800 114096
rect 0 112888 800 113008
rect 0 111800 800 111920
rect 0 110712 800 110832
rect 0 109624 800 109744
rect 0 108536 800 108656
rect 0 107448 800 107568
rect 0 106360 800 106480
rect 0 105272 800 105392
rect 0 104184 800 104304
rect 0 103096 800 103216
rect 0 102008 800 102128
rect 0 100920 800 101040
rect 0 99832 800 99952
rect 0 98744 800 98864
rect 0 97656 800 97776
rect 0 96568 800 96688
rect 0 95480 800 95600
rect 0 94392 800 94512
rect 0 93304 800 93424
rect 0 92216 800 92336
rect 0 91128 800 91248
rect 0 90040 800 90160
rect 0 88952 800 89072
rect 0 87864 800 87984
rect 0 86776 800 86896
rect 0 85688 800 85808
rect 0 84600 800 84720
rect 0 83512 800 83632
rect 0 82424 800 82544
rect 0 81336 800 81456
rect 0 80248 800 80368
rect 0 79160 800 79280
rect 0 78072 800 78192
rect 0 76984 800 77104
rect 0 75896 800 76016
rect 0 74808 800 74928
rect 0 73720 800 73840
rect 0 72632 800 72752
rect 0 71544 800 71664
rect 0 70456 800 70576
rect 0 69368 800 69488
rect 0 68280 800 68400
rect 0 67192 800 67312
rect 0 66104 800 66224
rect 0 65016 800 65136
rect 0 63928 800 64048
rect 0 62840 800 62960
rect 0 61752 800 61872
rect 0 60664 800 60784
rect 0 59576 800 59696
rect 0 58488 800 58608
rect 0 57400 800 57520
rect 0 56312 800 56432
rect 0 55224 800 55344
rect 0 54136 800 54256
rect 0 53048 800 53168
rect 0 51960 800 52080
rect 0 50872 800 50992
rect 0 49784 800 49904
rect 0 48696 800 48816
rect 0 47608 800 47728
rect 0 46520 800 46640
rect 0 45432 800 45552
rect 0 44344 800 44464
rect 0 43256 800 43376
rect 0 42168 800 42288
rect 0 41080 800 41200
rect 0 39992 800 40112
rect 0 38904 800 39024
rect 0 37816 800 37936
rect 0 36728 800 36848
rect 0 35640 800 35760
rect 0 34552 800 34672
rect 0 33464 800 33584
rect 0 32376 800 32496
rect 0 31288 800 31408
rect 0 30200 800 30320
rect 0 29112 800 29232
rect 0 28024 800 28144
rect 0 26936 800 27056
rect 0 25848 800 25968
rect 0 24760 800 24880
rect 0 23672 800 23792
rect 0 22584 800 22704
rect 0 21496 800 21616
rect 0 20408 800 20528
rect 0 19320 800 19440
rect 0 18232 800 18352
rect 0 17144 800 17264
rect 0 16056 800 16176
rect 0 14968 800 15088
rect 0 13880 800 14000
rect 0 12792 800 12912
rect 0 11704 800 11824
rect 0 10616 800 10736
rect 0 9528 800 9648
rect 0 8440 800 8560
rect 0 7352 800 7472
rect 0 6264 800 6384
rect 0 5176 800 5296
rect 0 4088 800 4208
rect 0 3000 800 3120
rect 0 1912 800 2032
rect 0 824 800 944
<< obsm3 >>
rect 880 138920 139367 139093
rect 606 138112 139367 138920
rect 880 137832 139367 138112
rect 606 137024 139367 137832
rect 880 136744 139367 137024
rect 606 135936 139367 136744
rect 880 135656 139367 135936
rect 606 134848 139367 135656
rect 880 134568 139367 134848
rect 606 133760 139367 134568
rect 880 133480 139367 133760
rect 606 132672 139367 133480
rect 880 132392 139367 132672
rect 606 131584 139367 132392
rect 880 131304 139367 131584
rect 606 130496 139367 131304
rect 880 130216 139367 130496
rect 606 129408 139367 130216
rect 880 129128 139367 129408
rect 606 128320 139367 129128
rect 880 128040 139367 128320
rect 606 127232 139367 128040
rect 880 126952 139367 127232
rect 606 126144 139367 126952
rect 880 125864 139367 126144
rect 606 125056 139367 125864
rect 880 124776 139367 125056
rect 606 123968 139367 124776
rect 880 123688 139367 123968
rect 606 122880 139367 123688
rect 880 122600 139367 122880
rect 606 121792 139367 122600
rect 880 121512 139367 121792
rect 606 120704 139367 121512
rect 880 120424 139367 120704
rect 606 119616 139367 120424
rect 880 119336 139367 119616
rect 606 118528 139367 119336
rect 880 118248 139367 118528
rect 606 117440 139367 118248
rect 880 117160 139367 117440
rect 606 116352 139367 117160
rect 880 116072 139367 116352
rect 606 115264 139367 116072
rect 880 114984 139367 115264
rect 606 114176 139367 114984
rect 880 113896 139367 114176
rect 606 113088 139367 113896
rect 880 112808 139367 113088
rect 606 112000 139367 112808
rect 880 111720 139367 112000
rect 606 110912 139367 111720
rect 880 110632 139367 110912
rect 606 109824 139367 110632
rect 880 109544 139367 109824
rect 606 108736 139367 109544
rect 880 108456 139367 108736
rect 606 107648 139367 108456
rect 880 107368 139367 107648
rect 606 106560 139367 107368
rect 880 106280 139367 106560
rect 606 105472 139367 106280
rect 880 105192 139367 105472
rect 606 104384 139367 105192
rect 880 104104 139367 104384
rect 606 103296 139367 104104
rect 880 103016 139367 103296
rect 606 102208 139367 103016
rect 880 101928 139367 102208
rect 606 101120 139367 101928
rect 880 100840 139367 101120
rect 606 100032 139367 100840
rect 880 99752 139367 100032
rect 606 98944 139367 99752
rect 880 98664 139367 98944
rect 606 97856 139367 98664
rect 880 97576 139367 97856
rect 606 96768 139367 97576
rect 880 96488 139367 96768
rect 606 95680 139367 96488
rect 880 95400 139367 95680
rect 606 94592 139367 95400
rect 880 94312 139367 94592
rect 606 93504 139367 94312
rect 880 93224 139367 93504
rect 606 92416 139367 93224
rect 880 92136 139367 92416
rect 606 91328 139367 92136
rect 880 91048 139367 91328
rect 606 90240 139367 91048
rect 880 89960 139367 90240
rect 606 89152 139367 89960
rect 880 88872 139367 89152
rect 606 88064 139367 88872
rect 880 87784 139367 88064
rect 606 86976 139367 87784
rect 880 86696 139367 86976
rect 606 85888 139367 86696
rect 880 85608 139367 85888
rect 606 84800 139367 85608
rect 880 84520 139367 84800
rect 606 83712 139367 84520
rect 880 83432 139367 83712
rect 606 82624 139367 83432
rect 880 82344 139367 82624
rect 606 81536 139367 82344
rect 880 81256 139367 81536
rect 606 80448 139367 81256
rect 880 80168 139367 80448
rect 606 79360 139367 80168
rect 880 79080 139367 79360
rect 606 78272 139367 79080
rect 880 77992 139367 78272
rect 606 77184 139367 77992
rect 880 76904 139367 77184
rect 606 76096 139367 76904
rect 880 75816 139367 76096
rect 606 75008 139367 75816
rect 880 74728 139367 75008
rect 606 73920 139367 74728
rect 880 73640 139367 73920
rect 606 72832 139367 73640
rect 880 72552 139367 72832
rect 606 71744 139367 72552
rect 880 71464 139367 71744
rect 606 70656 139367 71464
rect 880 70376 139367 70656
rect 606 69568 139367 70376
rect 880 69288 139367 69568
rect 606 68480 139367 69288
rect 880 68200 139367 68480
rect 606 67392 139367 68200
rect 880 67112 139367 67392
rect 606 66304 139367 67112
rect 880 66024 139367 66304
rect 606 65216 139367 66024
rect 880 64936 139367 65216
rect 606 64128 139367 64936
rect 880 63848 139367 64128
rect 606 63040 139367 63848
rect 880 62760 139367 63040
rect 606 61952 139367 62760
rect 880 61672 139367 61952
rect 606 60864 139367 61672
rect 880 60584 139367 60864
rect 606 59776 139367 60584
rect 880 59496 139367 59776
rect 606 58688 139367 59496
rect 880 58408 139367 58688
rect 606 57600 139367 58408
rect 880 57320 139367 57600
rect 606 56512 139367 57320
rect 880 56232 139367 56512
rect 606 55424 139367 56232
rect 880 55144 139367 55424
rect 606 54336 139367 55144
rect 880 54056 139367 54336
rect 606 53248 139367 54056
rect 880 52968 139367 53248
rect 606 52160 139367 52968
rect 880 51880 139367 52160
rect 606 51072 139367 51880
rect 880 50792 139367 51072
rect 606 49984 139367 50792
rect 880 49704 139367 49984
rect 606 48896 139367 49704
rect 880 48616 139367 48896
rect 606 47808 139367 48616
rect 880 47528 139367 47808
rect 606 46720 139367 47528
rect 880 46440 139367 46720
rect 606 45632 139367 46440
rect 880 45352 139367 45632
rect 606 44544 139367 45352
rect 880 44264 139367 44544
rect 606 43456 139367 44264
rect 880 43176 139367 43456
rect 606 42368 139367 43176
rect 880 42088 139367 42368
rect 606 41280 139367 42088
rect 880 41000 139367 41280
rect 606 40192 139367 41000
rect 880 39912 139367 40192
rect 606 39104 139367 39912
rect 880 38824 139367 39104
rect 606 38016 139367 38824
rect 880 37736 139367 38016
rect 606 36928 139367 37736
rect 880 36648 139367 36928
rect 606 35840 139367 36648
rect 880 35560 139367 35840
rect 606 34752 139367 35560
rect 880 34472 139367 34752
rect 606 33664 139367 34472
rect 880 33384 139367 33664
rect 606 32576 139367 33384
rect 880 32296 139367 32576
rect 606 31488 139367 32296
rect 880 31208 139367 31488
rect 606 30400 139367 31208
rect 880 30120 139367 30400
rect 606 29312 139367 30120
rect 880 29032 139367 29312
rect 606 28224 139367 29032
rect 880 27944 139367 28224
rect 606 27136 139367 27944
rect 880 26856 139367 27136
rect 606 26048 139367 26856
rect 880 25768 139367 26048
rect 606 24960 139367 25768
rect 880 24680 139367 24960
rect 606 23872 139367 24680
rect 880 23592 139367 23872
rect 606 22784 139367 23592
rect 880 22504 139367 22784
rect 606 21696 139367 22504
rect 880 21416 139367 21696
rect 606 20608 139367 21416
rect 880 20328 139367 20608
rect 606 19520 139367 20328
rect 880 19240 139367 19520
rect 606 18432 139367 19240
rect 880 18152 139367 18432
rect 606 17344 139367 18152
rect 880 17064 139367 17344
rect 606 16256 139367 17064
rect 880 15976 139367 16256
rect 606 15168 139367 15976
rect 880 14888 139367 15168
rect 606 14080 139367 14888
rect 880 13800 139367 14080
rect 606 12992 139367 13800
rect 880 12712 139367 12992
rect 606 11904 139367 12712
rect 880 11624 139367 11904
rect 606 10816 139367 11624
rect 880 10536 139367 10816
rect 606 9728 139367 10536
rect 880 9448 139367 9728
rect 606 8640 139367 9448
rect 880 8360 139367 8640
rect 606 7552 139367 8360
rect 880 7272 139367 7552
rect 606 6464 139367 7272
rect 880 6184 139367 6464
rect 606 5376 139367 6184
rect 880 5096 139367 5376
rect 606 4288 139367 5096
rect 880 4008 139367 4288
rect 606 3200 139367 4008
rect 880 2920 139367 3200
rect 606 2112 139367 2920
rect 880 1832 139367 2112
rect 606 1024 139367 1832
rect 880 851 139367 1024
<< metal4 >>
rect 1794 2128 2414 137680
rect 19794 2128 20414 137680
rect 37794 2128 38414 137680
rect 55794 2128 56414 137680
rect 73794 2128 74414 137680
rect 91794 2128 92414 137680
rect 109794 2128 110414 137680
rect 127794 2128 128414 137680
<< obsm4 >>
rect 611 2211 1714 137325
rect 2494 2211 19714 137325
rect 20494 2211 37714 137325
rect 38494 2211 55714 137325
rect 56494 2211 73714 137325
rect 74494 2211 91714 137325
rect 92494 2211 109714 137325
rect 110494 2211 127714 137325
rect 128494 2211 137389 137325
<< labels >>
rlabel metal2 s 3238 139200 3294 140000 6 CLK
port 1 nsew signal input
rlabel metal3 s 0 824 800 944 6 D1[0]
port 2 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 D1[10]
port 3 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 D1[11]
port 4 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 D1[12]
port 5 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 D1[13]
port 6 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 D1[14]
port 7 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 D1[15]
port 8 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 D1[16]
port 9 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 D1[17]
port 10 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 D1[18]
port 11 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 D1[19]
port 12 nsew signal output
rlabel metal3 s 0 1912 800 2032 6 D1[1]
port 13 nsew signal output
rlabel metal3 s 0 22584 800 22704 6 D1[20]
port 14 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 D1[21]
port 15 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 D1[22]
port 16 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 D1[23]
port 17 nsew signal output
rlabel metal3 s 0 26936 800 27056 6 D1[24]
port 18 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 D1[25]
port 19 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 D1[26]
port 20 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 D1[27]
port 21 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 D1[28]
port 22 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 D1[29]
port 23 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 D1[2]
port 24 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 D1[30]
port 25 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 D1[31]
port 26 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 D1[32]
port 27 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 D1[33]
port 28 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 D1[34]
port 29 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 D1[35]
port 30 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 D1[36]
port 31 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 D1[37]
port 32 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 D1[38]
port 33 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 D1[39]
port 34 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 D1[3]
port 35 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 D1[40]
port 36 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 D1[41]
port 37 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 D1[42]
port 38 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 D1[43]
port 39 nsew signal output
rlabel metal3 s 0 48696 800 48816 6 D1[44]
port 40 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 D1[45]
port 41 nsew signal output
rlabel metal3 s 0 50872 800 50992 6 D1[46]
port 42 nsew signal output
rlabel metal3 s 0 51960 800 52080 6 D1[47]
port 43 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 D1[48]
port 44 nsew signal output
rlabel metal3 s 0 54136 800 54256 6 D1[49]
port 45 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 D1[4]
port 46 nsew signal output
rlabel metal3 s 0 55224 800 55344 6 D1[50]
port 47 nsew signal output
rlabel metal3 s 0 56312 800 56432 6 D1[51]
port 48 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 D1[52]
port 49 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 D1[53]
port 50 nsew signal output
rlabel metal3 s 0 59576 800 59696 6 D1[54]
port 51 nsew signal output
rlabel metal3 s 0 60664 800 60784 6 D1[55]
port 52 nsew signal output
rlabel metal3 s 0 61752 800 61872 6 D1[56]
port 53 nsew signal output
rlabel metal3 s 0 62840 800 62960 6 D1[57]
port 54 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 D1[58]
port 55 nsew signal output
rlabel metal3 s 0 65016 800 65136 6 D1[59]
port 56 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 D1[5]
port 57 nsew signal output
rlabel metal3 s 0 66104 800 66224 6 D1[60]
port 58 nsew signal output
rlabel metal3 s 0 67192 800 67312 6 D1[61]
port 59 nsew signal output
rlabel metal3 s 0 68280 800 68400 6 D1[62]
port 60 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 D1[63]
port 61 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 D1[6]
port 62 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 D1[7]
port 63 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 D1[8]
port 64 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 D1[9]
port 65 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 D2[0]
port 66 nsew signal output
rlabel metal3 s 0 81336 800 81456 6 D2[10]
port 67 nsew signal output
rlabel metal3 s 0 82424 800 82544 6 D2[11]
port 68 nsew signal output
rlabel metal3 s 0 83512 800 83632 6 D2[12]
port 69 nsew signal output
rlabel metal3 s 0 84600 800 84720 6 D2[13]
port 70 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 D2[14]
port 71 nsew signal output
rlabel metal3 s 0 86776 800 86896 6 D2[15]
port 72 nsew signal output
rlabel metal3 s 0 87864 800 87984 6 D2[16]
port 73 nsew signal output
rlabel metal3 s 0 88952 800 89072 6 D2[17]
port 74 nsew signal output
rlabel metal3 s 0 90040 800 90160 6 D2[18]
port 75 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 D2[19]
port 76 nsew signal output
rlabel metal3 s 0 71544 800 71664 6 D2[1]
port 77 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 D2[20]
port 78 nsew signal output
rlabel metal3 s 0 93304 800 93424 6 D2[21]
port 79 nsew signal output
rlabel metal3 s 0 94392 800 94512 6 D2[22]
port 80 nsew signal output
rlabel metal3 s 0 95480 800 95600 6 D2[23]
port 81 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 D2[24]
port 82 nsew signal output
rlabel metal3 s 0 97656 800 97776 6 D2[25]
port 83 nsew signal output
rlabel metal3 s 0 98744 800 98864 6 D2[26]
port 84 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 D2[27]
port 85 nsew signal output
rlabel metal3 s 0 100920 800 101040 6 D2[28]
port 86 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 D2[29]
port 87 nsew signal output
rlabel metal3 s 0 72632 800 72752 6 D2[2]
port 88 nsew signal output
rlabel metal3 s 0 103096 800 103216 6 D2[30]
port 89 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 D2[31]
port 90 nsew signal output
rlabel metal3 s 0 105272 800 105392 6 D2[32]
port 91 nsew signal output
rlabel metal3 s 0 106360 800 106480 6 D2[33]
port 92 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 D2[34]
port 93 nsew signal output
rlabel metal3 s 0 108536 800 108656 6 D2[35]
port 94 nsew signal output
rlabel metal3 s 0 109624 800 109744 6 D2[36]
port 95 nsew signal output
rlabel metal3 s 0 110712 800 110832 6 D2[37]
port 96 nsew signal output
rlabel metal3 s 0 111800 800 111920 6 D2[38]
port 97 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 D2[39]
port 98 nsew signal output
rlabel metal3 s 0 73720 800 73840 6 D2[3]
port 99 nsew signal output
rlabel metal3 s 0 113976 800 114096 6 D2[40]
port 100 nsew signal output
rlabel metal3 s 0 115064 800 115184 6 D2[41]
port 101 nsew signal output
rlabel metal3 s 0 116152 800 116272 6 D2[42]
port 102 nsew signal output
rlabel metal3 s 0 117240 800 117360 6 D2[43]
port 103 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 D2[44]
port 104 nsew signal output
rlabel metal3 s 0 119416 800 119536 6 D2[45]
port 105 nsew signal output
rlabel metal3 s 0 120504 800 120624 6 D2[46]
port 106 nsew signal output
rlabel metal3 s 0 121592 800 121712 6 D2[47]
port 107 nsew signal output
rlabel metal3 s 0 122680 800 122800 6 D2[48]
port 108 nsew signal output
rlabel metal3 s 0 123768 800 123888 6 D2[49]
port 109 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 D2[4]
port 110 nsew signal output
rlabel metal3 s 0 124856 800 124976 6 D2[50]
port 111 nsew signal output
rlabel metal3 s 0 125944 800 126064 6 D2[51]
port 112 nsew signal output
rlabel metal3 s 0 127032 800 127152 6 D2[52]
port 113 nsew signal output
rlabel metal3 s 0 128120 800 128240 6 D2[53]
port 114 nsew signal output
rlabel metal3 s 0 129208 800 129328 6 D2[54]
port 115 nsew signal output
rlabel metal3 s 0 130296 800 130416 6 D2[55]
port 116 nsew signal output
rlabel metal3 s 0 131384 800 131504 6 D2[56]
port 117 nsew signal output
rlabel metal3 s 0 132472 800 132592 6 D2[57]
port 118 nsew signal output
rlabel metal3 s 0 133560 800 133680 6 D2[58]
port 119 nsew signal output
rlabel metal3 s 0 134648 800 134768 6 D2[59]
port 120 nsew signal output
rlabel metal3 s 0 75896 800 76016 6 D2[5]
port 121 nsew signal output
rlabel metal3 s 0 135736 800 135856 6 D2[60]
port 122 nsew signal output
rlabel metal3 s 0 136824 800 136944 6 D2[61]
port 123 nsew signal output
rlabel metal3 s 0 137912 800 138032 6 D2[62]
port 124 nsew signal output
rlabel metal3 s 0 139000 800 139120 6 D2[63]
port 125 nsew signal output
rlabel metal3 s 0 76984 800 77104 6 D2[6]
port 126 nsew signal output
rlabel metal3 s 0 78072 800 78192 6 D2[7]
port 127 nsew signal output
rlabel metal3 s 0 79160 800 79280 6 D2[8]
port 128 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 D2[9]
port 129 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 D3[0]
port 130 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 D3[10]
port 131 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 D3[11]
port 132 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 D3[12]
port 133 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 D3[13]
port 134 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 D3[14]
port 135 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 D3[15]
port 136 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 D3[16]
port 137 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 D3[17]
port 138 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 D3[18]
port 139 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 D3[19]
port 140 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 D3[1]
port 141 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 D3[20]
port 142 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 D3[21]
port 143 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 D3[22]
port 144 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 D3[23]
port 145 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 D3[24]
port 146 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 D3[25]
port 147 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 D3[26]
port 148 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 D3[27]
port 149 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 D3[28]
port 150 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 D3[29]
port 151 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 D3[2]
port 152 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 D3[30]
port 153 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 D3[31]
port 154 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 D3[32]
port 155 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 D3[33]
port 156 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 D3[34]
port 157 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 D3[35]
port 158 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 D3[36]
port 159 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 D3[37]
port 160 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 D3[38]
port 161 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 D3[39]
port 162 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 D3[3]
port 163 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 D3[40]
port 164 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 D3[41]
port 165 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 D3[42]
port 166 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 D3[43]
port 167 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 D3[44]
port 168 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 D3[45]
port 169 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 D3[46]
port 170 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 D3[47]
port 171 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 D3[48]
port 172 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 D3[49]
port 173 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 D3[4]
port 174 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 D3[50]
port 175 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 D3[51]
port 176 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 D3[52]
port 177 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 D3[53]
port 178 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 D3[54]
port 179 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 D3[55]
port 180 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 D3[56]
port 181 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 D3[57]
port 182 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 D3[58]
port 183 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 D3[59]
port 184 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 D3[5]
port 185 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 D3[60]
port 186 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 D3[61]
port 187 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 D3[62]
port 188 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 D3[63]
port 189 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 D3[6]
port 190 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 D3[7]
port 191 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 D3[8]
port 192 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 D3[9]
port 193 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 DW[0]
port 194 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 DW[10]
port 195 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 DW[11]
port 196 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 DW[12]
port 197 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 DW[13]
port 198 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 DW[14]
port 199 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 DW[15]
port 200 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 DW[16]
port 201 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 DW[17]
port 202 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 DW[18]
port 203 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 DW[19]
port 204 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 DW[1]
port 205 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 DW[20]
port 206 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 DW[21]
port 207 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 DW[22]
port 208 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 DW[23]
port 209 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 DW[24]
port 210 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 DW[25]
port 211 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 DW[26]
port 212 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 DW[27]
port 213 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 DW[28]
port 214 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 DW[29]
port 215 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 DW[2]
port 216 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 DW[30]
port 217 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 DW[31]
port 218 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 DW[32]
port 219 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 DW[33]
port 220 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 DW[34]
port 221 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 DW[35]
port 222 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 DW[36]
port 223 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 DW[37]
port 224 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 DW[38]
port 225 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 DW[39]
port 226 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 DW[3]
port 227 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 DW[40]
port 228 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 DW[41]
port 229 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 DW[42]
port 230 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 DW[43]
port 231 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 DW[44]
port 232 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 DW[45]
port 233 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 DW[46]
port 234 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 DW[47]
port 235 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 DW[48]
port 236 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 DW[49]
port 237 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 DW[4]
port 238 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 DW[50]
port 239 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 DW[51]
port 240 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 DW[52]
port 241 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 DW[53]
port 242 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 DW[54]
port 243 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 DW[55]
port 244 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 DW[56]
port 245 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 DW[57]
port 246 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 DW[58]
port 247 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 DW[59]
port 248 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 DW[5]
port 249 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 DW[60]
port 250 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 DW[61]
port 251 nsew signal input
rlabel metal2 s 133234 0 133290 800 6 DW[62]
port 252 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 DW[63]
port 253 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 DW[6]
port 254 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 DW[7]
port 255 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 DW[8]
port 256 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 DW[9]
port 257 nsew signal input
rlabel metal2 s 13910 139200 13966 140000 6 R1[0]
port 258 nsew signal input
rlabel metal2 s 19246 139200 19302 140000 6 R1[1]
port 259 nsew signal input
rlabel metal2 s 24582 139200 24638 140000 6 R1[2]
port 260 nsew signal input
rlabel metal2 s 29918 139200 29974 140000 6 R1[3]
port 261 nsew signal input
rlabel metal2 s 35254 139200 35310 140000 6 R1[4]
port 262 nsew signal input
rlabel metal2 s 40590 139200 40646 140000 6 R1[5]
port 263 nsew signal input
rlabel metal2 s 45926 139200 45982 140000 6 R2[0]
port 264 nsew signal input
rlabel metal2 s 51262 139200 51318 140000 6 R2[1]
port 265 nsew signal input
rlabel metal2 s 56598 139200 56654 140000 6 R2[2]
port 266 nsew signal input
rlabel metal2 s 61934 139200 61990 140000 6 R2[3]
port 267 nsew signal input
rlabel metal2 s 67270 139200 67326 140000 6 R2[4]
port 268 nsew signal input
rlabel metal2 s 72606 139200 72662 140000 6 R2[5]
port 269 nsew signal input
rlabel metal2 s 77942 139200 77998 140000 6 R3[0]
port 270 nsew signal input
rlabel metal2 s 83278 139200 83334 140000 6 R3[1]
port 271 nsew signal input
rlabel metal2 s 88614 139200 88670 140000 6 R3[2]
port 272 nsew signal input
rlabel metal2 s 93950 139200 94006 140000 6 R3[3]
port 273 nsew signal input
rlabel metal2 s 99286 139200 99342 140000 6 R3[4]
port 274 nsew signal input
rlabel metal2 s 104622 139200 104678 140000 6 R3[5]
port 275 nsew signal input
rlabel metal2 s 109958 139200 110014 140000 6 RW[0]
port 276 nsew signal input
rlabel metal2 s 115294 139200 115350 140000 6 RW[1]
port 277 nsew signal input
rlabel metal2 s 120630 139200 120686 140000 6 RW[2]
port 278 nsew signal input
rlabel metal2 s 125966 139200 126022 140000 6 RW[3]
port 279 nsew signal input
rlabel metal2 s 131302 139200 131358 140000 6 RW[4]
port 280 nsew signal input
rlabel metal2 s 136638 139200 136694 140000 6 RW[5]
port 281 nsew signal input
rlabel metal4 s 19794 2128 20414 137680 6 VGND
port 282 nsew ground bidirectional
rlabel metal4 s 55794 2128 56414 137680 6 VGND
port 282 nsew ground bidirectional
rlabel metal4 s 91794 2128 92414 137680 6 VGND
port 282 nsew ground bidirectional
rlabel metal4 s 127794 2128 128414 137680 6 VGND
port 282 nsew ground bidirectional
rlabel metal4 s 1794 2128 2414 137680 6 VPWR
port 283 nsew power bidirectional
rlabel metal4 s 37794 2128 38414 137680 6 VPWR
port 283 nsew power bidirectional
rlabel metal4 s 73794 2128 74414 137680 6 VPWR
port 283 nsew power bidirectional
rlabel metal4 s 109794 2128 110414 137680 6 VPWR
port 283 nsew power bidirectional
rlabel metal2 s 8574 139200 8630 140000 6 WE
port 284 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 140000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 66787478
string GDS_FILE /scratch/mpw7/caravel_user_project/openlane/Microwatt_FP_DFFRFile/runs/22_09_06_08_57/results/signoff/Microwatt_FP_DFFRFile.magic.gds
string GDS_START 339312
<< end >>

